// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Dec 29 2020 20:58:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    tx,
    rx,
    reset);

    output tx;
    input rx;
    input reset;

    wire N__30069;
    wire N__30068;
    wire N__30067;
    wire N__30060;
    wire N__30059;
    wire N__30058;
    wire N__30051;
    wire N__30050;
    wire N__30049;
    wire N__30032;
    wire N__30031;
    wire N__30030;
    wire N__30029;
    wire N__30028;
    wire N__30027;
    wire N__30026;
    wire N__30025;
    wire N__30022;
    wire N__30021;
    wire N__30020;
    wire N__30019;
    wire N__30018;
    wire N__30017;
    wire N__30016;
    wire N__30015;
    wire N__30014;
    wire N__30013;
    wire N__30008;
    wire N__30003;
    wire N__29998;
    wire N__29997;
    wire N__29996;
    wire N__29995;
    wire N__29994;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29986;
    wire N__29985;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29973;
    wire N__29970;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29962;
    wire N__29959;
    wire N__29958;
    wire N__29955;
    wire N__29948;
    wire N__29947;
    wire N__29946;
    wire N__29945;
    wire N__29944;
    wire N__29943;
    wire N__29942;
    wire N__29931;
    wire N__29928;
    wire N__29927;
    wire N__29924;
    wire N__29919;
    wire N__29916;
    wire N__29915;
    wire N__29914;
    wire N__29913;
    wire N__29912;
    wire N__29911;
    wire N__29910;
    wire N__29901;
    wire N__29890;
    wire N__29887;
    wire N__29882;
    wire N__29879;
    wire N__29878;
    wire N__29873;
    wire N__29866;
    wire N__29861;
    wire N__29860;
    wire N__29859;
    wire N__29858;
    wire N__29857;
    wire N__29856;
    wire N__29855;
    wire N__29854;
    wire N__29853;
    wire N__29852;
    wire N__29851;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29839;
    wire N__29826;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29803;
    wire N__29790;
    wire N__29777;
    wire N__29770;
    wire N__29767;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29734;
    wire N__29733;
    wire N__29732;
    wire N__29731;
    wire N__29730;
    wire N__29729;
    wire N__29728;
    wire N__29725;
    wire N__29724;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29704;
    wire N__29703;
    wire N__29702;
    wire N__29701;
    wire N__29700;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29642;
    wire N__29637;
    wire N__29632;
    wire N__29629;
    wire N__29624;
    wire N__29609;
    wire N__29608;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29600;
    wire N__29599;
    wire N__29598;
    wire N__29597;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29586;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29566;
    wire N__29565;
    wire N__29564;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29545;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29527;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29498;
    wire N__29493;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29471;
    wire N__29470;
    wire N__29469;
    wire N__29468;
    wire N__29465;
    wire N__29464;
    wire N__29461;
    wire N__29460;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29452;
    wire N__29449;
    wire N__29448;
    wire N__29447;
    wire N__29442;
    wire N__29441;
    wire N__29438;
    wire N__29435;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29411;
    wire N__29408;
    wire N__29407;
    wire N__29402;
    wire N__29399;
    wire N__29390;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29371;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29353;
    wire N__29350;
    wire N__29349;
    wire N__29346;
    wire N__29345;
    wire N__29344;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29319;
    wire N__29314;
    wire N__29311;
    wire N__29310;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29282;
    wire N__29279;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29271;
    wire N__29270;
    wire N__29269;
    wire N__29268;
    wire N__29267;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29253;
    wire N__29250;
    wire N__29249;
    wire N__29246;
    wire N__29241;
    wire N__29240;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29216;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29204;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29180;
    wire N__29179;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29171;
    wire N__29168;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29153;
    wire N__29150;
    wire N__29149;
    wire N__29148;
    wire N__29143;
    wire N__29140;
    wire N__29139;
    wire N__29138;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29119;
    wire N__29114;
    wire N__29109;
    wire N__29102;
    wire N__29095;
    wire N__29092;
    wire N__29081;
    wire N__29080;
    wire N__29079;
    wire N__29076;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29070;
    wire N__29067;
    wire N__29066;
    wire N__29065;
    wire N__29062;
    wire N__29061;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29040;
    wire N__29039;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29024;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__28997;
    wire N__28982;
    wire N__28979;
    wire N__28978;
    wire N__28977;
    wire N__28974;
    wire N__28973;
    wire N__28972;
    wire N__28971;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28950;
    wire N__28949;
    wire N__28946;
    wire N__28943;
    wire N__28940;
    wire N__28939;
    wire N__28938;
    wire N__28937;
    wire N__28936;
    wire N__28935;
    wire N__28930;
    wire N__28925;
    wire N__28922;
    wire N__28917;
    wire N__28914;
    wire N__28905;
    wire N__28904;
    wire N__28901;
    wire N__28898;
    wire N__28893;
    wire N__28888;
    wire N__28885;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28867;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28859;
    wire N__28858;
    wire N__28857;
    wire N__28854;
    wire N__28851;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28823;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28803;
    wire N__28800;
    wire N__28793;
    wire N__28790;
    wire N__28789;
    wire N__28788;
    wire N__28787;
    wire N__28786;
    wire N__28785;
    wire N__28784;
    wire N__28783;
    wire N__28782;
    wire N__28781;
    wire N__28778;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28763;
    wire N__28762;
    wire N__28759;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28731;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28716;
    wire N__28713;
    wire N__28704;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28686;
    wire N__28683;
    wire N__28678;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28657;
    wire N__28654;
    wire N__28653;
    wire N__28652;
    wire N__28649;
    wire N__28648;
    wire N__28639;
    wire N__28638;
    wire N__28637;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28626;
    wire N__28625;
    wire N__28624;
    wire N__28621;
    wire N__28620;
    wire N__28619;
    wire N__28618;
    wire N__28615;
    wire N__28610;
    wire N__28605;
    wire N__28590;
    wire N__28589;
    wire N__28588;
    wire N__28583;
    wire N__28582;
    wire N__28579;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28563;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28547;
    wire N__28544;
    wire N__28543;
    wire N__28542;
    wire N__28541;
    wire N__28540;
    wire N__28539;
    wire N__28538;
    wire N__28537;
    wire N__28536;
    wire N__28535;
    wire N__28534;
    wire N__28533;
    wire N__28532;
    wire N__28531;
    wire N__28530;
    wire N__28529;
    wire N__28528;
    wire N__28527;
    wire N__28526;
    wire N__28525;
    wire N__28524;
    wire N__28523;
    wire N__28522;
    wire N__28521;
    wire N__28520;
    wire N__28519;
    wire N__28518;
    wire N__28517;
    wire N__28516;
    wire N__28515;
    wire N__28514;
    wire N__28513;
    wire N__28512;
    wire N__28511;
    wire N__28510;
    wire N__28509;
    wire N__28508;
    wire N__28507;
    wire N__28506;
    wire N__28505;
    wire N__28504;
    wire N__28503;
    wire N__28502;
    wire N__28501;
    wire N__28500;
    wire N__28499;
    wire N__28498;
    wire N__28497;
    wire N__28496;
    wire N__28495;
    wire N__28494;
    wire N__28493;
    wire N__28492;
    wire N__28491;
    wire N__28490;
    wire N__28489;
    wire N__28488;
    wire N__28487;
    wire N__28486;
    wire N__28485;
    wire N__28484;
    wire N__28483;
    wire N__28482;
    wire N__28481;
    wire N__28480;
    wire N__28479;
    wire N__28478;
    wire N__28477;
    wire N__28476;
    wire N__28475;
    wire N__28474;
    wire N__28473;
    wire N__28472;
    wire N__28471;
    wire N__28470;
    wire N__28469;
    wire N__28468;
    wire N__28467;
    wire N__28466;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28300;
    wire N__28297;
    wire N__28296;
    wire N__28293;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28274;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28254;
    wire N__28251;
    wire N__28246;
    wire N__28243;
    wire N__28238;
    wire N__28237;
    wire N__28236;
    wire N__28235;
    wire N__28234;
    wire N__28233;
    wire N__28232;
    wire N__28231;
    wire N__28230;
    wire N__28227;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28213;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28154;
    wire N__28151;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28129;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28094;
    wire N__28089;
    wire N__28082;
    wire N__28073;
    wire N__28072;
    wire N__28071;
    wire N__28068;
    wire N__28067;
    wire N__28066;
    wire N__28061;
    wire N__28058;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28035;
    wire N__28032;
    wire N__28029;
    wire N__28028;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__27999;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27958;
    wire N__27957;
    wire N__27954;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27940;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27918;
    wire N__27915;
    wire N__27914;
    wire N__27913;
    wire N__27908;
    wire N__27905;
    wire N__27900;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27886;
    wire N__27885;
    wire N__27884;
    wire N__27883;
    wire N__27882;
    wire N__27879;
    wire N__27878;
    wire N__27877;
    wire N__27876;
    wire N__27875;
    wire N__27874;
    wire N__27869;
    wire N__27864;
    wire N__27859;
    wire N__27858;
    wire N__27857;
    wire N__27856;
    wire N__27855;
    wire N__27854;
    wire N__27851;
    wire N__27850;
    wire N__27847;
    wire N__27840;
    wire N__27835;
    wire N__27832;
    wire N__27825;
    wire N__27818;
    wire N__27815;
    wire N__27810;
    wire N__27807;
    wire N__27800;
    wire N__27797;
    wire N__27790;
    wire N__27785;
    wire N__27784;
    wire N__27783;
    wire N__27782;
    wire N__27781;
    wire N__27780;
    wire N__27775;
    wire N__27774;
    wire N__27771;
    wire N__27770;
    wire N__27767;
    wire N__27766;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27756;
    wire N__27755;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27694;
    wire N__27691;
    wire N__27690;
    wire N__27687;
    wire N__27676;
    wire N__27671;
    wire N__27668;
    wire N__27663;
    wire N__27656;
    wire N__27655;
    wire N__27654;
    wire N__27653;
    wire N__27652;
    wire N__27651;
    wire N__27650;
    wire N__27649;
    wire N__27644;
    wire N__27639;
    wire N__27634;
    wire N__27633;
    wire N__27632;
    wire N__27631;
    wire N__27630;
    wire N__27629;
    wire N__27626;
    wire N__27625;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27582;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27550;
    wire N__27549;
    wire N__27546;
    wire N__27545;
    wire N__27540;
    wire N__27539;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27517;
    wire N__27514;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27490;
    wire N__27483;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27461;
    wire N__27460;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27452;
    wire N__27449;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27441;
    wire N__27440;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27415;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27382;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27352;
    wire N__27351;
    wire N__27348;
    wire N__27347;
    wire N__27344;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27327;
    wire N__27326;
    wire N__27325;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27303;
    wire N__27298;
    wire N__27297;
    wire N__27296;
    wire N__27293;
    wire N__27292;
    wire N__27291;
    wire N__27290;
    wire N__27287;
    wire N__27280;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27255;
    wire N__27250;
    wire N__27245;
    wire N__27238;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27214;
    wire N__27213;
    wire N__27210;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27196;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27188;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27146;
    wire N__27141;
    wire N__27136;
    wire N__27125;
    wire N__27124;
    wire N__27121;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26995;
    wire N__26994;
    wire N__26993;
    wire N__26988;
    wire N__26985;
    wire N__26984;
    wire N__26983;
    wire N__26980;
    wire N__26979;
    wire N__26976;
    wire N__26975;
    wire N__26974;
    wire N__26973;
    wire N__26972;
    wire N__26969;
    wire N__26964;
    wire N__26961;
    wire N__26960;
    wire N__26959;
    wire N__26958;
    wire N__26955;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26941;
    wire N__26940;
    wire N__26935;
    wire N__26932;
    wire N__26927;
    wire N__26922;
    wire N__26919;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26869;
    wire N__26868;
    wire N__26865;
    wire N__26864;
    wire N__26861;
    wire N__26860;
    wire N__26859;
    wire N__26858;
    wire N__26857;
    wire N__26856;
    wire N__26855;
    wire N__26854;
    wire N__26839;
    wire N__26830;
    wire N__26829;
    wire N__26828;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26813;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26797;
    wire N__26796;
    wire N__26795;
    wire N__26790;
    wire N__26785;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26764;
    wire N__26763;
    wire N__26762;
    wire N__26761;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26753;
    wire N__26752;
    wire N__26751;
    wire N__26750;
    wire N__26749;
    wire N__26748;
    wire N__26747;
    wire N__26744;
    wire N__26741;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26711;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26699;
    wire N__26694;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26674;
    wire N__26667;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26644;
    wire N__26639;
    wire N__26636;
    wire N__26635;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26606;
    wire N__26605;
    wire N__26604;
    wire N__26603;
    wire N__26602;
    wire N__26591;
    wire N__26590;
    wire N__26589;
    wire N__26588;
    wire N__26587;
    wire N__26586;
    wire N__26585;
    wire N__26584;
    wire N__26583;
    wire N__26582;
    wire N__26581;
    wire N__26580;
    wire N__26579;
    wire N__26578;
    wire N__26577;
    wire N__26576;
    wire N__26575;
    wire N__26574;
    wire N__26573;
    wire N__26572;
    wire N__26571;
    wire N__26570;
    wire N__26569;
    wire N__26568;
    wire N__26567;
    wire N__26566;
    wire N__26565;
    wire N__26564;
    wire N__26563;
    wire N__26562;
    wire N__26561;
    wire N__26560;
    wire N__26559;
    wire N__26558;
    wire N__26557;
    wire N__26556;
    wire N__26555;
    wire N__26554;
    wire N__26553;
    wire N__26550;
    wire N__26541;
    wire N__26532;
    wire N__26531;
    wire N__26530;
    wire N__26529;
    wire N__26528;
    wire N__26527;
    wire N__26526;
    wire N__26525;
    wire N__26524;
    wire N__26523;
    wire N__26522;
    wire N__26521;
    wire N__26520;
    wire N__26519;
    wire N__26518;
    wire N__26517;
    wire N__26516;
    wire N__26513;
    wire N__26512;
    wire N__26511;
    wire N__26510;
    wire N__26509;
    wire N__26508;
    wire N__26507;
    wire N__26506;
    wire N__26503;
    wire N__26502;
    wire N__26501;
    wire N__26486;
    wire N__26473;
    wire N__26456;
    wire N__26455;
    wire N__26454;
    wire N__26453;
    wire N__26452;
    wire N__26451;
    wire N__26450;
    wire N__26449;
    wire N__26434;
    wire N__26429;
    wire N__26426;
    wire N__26415;
    wire N__26414;
    wire N__26413;
    wire N__26412;
    wire N__26411;
    wire N__26410;
    wire N__26409;
    wire N__26408;
    wire N__26407;
    wire N__26406;
    wire N__26405;
    wire N__26404;
    wire N__26403;
    wire N__26402;
    wire N__26401;
    wire N__26400;
    wire N__26399;
    wire N__26398;
    wire N__26397;
    wire N__26396;
    wire N__26395;
    wire N__26394;
    wire N__26393;
    wire N__26390;
    wire N__26373;
    wire N__26364;
    wire N__26351;
    wire N__26350;
    wire N__26349;
    wire N__26348;
    wire N__26347;
    wire N__26346;
    wire N__26345;
    wire N__26344;
    wire N__26343;
    wire N__26340;
    wire N__26335;
    wire N__26332;
    wire N__26327;
    wire N__26312;
    wire N__26309;
    wire N__26302;
    wire N__26287;
    wire N__26286;
    wire N__26285;
    wire N__26284;
    wire N__26283;
    wire N__26282;
    wire N__26281;
    wire N__26280;
    wire N__26279;
    wire N__26264;
    wire N__26247;
    wire N__26246;
    wire N__26245;
    wire N__26244;
    wire N__26243;
    wire N__26242;
    wire N__26241;
    wire N__26240;
    wire N__26239;
    wire N__26238;
    wire N__26235;
    wire N__26230;
    wire N__26227;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26197;
    wire N__26196;
    wire N__26195;
    wire N__26194;
    wire N__26193;
    wire N__26192;
    wire N__26189;
    wire N__26184;
    wire N__26167;
    wire N__26162;
    wire N__26159;
    wire N__26142;
    wire N__26129;
    wire N__26126;
    wire N__26115;
    wire N__26096;
    wire N__26093;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26078;
    wire N__26075;
    wire N__26074;
    wire N__26073;
    wire N__26072;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26061;
    wire N__26060;
    wire N__26059;
    wire N__26058;
    wire N__26057;
    wire N__26056;
    wire N__26055;
    wire N__26054;
    wire N__26053;
    wire N__26050;
    wire N__26049;
    wire N__26048;
    wire N__26047;
    wire N__26044;
    wire N__26039;
    wire N__26036;
    wire N__26035;
    wire N__26032;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26021;
    wire N__26020;
    wire N__26019;
    wire N__26016;
    wire N__26013;
    wire N__26012;
    wire N__26011;
    wire N__26010;
    wire N__26007;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25986;
    wire N__25983;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25968;
    wire N__25965;
    wire N__25960;
    wire N__25957;
    wire N__25954;
    wire N__25951;
    wire N__25948;
    wire N__25943;
    wire N__25928;
    wire N__25927;
    wire N__25926;
    wire N__25923;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25901;
    wire N__25898;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25870;
    wire N__25869;
    wire N__25868;
    wire N__25863;
    wire N__25860;
    wire N__25853;
    wire N__25850;
    wire N__25841;
    wire N__25830;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25771;
    wire N__25768;
    wire N__25767;
    wire N__25766;
    wire N__25765;
    wire N__25764;
    wire N__25763;
    wire N__25762;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25742;
    wire N__25735;
    wire N__25732;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25716;
    wire N__25713;
    wire N__25708;
    wire N__25703;
    wire N__25694;
    wire N__25693;
    wire N__25692;
    wire N__25689;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25681;
    wire N__25680;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25661;
    wire N__25660;
    wire N__25657;
    wire N__25652;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25623;
    wire N__25616;
    wire N__25615;
    wire N__25612;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25600;
    wire N__25595;
    wire N__25594;
    wire N__25589;
    wire N__25586;
    wire N__25585;
    wire N__25580;
    wire N__25577;
    wire N__25576;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25553;
    wire N__25550;
    wire N__25549;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25513;
    wire N__25512;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25504;
    wire N__25503;
    wire N__25502;
    wire N__25501;
    wire N__25500;
    wire N__25499;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25484;
    wire N__25479;
    wire N__25474;
    wire N__25473;
    wire N__25468;
    wire N__25467;
    wire N__25466;
    wire N__25461;
    wire N__25452;
    wire N__25451;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25408;
    wire N__25399;
    wire N__25394;
    wire N__25391;
    wire N__25390;
    wire N__25387;
    wire N__25384;
    wire N__25379;
    wire N__25376;
    wire N__25375;
    wire N__25374;
    wire N__25373;
    wire N__25370;
    wire N__25369;
    wire N__25366;
    wire N__25363;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25345;
    wire N__25340;
    wire N__25339;
    wire N__25336;
    wire N__25335;
    wire N__25330;
    wire N__25329;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25308;
    wire N__25303;
    wire N__25298;
    wire N__25295;
    wire N__25286;
    wire N__25283;
    wire N__25282;
    wire N__25277;
    wire N__25274;
    wire N__25273;
    wire N__25268;
    wire N__25265;
    wire N__25264;
    wire N__25259;
    wire N__25256;
    wire N__25255;
    wire N__25250;
    wire N__25247;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25211;
    wire N__25208;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25168;
    wire N__25167;
    wire N__25166;
    wire N__25161;
    wire N__25160;
    wire N__25159;
    wire N__25158;
    wire N__25157;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25146;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25131;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25116;
    wire N__25109;
    wire N__25106;
    wire N__25099;
    wire N__25094;
    wire N__25091;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25061;
    wire N__25060;
    wire N__25059;
    wire N__25056;
    wire N__25055;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25016;
    wire N__25011;
    wire N__25010;
    wire N__25009;
    wire N__25004;
    wire N__25001;
    wire N__24996;
    wire N__24993;
    wire N__24986;
    wire N__24983;
    wire N__24982;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24970;
    wire N__24965;
    wire N__24962;
    wire N__24961;
    wire N__24956;
    wire N__24953;
    wire N__24952;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24940;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24893;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24881;
    wire N__24880;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24862;
    wire N__24861;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24847;
    wire N__24846;
    wire N__24845;
    wire N__24844;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24826;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24811;
    wire N__24804;
    wire N__24801;
    wire N__24796;
    wire N__24791;
    wire N__24782;
    wire N__24779;
    wire N__24778;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24760;
    wire N__24759;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24747;
    wire N__24746;
    wire N__24743;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24724;
    wire N__24719;
    wire N__24714;
    wire N__24711;
    wire N__24704;
    wire N__24703;
    wire N__24698;
    wire N__24695;
    wire N__24694;
    wire N__24689;
    wire N__24686;
    wire N__24685;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24650;
    wire N__24649;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24592;
    wire N__24591;
    wire N__24590;
    wire N__24589;
    wire N__24588;
    wire N__24585;
    wire N__24580;
    wire N__24577;
    wire N__24572;
    wire N__24567;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24481;
    wire N__24480;
    wire N__24479;
    wire N__24478;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24457;
    wire N__24452;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24414;
    wire N__24409;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24370;
    wire N__24369;
    wire N__24366;
    wire N__24365;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24319;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24285;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24259;
    wire N__24258;
    wire N__24255;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24247;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24227;
    wire N__24226;
    wire N__24221;
    wire N__24220;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24190;
    wire N__24189;
    wire N__24186;
    wire N__24183;
    wire N__24178;
    wire N__24175;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24156;
    wire N__24143;
    wire N__24142;
    wire N__24141;
    wire N__24140;
    wire N__24139;
    wire N__24138;
    wire N__24137;
    wire N__24136;
    wire N__24135;
    wire N__24134;
    wire N__24131;
    wire N__24126;
    wire N__24119;
    wire N__24114;
    wire N__24109;
    wire N__24106;
    wire N__24103;
    wire N__24098;
    wire N__24095;
    wire N__24090;
    wire N__24087;
    wire N__24082;
    wire N__24079;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24043;
    wire N__24040;
    wire N__24039;
    wire N__24036;
    wire N__24035;
    wire N__24032;
    wire N__24031;
    wire N__24030;
    wire N__24029;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24000;
    wire N__23997;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23981;
    wire N__23980;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23958;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23932;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23924;
    wire N__23921;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23881;
    wire N__23880;
    wire N__23873;
    wire N__23870;
    wire N__23865;
    wire N__23862;
    wire N__23857;
    wire N__23854;
    wire N__23847;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23794;
    wire N__23793;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23776;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23707;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23667;
    wire N__23666;
    wire N__23665;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23637;
    wire N__23634;
    wire N__23633;
    wire N__23630;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23597;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23554;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23523;
    wire N__23520;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23475;
    wire N__23472;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23410;
    wire N__23407;
    wire N__23406;
    wire N__23403;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23385;
    wire N__23378;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23366;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23335;
    wire N__23334;
    wire N__23333;
    wire N__23332;
    wire N__23331;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23314;
    wire N__23309;
    wire N__23308;
    wire N__23307;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23279;
    wire N__23278;
    wire N__23275;
    wire N__23268;
    wire N__23263;
    wire N__23260;
    wire N__23259;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23244;
    wire N__23239;
    wire N__23236;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23212;
    wire N__23209;
    wire N__23208;
    wire N__23205;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23172;
    wire N__23169;
    wire N__23162;
    wire N__23159;
    wire N__23158;
    wire N__23157;
    wire N__23156;
    wire N__23155;
    wire N__23154;
    wire N__23151;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23116;
    wire N__23113;
    wire N__23112;
    wire N__23111;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23085;
    wire N__23082;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23024;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23012;
    wire N__23009;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22997;
    wire N__22994;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22982;
    wire N__22979;
    wire N__22978;
    wire N__22977;
    wire N__22976;
    wire N__22975;
    wire N__22974;
    wire N__22973;
    wire N__22972;
    wire N__22971;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22957;
    wire N__22952;
    wire N__22945;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22906;
    wire N__22905;
    wire N__22902;
    wire N__22897;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22882;
    wire N__22881;
    wire N__22880;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22872;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22857;
    wire N__22854;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22840;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22798;
    wire N__22793;
    wire N__22790;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22765;
    wire N__22764;
    wire N__22763;
    wire N__22762;
    wire N__22761;
    wire N__22760;
    wire N__22759;
    wire N__22758;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22750;
    wire N__22747;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22732;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22711;
    wire N__22710;
    wire N__22709;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22674;
    wire N__22669;
    wire N__22666;
    wire N__22661;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22549;
    wire N__22548;
    wire N__22547;
    wire N__22546;
    wire N__22545;
    wire N__22544;
    wire N__22543;
    wire N__22542;
    wire N__22541;
    wire N__22540;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22529;
    wire N__22528;
    wire N__22527;
    wire N__22524;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22512;
    wire N__22511;
    wire N__22510;
    wire N__22509;
    wire N__22508;
    wire N__22507;
    wire N__22506;
    wire N__22505;
    wire N__22504;
    wire N__22503;
    wire N__22502;
    wire N__22501;
    wire N__22498;
    wire N__22497;
    wire N__22496;
    wire N__22493;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22485;
    wire N__22482;
    wire N__22481;
    wire N__22480;
    wire N__22479;
    wire N__22474;
    wire N__22469;
    wire N__22466;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22450;
    wire N__22447;
    wire N__22432;
    wire N__22415;
    wire N__22412;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22398;
    wire N__22389;
    wire N__22384;
    wire N__22379;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22361;
    wire N__22358;
    wire N__22353;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22327;
    wire N__22326;
    wire N__22323;
    wire N__22322;
    wire N__22321;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22313;
    wire N__22312;
    wire N__22311;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22303;
    wire N__22300;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22269;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22258;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22210;
    wire N__22203;
    wire N__22196;
    wire N__22187;
    wire N__22186;
    wire N__22183;
    wire N__22182;
    wire N__22179;
    wire N__22174;
    wire N__22171;
    wire N__22170;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22151;
    wire N__22150;
    wire N__22147;
    wire N__22146;
    wire N__22145;
    wire N__22144;
    wire N__22143;
    wire N__22142;
    wire N__22141;
    wire N__22140;
    wire N__22139;
    wire N__22136;
    wire N__22135;
    wire N__22134;
    wire N__22131;
    wire N__22126;
    wire N__22123;
    wire N__22116;
    wire N__22111;
    wire N__22110;
    wire N__22109;
    wire N__22108;
    wire N__22107;
    wire N__22104;
    wire N__22099;
    wire N__22094;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22078;
    wire N__22077;
    wire N__22074;
    wire N__22069;
    wire N__22064;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22049;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22033;
    wire N__22030;
    wire N__22019;
    wire N__22018;
    wire N__22013;
    wire N__22010;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21988;
    wire N__21985;
    wire N__21982;
    wire N__21977;
    wire N__21974;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21899;
    wire N__21896;
    wire N__21895;
    wire N__21894;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21876;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21868;
    wire N__21867;
    wire N__21866;
    wire N__21865;
    wire N__21864;
    wire N__21861;
    wire N__21856;
    wire N__21851;
    wire N__21846;
    wire N__21841;
    wire N__21836;
    wire N__21835;
    wire N__21834;
    wire N__21831;
    wire N__21830;
    wire N__21827;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21798;
    wire N__21795;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21734;
    wire N__21733;
    wire N__21728;
    wire N__21725;
    wire N__21724;
    wire N__21719;
    wire N__21716;
    wire N__21715;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21692;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21677;
    wire N__21674;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21662;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21647;
    wire N__21644;
    wire N__21643;
    wire N__21638;
    wire N__21635;
    wire N__21634;
    wire N__21633;
    wire N__21632;
    wire N__21631;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21612;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21600;
    wire N__21599;
    wire N__21596;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21566;
    wire N__21557;
    wire N__21554;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21542;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21530;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21509;
    wire N__21506;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21494;
    wire N__21493;
    wire N__21488;
    wire N__21485;
    wire N__21484;
    wire N__21479;
    wire N__21476;
    wire N__21475;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21425;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21413;
    wire N__21412;
    wire N__21407;
    wire N__21404;
    wire N__21403;
    wire N__21398;
    wire N__21395;
    wire N__21394;
    wire N__21389;
    wire N__21386;
    wire N__21385;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21373;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21314;
    wire N__21313;
    wire N__21312;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21184;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21142;
    wire N__21141;
    wire N__21140;
    wire N__21137;
    wire N__21136;
    wire N__21135;
    wire N__21132;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21115;
    wire N__21112;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21107;
    wire N__21104;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21084;
    wire N__21081;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21056;
    wire N__21047;
    wire N__21044;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21026;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20908;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20842;
    wire N__20841;
    wire N__20840;
    wire N__20839;
    wire N__20838;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20822;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20767;
    wire N__20766;
    wire N__20765;
    wire N__20764;
    wire N__20763;
    wire N__20762;
    wire N__20757;
    wire N__20752;
    wire N__20751;
    wire N__20750;
    wire N__20749;
    wire N__20748;
    wire N__20745;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20725;
    wire N__20722;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20588;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20576;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20564;
    wire N__20561;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20549;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20537;
    wire N__20536;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20513;
    wire N__20512;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20489;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20453;
    wire N__20450;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20438;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20420;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20405;
    wire N__20402;
    wire N__20401;
    wire N__20396;
    wire N__20393;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20381;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20366;
    wire N__20365;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20314;
    wire N__20313;
    wire N__20312;
    wire N__20311;
    wire N__20304;
    wire N__20299;
    wire N__20298;
    wire N__20297;
    wire N__20296;
    wire N__20295;
    wire N__20294;
    wire N__20293;
    wire N__20292;
    wire N__20291;
    wire N__20286;
    wire N__20281;
    wire N__20280;
    wire N__20279;
    wire N__20278;
    wire N__20277;
    wire N__20276;
    wire N__20273;
    wire N__20272;
    wire N__20271;
    wire N__20270;
    wire N__20269;
    wire N__20268;
    wire N__20267;
    wire N__20266;
    wire N__20265;
    wire N__20254;
    wire N__20249;
    wire N__20246;
    wire N__20245;
    wire N__20244;
    wire N__20241;
    wire N__20240;
    wire N__20239;
    wire N__20238;
    wire N__20233;
    wire N__20232;
    wire N__20231;
    wire N__20230;
    wire N__20229;
    wire N__20228;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20213;
    wire N__20208;
    wire N__20201;
    wire N__20196;
    wire N__20195;
    wire N__20194;
    wire N__20183;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20168;
    wire N__20167;
    wire N__20166;
    wire N__20165;
    wire N__20164;
    wire N__20163;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20151;
    wire N__20146;
    wire N__20145;
    wire N__20140;
    wire N__20133;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20125;
    wire N__20124;
    wire N__20123;
    wire N__20122;
    wire N__20121;
    wire N__20120;
    wire N__20119;
    wire N__20118;
    wire N__20115;
    wire N__20108;
    wire N__20105;
    wire N__20090;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20071;
    wire N__20060;
    wire N__20051;
    wire N__20046;
    wire N__20043;
    wire N__20034;
    wire N__20031;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19903;
    wire N__19902;
    wire N__19901;
    wire N__19898;
    wire N__19897;
    wire N__19896;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19856;
    wire N__19853;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19831;
    wire N__19828;
    wire N__19823;
    wire N__19818;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19744;
    wire N__19739;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19699;
    wire N__19694;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19682;
    wire N__19681;
    wire N__19680;
    wire N__19677;
    wire N__19672;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19642;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19600;
    wire N__19599;
    wire N__19598;
    wire N__19597;
    wire N__19596;
    wire N__19595;
    wire N__19594;
    wire N__19593;
    wire N__19592;
    wire N__19591;
    wire N__19590;
    wire N__19589;
    wire N__19588;
    wire N__19587;
    wire N__19586;
    wire N__19579;
    wire N__19568;
    wire N__19561;
    wire N__19550;
    wire N__19545;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19333;
    wire N__19330;
    wire N__19325;
    wire N__19324;
    wire N__19323;
    wire N__19320;
    wire N__19315;
    wire N__19312;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19258;
    wire N__19257;
    wire N__19256;
    wire N__19255;
    wire N__19252;
    wire N__19247;
    wire N__19246;
    wire N__19245;
    wire N__19244;
    wire N__19241;
    wire N__19240;
    wire N__19239;
    wire N__19238;
    wire N__19237;
    wire N__19236;
    wire N__19233;
    wire N__19232;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19217;
    wire N__19216;
    wire N__19215;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19200;
    wire N__19199;
    wire N__19198;
    wire N__19191;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19168;
    wire N__19167;
    wire N__19166;
    wire N__19163;
    wire N__19158;
    wire N__19155;
    wire N__19154;
    wire N__19153;
    wire N__19148;
    wire N__19143;
    wire N__19140;
    wire N__19135;
    wire N__19130;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19102;
    wire N__19097;
    wire N__19092;
    wire N__19073;
    wire N__19072;
    wire N__19071;
    wire N__19070;
    wire N__19067;
    wire N__19066;
    wire N__19061;
    wire N__19060;
    wire N__19059;
    wire N__19058;
    wire N__19057;
    wire N__19056;
    wire N__19055;
    wire N__19054;
    wire N__19053;
    wire N__19052;
    wire N__19051;
    wire N__19050;
    wire N__19049;
    wire N__19048;
    wire N__19047;
    wire N__19046;
    wire N__19045;
    wire N__19044;
    wire N__19043;
    wire N__19042;
    wire N__19039;
    wire N__19038;
    wire N__19037;
    wire N__19032;
    wire N__19029;
    wire N__19024;
    wire N__19019;
    wire N__19018;
    wire N__19017;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__18999;
    wire N__18994;
    wire N__18987;
    wire N__18984;
    wire N__18983;
    wire N__18980;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18963;
    wire N__18962;
    wire N__18955;
    wire N__18950;
    wire N__18947;
    wire N__18942;
    wire N__18937;
    wire N__18932;
    wire N__18925;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18910;
    wire N__18909;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18884;
    wire N__18881;
    wire N__18876;
    wire N__18871;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18851;
    wire N__18836;
    wire N__18835;
    wire N__18834;
    wire N__18833;
    wire N__18832;
    wire N__18831;
    wire N__18830;
    wire N__18827;
    wire N__18822;
    wire N__18819;
    wire N__18818;
    wire N__18817;
    wire N__18816;
    wire N__18815;
    wire N__18808;
    wire N__18805;
    wire N__18804;
    wire N__18799;
    wire N__18792;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18778;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18766;
    wire N__18765;
    wire N__18762;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18750;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18727;
    wire N__18724;
    wire N__18713;
    wire N__18710;
    wire N__18709;
    wire N__18704;
    wire N__18701;
    wire N__18700;
    wire N__18695;
    wire N__18692;
    wire N__18691;
    wire N__18686;
    wire N__18683;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18665;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18653;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18641;
    wire N__18638;
    wire N__18637;
    wire N__18632;
    wire N__18629;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18617;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18605;
    wire N__18604;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18592;
    wire N__18589;
    wire N__18586;
    wire N__18581;
    wire N__18580;
    wire N__18575;
    wire N__18572;
    wire N__18571;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18559;
    wire N__18554;
    wire N__18551;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18536;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18524;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18452;
    wire N__18451;
    wire N__18446;
    wire N__18443;
    wire N__18442;
    wire N__18437;
    wire N__18434;
    wire N__18433;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18421;
    wire N__18420;
    wire N__18415;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18385;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18367;
    wire N__18362;
    wire N__18361;
    wire N__18360;
    wire N__18359;
    wire N__18358;
    wire N__18357;
    wire N__18356;
    wire N__18355;
    wire N__18354;
    wire N__18353;
    wire N__18352;
    wire N__18351;
    wire N__18350;
    wire N__18347;
    wire N__18342;
    wire N__18341;
    wire N__18340;
    wire N__18339;
    wire N__18336;
    wire N__18335;
    wire N__18334;
    wire N__18331;
    wire N__18322;
    wire N__18319;
    wire N__18318;
    wire N__18317;
    wire N__18316;
    wire N__18315;
    wire N__18314;
    wire N__18313;
    wire N__18308;
    wire N__18307;
    wire N__18306;
    wire N__18305;
    wire N__18304;
    wire N__18301;
    wire N__18296;
    wire N__18295;
    wire N__18294;
    wire N__18293;
    wire N__18284;
    wire N__18283;
    wire N__18282;
    wire N__18281;
    wire N__18280;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18268;
    wire N__18263;
    wire N__18262;
    wire N__18259;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18251;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18218;
    wire N__18215;
    wire N__18214;
    wire N__18213;
    wire N__18210;
    wire N__18209;
    wire N__18208;
    wire N__18205;
    wire N__18202;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18194;
    wire N__18193;
    wire N__18192;
    wire N__18189;
    wire N__18182;
    wire N__18179;
    wire N__18164;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18144;
    wire N__18141;
    wire N__18128;
    wire N__18115;
    wire N__18110;
    wire N__18103;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18073;
    wire N__18072;
    wire N__18069;
    wire N__18064;
    wire N__18059;
    wire N__18058;
    wire N__18055;
    wire N__18054;
    wire N__18053;
    wire N__18052;
    wire N__18051;
    wire N__18048;
    wire N__18047;
    wire N__18046;
    wire N__18043;
    wire N__18038;
    wire N__18035;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18027;
    wire N__18026;
    wire N__18025;
    wire N__18024;
    wire N__18023;
    wire N__18022;
    wire N__18021;
    wire N__18020;
    wire N__18019;
    wire N__18018;
    wire N__18017;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18003;
    wire N__18002;
    wire N__17999;
    wire N__17998;
    wire N__17997;
    wire N__17996;
    wire N__17991;
    wire N__17986;
    wire N__17983;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17975;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17967;
    wire N__17966;
    wire N__17965;
    wire N__17964;
    wire N__17963;
    wire N__17962;
    wire N__17951;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17934;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17926;
    wire N__17921;
    wire N__17918;
    wire N__17905;
    wire N__17902;
    wire N__17889;
    wire N__17886;
    wire N__17881;
    wire N__17878;
    wire N__17869;
    wire N__17864;
    wire N__17857;
    wire N__17848;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17812;
    wire N__17809;
    wire N__17808;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17794;
    wire N__17791;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17774;
    wire N__17771;
    wire N__17770;
    wire N__17769;
    wire N__17768;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17749;
    wire N__17746;
    wire N__17745;
    wire N__17742;
    wire N__17737;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17677;
    wire N__17674;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17614;
    wire N__17613;
    wire N__17612;
    wire N__17611;
    wire N__17610;
    wire N__17607;
    wire N__17602;
    wire N__17599;
    wire N__17598;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17582;
    wire N__17579;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17530;
    wire N__17529;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17517;
    wire N__17514;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17491;
    wire N__17488;
    wire N__17487;
    wire N__17484;
    wire N__17483;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17468;
    wire N__17459;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17416;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17344;
    wire N__17343;
    wire N__17340;
    wire N__17335;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17306;
    wire N__17305;
    wire N__17304;
    wire N__17297;
    wire N__17294;
    wire N__17293;
    wire N__17290;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17201;
    wire N__17198;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17159;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17151;
    wire N__17148;
    wire N__17145;
    wire N__17142;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17107;
    wire N__17102;
    wire N__17101;
    wire N__17098;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17083;
    wire N__17078;
    wire N__17077;
    wire N__17076;
    wire N__17073;
    wire N__17068;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17058;
    wire N__17053;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16990;
    wire N__16987;
    wire N__16984;
    wire N__16981;
    wire N__16976;
    wire N__16975;
    wire N__16974;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16949;
    wire N__16948;
    wire N__16945;
    wire N__16944;
    wire N__16943;
    wire N__16942;
    wire N__16941;
    wire N__16940;
    wire N__16939;
    wire N__16936;
    wire N__16935;
    wire N__16934;
    wire N__16933;
    wire N__16932;
    wire N__16931;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16923;
    wire N__16922;
    wire N__16917;
    wire N__16912;
    wire N__16909;
    wire N__16902;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16882;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16858;
    wire N__16857;
    wire N__16856;
    wire N__16855;
    wire N__16854;
    wire N__16853;
    wire N__16850;
    wire N__16849;
    wire N__16848;
    wire N__16845;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16837;
    wire N__16828;
    wire N__16821;
    wire N__16812;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16798;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16780;
    wire N__16777;
    wire N__16774;
    wire N__16771;
    wire N__16770;
    wire N__16769;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16736;
    wire N__16735;
    wire N__16734;
    wire N__16733;
    wire N__16732;
    wire N__16731;
    wire N__16730;
    wire N__16729;
    wire N__16720;
    wire N__16713;
    wire N__16710;
    wire N__16703;
    wire N__16702;
    wire N__16701;
    wire N__16700;
    wire N__16699;
    wire N__16698;
    wire N__16697;
    wire N__16694;
    wire N__16693;
    wire N__16684;
    wire N__16677;
    wire N__16674;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16657;
    wire N__16654;
    wire N__16651;
    wire N__16648;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16632;
    wire N__16631;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16615;
    wire N__16610;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16594;
    wire N__16589;
    wire N__16586;
    wire N__16585;
    wire N__16584;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16565;
    wire N__16562;
    wire N__16561;
    wire N__16556;
    wire N__16553;
    wire N__16552;
    wire N__16547;
    wire N__16544;
    wire N__16543;
    wire N__16538;
    wire N__16535;
    wire N__16534;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16498;
    wire N__16497;
    wire N__16494;
    wire N__16493;
    wire N__16492;
    wire N__16489;
    wire N__16488;
    wire N__16485;
    wire N__16484;
    wire N__16481;
    wire N__16480;
    wire N__16477;
    wire N__16476;
    wire N__16473;
    wire N__16470;
    wire N__16463;
    wire N__16460;
    wire N__16451;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16435;
    wire N__16434;
    wire N__16433;
    wire N__16432;
    wire N__16429;
    wire N__16422;
    wire N__16419;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16390;
    wire N__16387;
    wire N__16384;
    wire N__16383;
    wire N__16382;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16370;
    wire N__16369;
    wire N__16366;
    wire N__16361;
    wire N__16358;
    wire N__16357;
    wire N__16354;
    wire N__16353;
    wire N__16348;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16316;
    wire N__16313;
    wire N__16312;
    wire N__16311;
    wire N__16310;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16298;
    wire N__16295;
    wire N__16294;
    wire N__16293;
    wire N__16290;
    wire N__16285;
    wire N__16282;
    wire N__16281;
    wire N__16278;
    wire N__16275;
    wire N__16268;
    wire N__16265;
    wire N__16256;
    wire N__16253;
    wire N__16252;
    wire N__16251;
    wire N__16248;
    wire N__16243;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16228;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16204;
    wire N__16203;
    wire N__16202;
    wire N__16201;
    wire N__16198;
    wire N__16197;
    wire N__16196;
    wire N__16195;
    wire N__16194;
    wire N__16191;
    wire N__16186;
    wire N__16173;
    wire N__16172;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16164;
    wire N__16163;
    wire N__16162;
    wire N__16159;
    wire N__16154;
    wire N__16149;
    wire N__16144;
    wire N__16141;
    wire N__16136;
    wire N__16135;
    wire N__16134;
    wire N__16127;
    wire N__16124;
    wire N__16119;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16105;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16083;
    wire N__16080;
    wire N__16073;
    wire N__16072;
    wire N__16071;
    wire N__16068;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16053;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16024;
    wire N__16021;
    wire N__16018;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15991;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15981;
    wire N__15978;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15964;
    wire N__15963;
    wire N__15962;
    wire N__15961;
    wire N__15960;
    wire N__15957;
    wire N__15954;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15911;
    wire N__15908;
    wire N__15905;
    wire N__15900;
    wire N__15893;
    wire N__15890;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15882;
    wire N__15879;
    wire N__15876;
    wire N__15875;
    wire N__15874;
    wire N__15873;
    wire N__15870;
    wire N__15865;
    wire N__15862;
    wire N__15861;
    wire N__15860;
    wire N__15857;
    wire N__15854;
    wire N__15851;
    wire N__15846;
    wire N__15843;
    wire N__15840;
    wire N__15835;
    wire N__15830;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15814;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15766;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15737;
    wire N__15734;
    wire N__15731;
    wire N__15728;
    wire N__15727;
    wire N__15726;
    wire N__15723;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15673;
    wire N__15672;
    wire N__15671;
    wire N__15668;
    wire N__15667;
    wire N__15664;
    wire N__15663;
    wire N__15660;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15640;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15628;
    wire N__15627;
    wire N__15626;
    wire N__15625;
    wire N__15624;
    wire N__15623;
    wire N__15622;
    wire N__15621;
    wire N__15620;
    wire N__15619;
    wire N__15612;
    wire N__15595;
    wire N__15594;
    wire N__15591;
    wire N__15590;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15575;
    wire N__15566;
    wire N__15563;
    wire N__15562;
    wire N__15561;
    wire N__15560;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15544;
    wire N__15543;
    wire N__15542;
    wire N__15539;
    wire N__15536;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15528;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15517;
    wire N__15512;
    wire N__15509;
    wire N__15508;
    wire N__15505;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15489;
    wire N__15486;
    wire N__15483;
    wire N__15476;
    wire N__15471;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15451;
    wire N__15450;
    wire N__15447;
    wire N__15442;
    wire N__15437;
    wire N__15434;
    wire N__15433;
    wire N__15432;
    wire N__15425;
    wire N__15424;
    wire N__15423;
    wire N__15420;
    wire N__15419;
    wire N__15418;
    wire N__15417;
    wire N__15412;
    wire N__15409;
    wire N__15402;
    wire N__15395;
    wire N__15392;
    wire N__15391;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15379;
    wire N__15376;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15355;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15337;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15325;
    wire N__15324;
    wire N__15317;
    wire N__15314;
    wire N__15313;
    wire N__15312;
    wire N__15311;
    wire N__15308;
    wire N__15303;
    wire N__15300;
    wire N__15295;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15274;
    wire N__15271;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15235;
    wire N__15234;
    wire N__15233;
    wire N__15232;
    wire N__15231;
    wire N__15230;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15196;
    wire N__15187;
    wire N__15186;
    wire N__15185;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15169;
    wire N__15164;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15142;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15127;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15094;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15076;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15055;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15040;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15019;
    wire N__15018;
    wire N__15017;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14977;
    wire N__14976;
    wire N__14973;
    wire N__14968;
    wire N__14967;
    wire N__14964;
    wire N__14961;
    wire N__14958;
    wire N__14953;
    wire N__14948;
    wire N__14945;
    wire N__14944;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14850;
    wire N__14849;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14833;
    wire N__14830;
    wire N__14827;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14778;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14768;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14752;
    wire N__14749;
    wire N__14746;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14697;
    wire N__14696;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14665;
    wire N__14662;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14622;
    wire N__14619;
    wire N__14616;
    wire N__14615;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14594;
    wire N__14591;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14553;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14534;
    wire N__14531;
    wire N__14526;
    wire N__14523;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14494;
    wire N__14489;
    wire N__14486;
    wire N__14485;
    wire N__14480;
    wire N__14477;
    wire N__14476;
    wire N__14471;
    wire N__14468;
    wire N__14467;
    wire N__14462;
    wire N__14459;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14449;
    wire N__14444;
    wire N__14441;
    wire N__14440;
    wire N__14435;
    wire N__14432;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14422;
    wire N__14417;
    wire N__14416;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14374;
    wire N__14373;
    wire N__14372;
    wire N__14371;
    wire N__14370;
    wire N__14369;
    wire N__14368;
    wire N__14367;
    wire N__14366;
    wire N__14365;
    wire N__14362;
    wire N__14357;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14321;
    wire N__14318;
    wire N__14313;
    wire N__14306;
    wire N__14303;
    wire N__14300;
    wire N__14297;
    wire N__14294;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14270;
    wire N__14269;
    wire N__14266;
    wire N__14265;
    wire N__14264;
    wire N__14261;
    wire N__14260;
    wire N__14257;
    wire N__14256;
    wire N__14255;
    wire N__14252;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14220;
    wire N__14213;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14197;
    wire N__14196;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14188;
    wire N__14187;
    wire N__14186;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14174;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14124;
    wire N__14117;
    wire N__14114;
    wire N__14113;
    wire N__14112;
    wire N__14109;
    wire N__14106;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14094;
    wire N__14091;
    wire N__14084;
    wire N__14083;
    wire N__14080;
    wire N__14079;
    wire N__14076;
    wire N__14071;
    wire N__14070;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14054;
    wire N__14053;
    wire N__14048;
    wire N__14045;
    wire N__14044;
    wire N__14041;
    wire N__14040;
    wire N__14039;
    wire N__14038;
    wire N__14037;
    wire N__14036;
    wire N__14035;
    wire N__14034;
    wire N__14033;
    wire N__14032;
    wire N__14031;
    wire N__14030;
    wire N__14029;
    wire N__14028;
    wire N__14027;
    wire N__14026;
    wire N__14025;
    wire N__14024;
    wire N__14023;
    wire N__14022;
    wire N__14021;
    wire N__14020;
    wire N__14019;
    wire N__14018;
    wire N__14017;
    wire N__14016;
    wire N__14015;
    wire N__14014;
    wire N__14013;
    wire N__14012;
    wire N__14011;
    wire N__14010;
    wire N__14009;
    wire N__14008;
    wire N__14007;
    wire N__14006;
    wire N__14005;
    wire N__14004;
    wire N__14003;
    wire N__14002;
    wire N__14001;
    wire N__14000;
    wire N__13999;
    wire N__13998;
    wire N__13997;
    wire N__13996;
    wire N__13995;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13983;
    wire N__13980;
    wire N__13979;
    wire N__13978;
    wire N__13977;
    wire N__13976;
    wire N__13963;
    wire N__13950;
    wire N__13943;
    wire N__13930;
    wire N__13921;
    wire N__13908;
    wire N__13907;
    wire N__13906;
    wire N__13905;
    wire N__13904;
    wire N__13903;
    wire N__13902;
    wire N__13901;
    wire N__13900;
    wire N__13899;
    wire N__13898;
    wire N__13897;
    wire N__13896;
    wire N__13893;
    wire N__13880;
    wire N__13867;
    wire N__13864;
    wire N__13859;
    wire N__13856;
    wire N__13847;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13833;
    wire N__13830;
    wire N__13817;
    wire N__13804;
    wire N__13801;
    wire N__13794;
    wire N__13785;
    wire N__13778;
    wire N__13773;
    wire N__13770;
    wire N__13765;
    wire N__13762;
    wire N__13757;
    wire N__13748;
    wire N__13747;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13721;
    wire N__13720;
    wire N__13717;
    wire N__13716;
    wire N__13715;
    wire N__13714;
    wire N__13713;
    wire N__13712;
    wire N__13711;
    wire N__13708;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13696;
    wire N__13695;
    wire N__13694;
    wire N__13693;
    wire N__13692;
    wire N__13691;
    wire N__13690;
    wire N__13689;
    wire N__13688;
    wire N__13687;
    wire N__13686;
    wire N__13685;
    wire N__13684;
    wire N__13683;
    wire N__13682;
    wire N__13681;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13671;
    wire N__13670;
    wire N__13669;
    wire N__13668;
    wire N__13667;
    wire N__13666;
    wire N__13665;
    wire N__13664;
    wire N__13663;
    wire N__13658;
    wire N__13649;
    wire N__13648;
    wire N__13647;
    wire N__13646;
    wire N__13645;
    wire N__13644;
    wire N__13643;
    wire N__13642;
    wire N__13639;
    wire N__13636;
    wire N__13635;
    wire N__13634;
    wire N__13633;
    wire N__13632;
    wire N__13631;
    wire N__13628;
    wire N__13627;
    wire N__13624;
    wire N__13623;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13612;
    wire N__13611;
    wire N__13610;
    wire N__13609;
    wire N__13608;
    wire N__13607;
    wire N__13606;
    wire N__13605;
    wire N__13604;
    wire N__13603;
    wire N__13602;
    wire N__13601;
    wire N__13600;
    wire N__13599;
    wire N__13590;
    wire N__13583;
    wire N__13570;
    wire N__13557;
    wire N__13552;
    wire N__13551;
    wire N__13550;
    wire N__13549;
    wire N__13546;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13520;
    wire N__13515;
    wire N__13512;
    wire N__13503;
    wire N__13492;
    wire N__13479;
    wire N__13466;
    wire N__13463;
    wire N__13454;
    wire N__13447;
    wire N__13444;
    wire N__13439;
    wire N__13436;
    wire N__13415;
    wire N__13412;
    wire N__13407;
    wire N__13404;
    wire N__13397;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13384;
    wire N__13381;
    wire N__13376;
    wire N__13373;
    wire N__13372;
    wire N__13371;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13363;
    wire N__13362;
    wire N__13361;
    wire N__13360;
    wire N__13357;
    wire N__13354;
    wire N__13349;
    wire N__13346;
    wire N__13345;
    wire N__13342;
    wire N__13339;
    wire N__13336;
    wire N__13331;
    wire N__13330;
    wire N__13329;
    wire N__13328;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13290;
    wire N__13285;
    wire N__13276;
    wire N__13273;
    wire N__13262;
    wire N__13261;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13130;
    wire N__13129;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13090;
    wire N__13087;
    wire N__13086;
    wire N__13083;
    wire N__13080;
    wire N__13077;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13065;
    wire N__13062;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13048;
    wire N__13045;
    wire N__13042;
    wire N__13041;
    wire N__13040;
    wire N__13037;
    wire N__13032;
    wire N__13029;
    wire N__13022;
    wire N__13019;
    wire N__13018;
    wire N__13015;
    wire N__13014;
    wire N__13013;
    wire N__13010;
    wire N__13007;
    wire N__13002;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12988;
    wire N__12987;
    wire N__12984;
    wire N__12983;
    wire N__12978;
    wire N__12975;
    wire N__12972;
    wire N__12967;
    wire N__12962;
    wire N__12959;
    wire N__12958;
    wire N__12957;
    wire N__12954;
    wire N__12949;
    wire N__12948;
    wire N__12943;
    wire N__12940;
    wire N__12937;
    wire N__12932;
    wire N__12929;
    wire N__12928;
    wire N__12927;
    wire N__12926;
    wire N__12925;
    wire N__12924;
    wire N__12923;
    wire N__12920;
    wire N__12907;
    wire N__12904;
    wire N__12901;
    wire N__12898;
    wire N__12893;
    wire N__12890;
    wire N__12887;
    wire N__12886;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12871;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12838;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12826;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12808;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12796;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12784;
    wire N__12781;
    wire N__12780;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12768;
    wire N__12765;
    wire N__12758;
    wire N__12757;
    wire N__12756;
    wire N__12753;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12729;
    wire N__12726;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12712;
    wire N__12711;
    wire N__12710;
    wire N__12707;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12686;
    wire N__12683;
    wire N__12682;
    wire N__12681;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12669;
    wire N__12666;
    wire N__12659;
    wire N__12658;
    wire N__12655;
    wire N__12654;
    wire N__12651;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12633;
    wire N__12630;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12616;
    wire N__12613;
    wire N__12612;
    wire N__12611;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12595;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12559;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12544;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12466;
    wire N__12465;
    wire N__12464;
    wire N__12455;
    wire N__12452;
    wire N__12451;
    wire N__12450;
    wire N__12447;
    wire N__12446;
    wire N__12441;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12425;
    wire N__12422;
    wire N__12421;
    wire N__12420;
    wire N__12419;
    wire N__12416;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12398;
    wire N__12389;
    wire N__12388;
    wire N__12383;
    wire N__12380;
    wire N__12379;
    wire N__12378;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12364;
    wire N__12359;
    wire N__12358;
    wire N__12357;
    wire N__12356;
    wire N__12355;
    wire N__12354;
    wire N__12353;
    wire N__12348;
    wire N__12345;
    wire N__12336;
    wire N__12329;
    wire N__12328;
    wire N__12327;
    wire N__12326;
    wire N__12317;
    wire N__12314;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12302;
    wire N__12299;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12133;
    wire N__12132;
    wire N__12129;
    wire N__12128;
    wire N__12121;
    wire N__12118;
    wire N__12115;
    wire N__12112;
    wire N__12109;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12048;
    wire N__12041;
    wire N__12040;
    wire N__12039;
    wire N__12036;
    wire N__12031;
    wire N__12028;
    wire N__12023;
    wire N__12022;
    wire N__12021;
    wire N__12014;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__11999;
    wire N__11996;
    wire N__11995;
    wire N__11992;
    wire N__11989;
    wire N__11984;
    wire N__11981;
    wire N__11980;
    wire N__11977;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11900;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11888;
    wire N__11887;
    wire N__11886;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11876;
    wire N__11871;
    wire N__11868;
    wire N__11861;
    wire N__11858;
    wire N__11855;
    wire N__11854;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11846;
    wire N__11845;
    wire N__11844;
    wire N__11843;
    wire N__11830;
    wire N__11827;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11800;
    wire N__11795;
    wire N__11794;
    wire N__11793;
    wire N__11792;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11777;
    wire N__11774;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11743;
    wire N__11738;
    wire N__11735;
    wire N__11734;
    wire N__11729;
    wire N__11726;
    wire N__11725;
    wire N__11720;
    wire N__11717;
    wire N__11716;
    wire N__11711;
    wire N__11708;
    wire N__11707;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11692;
    wire N__11689;
    wire N__11686;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11657;
    wire N__11656;
    wire N__11651;
    wire N__11648;
    wire N__11647;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11605;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11585;
    wire N__11584;
    wire N__11583;
    wire N__11580;
    wire N__11579;
    wire N__11576;
    wire N__11571;
    wire N__11568;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11503;
    wire N__11500;
    wire N__11499;
    wire N__11492;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11444;
    wire N__11443;
    wire N__11438;
    wire N__11435;
    wire N__11432;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11408;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11314;
    wire N__11309;
    wire N__11306;
    wire N__11305;
    wire N__11300;
    wire N__11297;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11246;
    wire N__11243;
    wire N__11242;
    wire N__11241;
    wire N__11240;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11222;
    wire N__11219;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11207;
    wire N__11204;
    wire N__11203;
    wire N__11202;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11188;
    wire N__11187;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11171;
    wire N__11170;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11158;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11135;
    wire N__11132;
    wire N__11131;
    wire N__11130;
    wire N__11127;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11069;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11057;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11042;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11025;
    wire N__11018;
    wire N__11015;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11003;
    wire N__11002;
    wire N__10999;
    wire N__10996;
    wire N__10991;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10979;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10967;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10922;
    wire N__10919;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10907;
    wire N__10906;
    wire N__10903;
    wire N__10900;
    wire N__10895;
    wire N__10894;
    wire N__10891;
    wire N__10888;
    wire N__10885;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10850;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10838;
    wire N__10837;
    wire N__10834;
    wire N__10831;
    wire N__10828;
    wire N__10823;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10804;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10783;
    wire N__10778;
    wire N__10777;
    wire N__10774;
    wire N__10771;
    wire N__10766;
    wire N__10763;
    wire N__10762;
    wire N__10757;
    wire N__10754;
    wire N__10753;
    wire N__10748;
    wire N__10745;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10727;
    wire N__10724;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10687;
    wire N__10684;
    wire N__10681;
    wire N__10676;
    wire N__10675;
    wire N__10670;
    wire N__10667;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10655;
    wire N__10652;
    wire N__10651;
    wire N__10646;
    wire N__10643;
    wire N__10642;
    wire N__10637;
    wire N__10634;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10613;
    wire N__10610;
    wire N__10609;
    wire N__10606;
    wire N__10603;
    wire N__10600;
    wire N__10595;
    wire N__10592;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10580;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10559;
    wire N__10556;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10544;
    wire N__10541;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10531;
    wire N__10526;
    wire N__10523;
    wire N__10522;
    wire N__10519;
    wire N__10516;
    wire N__10511;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10498;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10486;
    wire N__10483;
    wire N__10480;
    wire N__10475;
    wire N__10474;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10454;
    wire N__10451;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10439;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10427;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10415;
    wire N__10412;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10400;
    wire N__10397;
    wire N__10396;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10373;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10361;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10348;
    wire N__10343;
    wire N__10342;
    wire N__10339;
    wire N__10336;
    wire N__10333;
    wire N__10330;
    wire N__10325;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10313;
    wire N__10312;
    wire N__10309;
    wire N__10304;
    wire N__10301;
    wire N__10300;
    wire N__10295;
    wire N__10292;
    wire N__10291;
    wire N__10286;
    wire N__10283;
    wire N__10282;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10259;
    wire N__10258;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10195;
    wire N__10190;
    wire N__10187;
    wire N__10186;
    wire N__10183;
    wire N__10180;
    wire N__10175;
    wire N__10172;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10157;
    wire N__10154;
    wire N__10153;
    wire N__10148;
    wire N__10145;
    wire N__10144;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10126;
    wire N__10121;
    wire N__10118;
    wire N__10117;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10103;
    wire N__10102;
    wire N__10097;
    wire N__10094;
    wire N__10093;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10081;
    wire N__10078;
    wire N__10075;
    wire VCCG0;
    wire \tok.C_stk.n5447_cascade_ ;
    wire \tok.C_stk.tail_3 ;
    wire \tok.tail_11 ;
    wire \tok.C_stk.tail_19 ;
    wire \tok.tail_27 ;
    wire \tok.C_stk.tail_35 ;
    wire \tok.C_stk.n5456_cascade_ ;
    wire \tok.C_stk.tail_0 ;
    wire \tok.tail_8 ;
    wire \tok.C_stk.tail_16 ;
    wire \tok.tail_24 ;
    wire \tok.C_stk.tail_32 ;
    wire bfn_1_3_0_;
    wire \tok.uart.n4827 ;
    wire \tok.uart.n4828 ;
    wire \tok.uart.n4829 ;
    wire \tok.uart.n4830 ;
    wire \tok.uart.n4831 ;
    wire \tok.uart.n4832 ;
    wire bfn_1_4_0_;
    wire \tok.uart.n4814 ;
    wire \tok.uart.n4815 ;
    wire \tok.uart.n4816 ;
    wire \tok.uart.n4817 ;
    wire \tok.uart.n4818 ;
    wire \tok.uart.n4819 ;
    wire \tok.uart.n4820 ;
    wire \tok.uart.n4821 ;
    wire bfn_1_5_0_;
    wire \tok.C_stk.n5453_cascade_ ;
    wire \tok.C_stk.tail_1 ;
    wire \tok.tail_9 ;
    wire \tok.C_stk.tail_17 ;
    wire \tok.tail_25 ;
    wire \tok.C_stk.tail_33 ;
    wire \tok.C_stk.n5450_cascade_ ;
    wire \tok.C_stk.tail_2 ;
    wire \tok.tail_10 ;
    wire \tok.C_stk.tail_18 ;
    wire \tok.tail_26 ;
    wire \tok.C_stk.tail_34 ;
    wire \tok.tail_43 ;
    wire \tok.tail_42 ;
    wire \tok.tail_41 ;
    wire \tok.tail_40 ;
    wire \tok.tail_60 ;
    wire \tok.tail_51 ;
    wire \tok.tail_59 ;
    wire \tok.tail_50 ;
    wire \tok.tail_58 ;
    wire \tok.tail_49 ;
    wire \tok.tail_57 ;
    wire \tok.tail_48 ;
    wire \tok.tail_56 ;
    wire \tok.tail_63 ;
    wire \tok.C_stk.n5435_cascade_ ;
    wire \tok.C_stk.tail_7 ;
    wire \tok.tail_15 ;
    wire \tok.C_stk.tail_23 ;
    wire \tok.tail_31 ;
    wire \tok.C_stk.tail_39 ;
    wire \tok.tail_55 ;
    wire \tok.tail_47 ;
    wire \tok.tail_12 ;
    wire \tok.C_stk.tail_20 ;
    wire \tok.tail_28 ;
    wire \tok.C_stk.tail_36 ;
    wire \tok.tail_52 ;
    wire \tok.tail_44 ;
    wire bfn_2_2_0_;
    wire \tok.uart.n4822 ;
    wire \tok.uart.n4823 ;
    wire \tok.uart.n4824 ;
    wire \tok.uart.n4825 ;
    wire \tok.uart.n4826 ;
    wire \tok.uart.rxclkcounter_5 ;
    wire \tok.uart.rxclkcounter_3 ;
    wire \tok.uart.rxclkcounter_2 ;
    wire n813_cascade_;
    wire n971;
    wire \tok.uart.rxclkcounter_6 ;
    wire \tok.uart.rxclkcounter_0 ;
    wire \tok.uart.rxclkcounter_4 ;
    wire \tok.uart.rxclkcounter_1 ;
    wire \tok.uart.n12_adj_640 ;
    wire \tok.uart.sentbits_3 ;
    wire \tok.uart.txclkcounter_5 ;
    wire \tok.uart.txclkcounter_2 ;
    wire \tok.uart.txclkcounter_8 ;
    wire \tok.uart.txclkcounter_3 ;
    wire \tok.uart.sentbits_2 ;
    wire \tok.uart.txclkcounter_4 ;
    wire \tok.uart.txclkcounter_7 ;
    wire \tok.uart.txclkcounter_6 ;
    wire \tok.uart.txclkcounter_0 ;
    wire \tok.uart.txclkcounter_1 ;
    wire \tok.uart.n5418_cascade_ ;
    wire \tok.uart.n12 ;
    wire txtick_cascade_;
    wire \tok.tail_61 ;
    wire \tok.uart.n2_cascade_ ;
    wire \tok.uart.rxclkcounter_6__N_477 ;
    wire \tok.uart.bytephase_2 ;
    wire \tok.uart.n13_cascade_ ;
    wire \tok.uart.bytephase_4 ;
    wire bytephase_5__N_510;
    wire \tok.uart.bytephase_0 ;
    wire n813;
    wire \tok.uart.bytephase_1 ;
    wire \tok.c_stk_r_2 ;
    wire \tok.ram.n5585 ;
    wire \tok.n3_adj_645_cascade_ ;
    wire \tok.n83 ;
    wire \tok.n5603 ;
    wire \tok.n31_adj_795_cascade_ ;
    wire \tok.n5473 ;
    wire \tok.C_stk.n5441_cascade_ ;
    wire \tok.C_stk.tail_5 ;
    wire \tok.tail_13 ;
    wire \tok.C_stk.tail_21 ;
    wire \tok.tail_29 ;
    wire \tok.C_stk.tail_37 ;
    wire \tok.tail_53 ;
    wire \tok.tail_45 ;
    wire \tok.tc_0 ;
    wire n92;
    wire n92_cascade_;
    wire \tok.tc_3 ;
    wire \tok.n13_adj_646 ;
    wire n10_cascade_;
    wire \tok.tc_2 ;
    wire n10;
    wire \tok.n36_cascade_ ;
    wire \tok.n83_adj_842_cascade_ ;
    wire \tok.ram.n5597_cascade_ ;
    wire \tok.c_stk_r_0 ;
    wire \tok.n5583 ;
    wire \tok.n3_adj_863_cascade_ ;
    wire \tok.n5_adj_864 ;
    wire \tok.n83_adj_714_cascade_ ;
    wire \tok.tc_7 ;
    wire \tok.ram.n5600_cascade_ ;
    wire \tok.c_stk_r_7 ;
    wire \tok.n5511 ;
    wire \tok.n3_adj_719_cascade_ ;
    wire \tok.n5_adj_720_cascade_ ;
    wire n92_adj_869;
    wire n92_adj_869_cascade_;
    wire \tok.n5507 ;
    wire \tok.C_stk.tail_4 ;
    wire \tok.tail_62 ;
    wire \tok.C_stk.n5444 ;
    wire \tok.tail_54 ;
    wire \tok.C_stk.tail_38 ;
    wire \tok.tail_46 ;
    wire sender_1;
    wire tx_c;
    wire \tok.A_stk.tail_17 ;
    wire \tok.A_stk.tail_33 ;
    wire \tok.A_stk.tail_49 ;
    wire \tok.A_stk.tail_65 ;
    wire \tok.A_stk.tail_81 ;
    wire \tok.A_stk.tail_1 ;
    wire \tok.A_stk_delta_1__N_4_cascade_ ;
    wire \tok.depth_1_cascade_ ;
    wire \tok.n37 ;
    wire \tok.n2585_cascade_ ;
    wire \tok.n59 ;
    wire \tok.depth_3 ;
    wire \tok.n60 ;
    wire \tok.depth_2 ;
    wire \tok.n807 ;
    wire n23_cascade_;
    wire txtick;
    wire \tok.uart.sentbits_0 ;
    wire \tok.uart.sentbits_1 ;
    wire \tok.uart.n1023 ;
    wire \tok.uart.n1093 ;
    wire \tok.n4_adj_707 ;
    wire \tok.n42 ;
    wire \tok.n5287 ;
    wire \tok.n5287_cascade_ ;
    wire \tok.n7 ;
    wire \tok.n5312_cascade_ ;
    wire \tok.n15_adj_817_cascade_ ;
    wire \tok.n898 ;
    wire \tok.n898_cascade_ ;
    wire \tok.uart.n6 ;
    wire \tok.ram.n5608_cascade_ ;
    wire \tok.c_stk_r_5 ;
    wire \tok.n83_adj_678_cascade_ ;
    wire \tok.n3_adj_683 ;
    wire \tok.n5483_cascade_ ;
    wire \tok.n5_adj_684_cascade_ ;
    wire n92_adj_868_cascade_;
    wire \tok.tc_5 ;
    wire n92_adj_868;
    wire \tok.table_wr_data_4 ;
    wire \tok.table_wr_data_15 ;
    wire \tok.table_wr_data_14 ;
    wire \tok.table_wr_data_3 ;
    wire \tok.table_wr_data_2 ;
    wire \tok.table_wr_data_1 ;
    wire \tok.table_wr_data_5 ;
    wire \tok.table_wr_data_7 ;
    wire \tok.table_wr_data_13 ;
    wire \tok.table_wr_data_12 ;
    wire \tok.table_wr_data_11 ;
    wire \tok.table_wr_data_10 ;
    wire \tok.table_wr_data_9 ;
    wire \tok.table_wr_data_8 ;
    wire \tok.table_wr_data_0 ;
    wire \tok.n8_adj_790 ;
    wire \tok.n14_adj_644_cascade_ ;
    wire \tok.n7_adj_785 ;
    wire tail_97;
    wire tail_113;
    wire \tok.n27_adj_828_cascade_ ;
    wire \tok.n27_adj_831_cascade_ ;
    wire \tok.n27_adj_833_cascade_ ;
    wire \tok.n27_adj_825 ;
    wire \tok.n5285_cascade_ ;
    wire \tok.n1_adj_715_cascade_ ;
    wire \tok.n190 ;
    wire \tok.n890 ;
    wire \tok.n10_adj_763_cascade_ ;
    wire \tok.n5338 ;
    wire \tok.n5340 ;
    wire \tok.A_stk_delta_1__N_4 ;
    wire \tok.n61 ;
    wire \tok.n4_adj_813 ;
    wire \tok.n13_adj_691_cascade_ ;
    wire n10_adj_871_cascade_;
    wire \tok.tc_6 ;
    wire \tok.ram.n5605_cascade_ ;
    wire \tok.n3_adj_690 ;
    wire \tok.n83_adj_687_cascade_ ;
    wire \tok.n5505 ;
    wire n10_adj_871;
    wire \tok.n83_adj_848_cascade_ ;
    wire \tok.c_stk_r_1 ;
    wire \tok.ram.n5594_cascade_ ;
    wire \tok.n5610 ;
    wire \tok.n3_cascade_ ;
    wire \tok.n13_cascade_ ;
    wire \tok.uart.n5 ;
    wire \tok.key_rd_10 ;
    wire \tok.key_rd_12 ;
    wire \tok.n21_adj_733_cascade_ ;
    wire \tok.key_rd_7 ;
    wire \tok.key_rd_2 ;
    wire \tok.n22_adj_721 ;
    wire \tok.n23_adj_731 ;
    wire \tok.n24_adj_651 ;
    wire \tok.key_rd_14 ;
    wire \tok.key_rd_15 ;
    wire \tok.key_rd_9 ;
    wire \tok.key_rd_11 ;
    wire tc_0;
    wire \tok.tc_plus_1_0 ;
    wire bfn_5_8_0_;
    wire \tok.tc_plus_1_1 ;
    wire \tok.n4754 ;
    wire tc_2;
    wire \tok.tc_plus_1_2 ;
    wire \tok.n4755 ;
    wire tc_3;
    wire \tok.n4756 ;
    wire \tok.n4757 ;
    wire tc_5;
    wire \tok.tc_plus_1_5 ;
    wire \tok.n4758 ;
    wire \tok.n4759 ;
    wire tc_7;
    wire \tok.n4760 ;
    wire \tok.tc_plus_1_7 ;
    wire \tok.n9_adj_798 ;
    wire \tok.n5293 ;
    wire \tok.n5391 ;
    wire \tok.n14_adj_688_cascade_ ;
    wire \tok.n2735_cascade_ ;
    wire \tok.n1_adj_850_cascade_ ;
    wire \tok.n26_adj_750 ;
    wire \tok.n5380 ;
    wire \tok.n8_adj_805 ;
    wire \tok.n11_adj_793 ;
    wire \tok.n5271_cascade_ ;
    wire \tok.n5318 ;
    wire \tok.n11_adj_694 ;
    wire \tok.n15_adj_695 ;
    wire uart_rx_data_4;
    wire \tok.n12_adj_826 ;
    wire \tok.n11_adj_788 ;
    wire sender_2;
    wire \tok.uart.sender_3 ;
    wire \tok.uart.sender_4 ;
    wire \tok.uart.sender_5 ;
    wire \tok.uart.sender_6 ;
    wire \tok.uart.sender_7 ;
    wire sender_9;
    wire n23;
    wire \tok.uart.sender_8 ;
    wire \tok.uart.n1017 ;
    wire \tok.C_stk.n602 ;
    wire \tok.n241 ;
    wire \tok.C_stk.n5438_cascade_ ;
    wire tc_6;
    wire \tok.c_stk_r_6 ;
    wire \tok.C_stk.tail_6 ;
    wire \tok.n2515 ;
    wire \tok.tail_14 ;
    wire \tok.tail_30 ;
    wire \tok.n29_adj_787 ;
    wire \tok.C_stk.tail_22 ;
    wire \tok.C_stk_delta_0 ;
    wire reset_c;
    wire \tok.A_stk.tail_16 ;
    wire \tok.A_stk.tail_32 ;
    wire \tok.A_stk.tail_48 ;
    wire \tok.A_stk.tail_64 ;
    wire tail_112;
    wire \tok.A_stk.tail_80 ;
    wire tail_96;
    wire \tok.A_stk.tail_0 ;
    wire bfn_6_3_0_;
    wire \tok.n4747 ;
    wire \tok.n4748 ;
    wire \tok.n4749 ;
    wire \tok.idx_4 ;
    wire \tok.n33_adj_819 ;
    wire \tok.n4750 ;
    wire \tok.idx_5 ;
    wire \tok.n33_adj_811 ;
    wire \tok.n4751 ;
    wire \tok.idx_6 ;
    wire \tok.n33_adj_804 ;
    wire \tok.n4752 ;
    wire \tok.idx_7 ;
    wire \tok.n4753 ;
    wire \tok.n33_adj_801 ;
    wire \tok.n5_cascade_ ;
    wire \tok.n5 ;
    wire \tok.n33 ;
    wire \tok.n27_cascade_ ;
    wire \tok.idx_0 ;
    wire \tok.n83_adj_652_cascade_ ;
    wire \tok.c_stk_r_3 ;
    wire \tok.ram.n5580_cascade_ ;
    wire \tok.n5460 ;
    wire \tok.n3_adj_659_cascade_ ;
    wire \tok.tc_plus_1_3 ;
    wire \tok.n13_adj_660_cascade_ ;
    wire n92_adj_867;
    wire \tok.n17_adj_777 ;
    wire \tok.n4_adj_778_cascade_ ;
    wire \tok.n26_adj_760_cascade_ ;
    wire \tok.n30_adj_761 ;
    wire \tok.n5587_cascade_ ;
    wire \tok.key_rd_8 ;
    wire \tok.n28_adj_755 ;
    wire \tok.n26_adj_756_cascade_ ;
    wire \tok.n27_adj_757 ;
    wire \tok.found_slot_N_145 ;
    wire \tok.found_slot ;
    wire \tok.write_slot ;
    wire \tok.key_rd_3 ;
    wire \tok.key_rd_5 ;
    wire \tok.n20 ;
    wire \tok.n18_adj_759 ;
    wire \tok.key_rd_1 ;
    wire \tok.key_rd_4 ;
    wire \tok.n25_adj_758 ;
    wire \tok.key_rd_0 ;
    wire \tok.key_rd_6 ;
    wire \tok.n5590 ;
    wire uart_rx_data_6;
    wire \tok.n6_adj_843 ;
    wire \tok.n31_adj_844_cascade_ ;
    wire uart_rx_data_3;
    wire capture_4;
    wire \tok.tc_plus_1_6 ;
    wire \tok.table_wr_data_6 ;
    wire \tok.n10_adj_747 ;
    wire \tok.n2635 ;
    wire \tok.n11 ;
    wire \tok.n2697 ;
    wire \tok.n15_adj_789 ;
    wire \tok.n2520 ;
    wire \tok.n10_adj_803 ;
    wire \tok.n2520_cascade_ ;
    wire \tok.n9_adj_802 ;
    wire \tok.table_rd_3 ;
    wire \tok.n2661_cascade_ ;
    wire \tok.n10_adj_845 ;
    wire \tok.n9_adj_847_cascade_ ;
    wire \tok.n14_adj_701 ;
    wire \tok.n5429 ;
    wire \tok.n5406 ;
    wire \tok.n5433_cascade_ ;
    wire \tok.n5272 ;
    wire \tok.n10_adj_796 ;
    wire \tok.n14_adj_807 ;
    wire \tok.n5175 ;
    wire n10_adj_866;
    wire tc_1;
    wire \tok.tc_1 ;
    wire \tok.n2_adj_808 ;
    wire \tok.n5423 ;
    wire \tok.n42_adj_751 ;
    wire capture_9;
    wire \tok.n2609 ;
    wire \tok.n4_adj_712 ;
    wire \tok.ram.n5577_cascade_ ;
    wire \tok.n101 ;
    wire \tok.n3_adj_672 ;
    wire \tok.n820 ;
    wire \tok.n5298 ;
    wire \tok.n13_adj_673_cascade_ ;
    wire \tok.tc_plus_1_4 ;
    wire n10_adj_870_cascade_;
    wire \tok.tc_4 ;
    wire stall_;
    wire n10_adj_870;
    wire tc_4;
    wire \tok.c_stk_r_4 ;
    wire \tok.n83_adj_665_cascade_ ;
    wire \tok.n5487 ;
    wire \tok.A_stk.tail_94 ;
    wire \tok.A_stk.tail_78 ;
    wire \tok.A_stk.tail_62 ;
    wire \tok.A_stk.tail_46 ;
    wire \tok.A_stk.tail_30 ;
    wire tail_127;
    wire \tok.n33_adj_814 ;
    wire \tok.n62 ;
    wire \tok.n1_adj_715 ;
    wire \tok.depth_0_cascade_ ;
    wire \tok.n5408 ;
    wire \tok.n33_adj_816 ;
    wire \tok.n27_adj_818_cascade_ ;
    wire \tok.idx_2 ;
    wire \tok.stall ;
    wire \tok.n33_adj_821 ;
    wire \tok.search_clk ;
    wire \tok.n27_adj_822_cascade_ ;
    wire \tok.idx_3 ;
    wire \tok.n2699 ;
    wire \tok.n5282 ;
    wire \tok.n27_adj_815 ;
    wire \tok.idx_1 ;
    wire rd_15__N_301_cascade_;
    wire \tok.n797 ;
    wire \tok.n2585 ;
    wire A_stk_delta_1_cascade_;
    wire tail_110;
    wire tail_126;
    wire tail_111;
    wire rx_c;
    wire \tok.uart.n5235 ;
    wire \tok.uart.bytephase_5 ;
    wire \tok.uart.bytephase_3 ;
    wire \tok.uart.n5374 ;
    wire \tok.key_rd_13 ;
    wire \tok.n14_adj_647 ;
    wire capture_0;
    wire capture_1;
    wire uart_rx_data_0;
    wire \tok.n6_adj_794_cascade_ ;
    wire \tok.table_rd_6 ;
    wire \tok.n5553_cascade_ ;
    wire \tok.table_rd_14 ;
    wire \tok.table_rd_12 ;
    wire \tok.n14_adj_735_cascade_ ;
    wire \tok.n6_adj_754 ;
    wire \tok.table_rd_4 ;
    wire \tok.n16_adj_851_cascade_ ;
    wire \tok.n17_adj_853 ;
    wire \tok.n5562_cascade_ ;
    wire \tok.n13_adj_852 ;
    wire \tok.n14_adj_854 ;
    wire capture_3;
    wire \tok.table_rd_0 ;
    wire \tok.n31 ;
    wire \tok.n5463_cascade_ ;
    wire \tok.n2607 ;
    wire \tok.n14_adj_765 ;
    wire \tok.table_rd_1 ;
    wire \tok.n5334_cascade_ ;
    wire \tok.n5462 ;
    wire \tok.n5566 ;
    wire \tok.n5561 ;
    wire \tok.n9_adj_766 ;
    wire \tok.n10_adj_643 ;
    wire \tok.uart_tx_busy ;
    wire \tok.n15_adj_655_cascade_ ;
    wire \tok.uart_stall ;
    wire \tok.uart_rx_valid ;
    wire \tok.uart.n953 ;
    wire \tok.n15_adj_667_cascade_ ;
    wire \tok.table_rd_2 ;
    wire \tok.n28_adj_771_cascade_ ;
    wire \tok.n5470 ;
    wire \tok.n5467_cascade_ ;
    wire \tok.n34 ;
    wire \tok.n82_cascade_ ;
    wire \tok.n878 ;
    wire \tok.n8_adj_846 ;
    wire \tok.n41 ;
    wire bfn_7_13_0_;
    wire \tok.T_1 ;
    wire \tok.n4761 ;
    wire \tok.n15_adj_664 ;
    wire \tok.n4762 ;
    wire \tok.n82 ;
    wire \tok.T_3 ;
    wire \tok.n11_adj_830 ;
    wire \tok.n4763 ;
    wire \tok.n212 ;
    wire \tok.n4764 ;
    wire \tok.n4765 ;
    wire \tok.n210 ;
    wire \tok.n4766 ;
    wire \tok.n4767 ;
    wire \tok.n4768 ;
    wire bfn_7_14_0_;
    wire tail_121;
    wire tail_105;
    wire \tok.A_stk.tail_89 ;
    wire \tok.A_stk.tail_73 ;
    wire \tok.A_stk.tail_57 ;
    wire \tok.A_stk.tail_41 ;
    wire \tok.A_stk.tail_25 ;
    wire \tok.A_stk.tail_9 ;
    wire tail_115;
    wire tail_99;
    wire \tok.A_stk.tail_84 ;
    wire \tok.A_stk.tail_68 ;
    wire \tok.A_stk.tail_52 ;
    wire \tok.A_stk.tail_36 ;
    wire tail_119;
    wire \tok.A_stk.tail_20 ;
    wire tail_103;
    wire \tok.A_stk.tail_71 ;
    wire \tok.A_stk.tail_87 ;
    wire tail_120;
    wire \tok.A_stk.tail_88 ;
    wire tail_104;
    wire \tok.n9_adj_786 ;
    wire \tok.table_rd_7 ;
    wire \tok.n5548_cascade_ ;
    wire \tok.n285_cascade_ ;
    wire \tok.n12_adj_824 ;
    wire \tok.n1_adj_862_cascade_ ;
    wire \tok.T_6 ;
    wire \tok.T_4 ;
    wire \tok.T_5 ;
    wire \tok.n6_adj_650_cascade_ ;
    wire \tok.n13_adj_654_cascade_ ;
    wire \tok.n5547 ;
    wire \tok.n5546_cascade_ ;
    wire \tok.n14 ;
    wire \tok.n17 ;
    wire \tok.n13_adj_641_cascade_ ;
    wire \tok.n5552 ;
    wire \tok.n5551_cascade_ ;
    wire \tok.n5465 ;
    wire bfn_8_7_0_;
    wire \tok.n4784 ;
    wire \tok.n4785 ;
    wire \tok.n4_adj_806 ;
    wire \tok.n4786 ;
    wire \tok.n5564 ;
    wire \tok.n4787 ;
    wire \tok.n4788 ;
    wire \tok.n5554 ;
    wire \tok.n4789 ;
    wire \tok.n5549 ;
    wire \tok.n4790 ;
    wire \tok.n4791 ;
    wire bfn_8_8_0_;
    wire \tok.n4792 ;
    wire \tok.n4793 ;
    wire \tok.n4794 ;
    wire \tok.n5_adj_734 ;
    wire \tok.n4795 ;
    wire \tok.n4796 ;
    wire \tok.n5_adj_716 ;
    wire \tok.n4797 ;
    wire \tok.n399 ;
    wire \tok.n4798 ;
    wire \tok.n8_adj_837 ;
    wire \tok.n5574 ;
    wire \tok.n5334 ;
    wire \tok.n5254 ;
    wire \tok.n5414_cascade_ ;
    wire \tok.n8_adj_767 ;
    wire \tok.n904_cascade_ ;
    wire \tok.n11_adj_840 ;
    wire \tok.n5346_cascade_ ;
    wire \tok.n16_adj_810 ;
    wire \tok.n14_adj_841_cascade_ ;
    wire \tok.n5571 ;
    wire \tok.n5569 ;
    wire \tok.n45_adj_849 ;
    wire \tok.n4848 ;
    wire \tok.table_rd_9 ;
    wire \tok.n45_cascade_ ;
    wire \tok.n39 ;
    wire \tok.n11_adj_680 ;
    wire \tok.table_rd_10 ;
    wire \tok.n14_adj_679 ;
    wire \tok.n45_adj_696 ;
    wire \tok.n39_adj_697_cascade_ ;
    wire \tok.n10_adj_700_cascade_ ;
    wire \tok.n5536 ;
    wire \tok.n11_adj_730 ;
    wire \tok.n26_cascade_ ;
    wire \tok.tc__7__N_134 ;
    wire \tok.n25_adj_710 ;
    wire \tok.n28_adj_708 ;
    wire \tok.n27_adj_709 ;
    wire \tok.n14_adj_764 ;
    wire \tok.T_0 ;
    wire \tok.n10_adj_858 ;
    wire \tok.table_rd_13 ;
    wire \tok.n5_adj_732 ;
    wire \tok.n12_adj_779 ;
    wire \tok.n14_adj_776_cascade_ ;
    wire \tok.n13_adj_780 ;
    wire \tok.n20_adj_784_cascade_ ;
    wire \tok.n9_adj_781 ;
    wire \tok.n5_adj_713 ;
    wire \tok.table_rd_15 ;
    wire \tok.n16_adj_782 ;
    wire \tok.n209 ;
    wire \tok.n14_adj_658 ;
    wire \tok.n2_adj_775 ;
    wire tail_118;
    wire tail_100;
    wire tail_116;
    wire tail_114;
    wire tail_98;
    wire \tok.A_stk.tail_82 ;
    wire \tok.A_stk.tail_72 ;
    wire tail_102;
    wire \tok.A_stk.tail_70 ;
    wire \tok.A_stk.tail_86 ;
    wire \tok.A_stk.tail_55 ;
    wire \tok.A_stk.tail_39 ;
    wire \tok.A_stk.tail_83 ;
    wire \tok.A_stk.tail_4 ;
    wire \tok.A_stk.tail_6 ;
    wire \tok.A_stk.tail_54 ;
    wire \tok.A_stk.tail_22 ;
    wire \tok.A_stk.tail_38 ;
    wire \tok.A_stk.tail_23 ;
    wire \tok.n3_adj_692 ;
    wire bfn_9_6_0_;
    wire \tok.n4799 ;
    wire \tok.n4800 ;
    wire \tok.n22_adj_829 ;
    wire \tok.n4801 ;
    wire \tok.n10_adj_827 ;
    wire \tok.n4802 ;
    wire \tok.n4803 ;
    wire \tok.n10_adj_820 ;
    wire \tok.n4804 ;
    wire \tok.n10_adj_653 ;
    wire \tok.n4805 ;
    wire \tok.n4806 ;
    wire bfn_9_7_0_;
    wire \tok.n4807 ;
    wire \tok.n20_adj_663 ;
    wire \tok.n4808 ;
    wire \tok.n4809 ;
    wire \tok.n10_adj_738 ;
    wire \tok.n4810 ;
    wire \tok.n4811 ;
    wire \tok.n10_adj_768 ;
    wire \tok.n4812 ;
    wire \tok.write_flag ;
    wire \tok.n4813 ;
    wire \tok.n5516 ;
    wire \tok.n18_adj_739 ;
    wire \tok.n12_adj_737_cascade_ ;
    wire \tok.n1_cascade_ ;
    wire \tok.n17_adj_656 ;
    wire \tok.n12 ;
    wire uart_rx_data_7;
    wire \tok.n177 ;
    wire \tok.n17_adj_812 ;
    wire \tok.n9_adj_838 ;
    wire \tok.n23_adj_682 ;
    wire \tok.n25 ;
    wire \tok.n4_cascade_ ;
    wire \tok.n5350 ;
    wire capture_2;
    wire \tok.n9 ;
    wire \tok.n5342_cascade_ ;
    wire \tok.n10_adj_686 ;
    wire \tok.A_low_1 ;
    wire \tok.n5336 ;
    wire \tok.table_rd_11 ;
    wire \tok.n5_adj_726 ;
    wire \tok.n13_adj_724_cascade_ ;
    wire \tok.n12_adj_723 ;
    wire \tok.n5534 ;
    wire \tok.n16 ;
    wire \tok.n20_adj_729_cascade_ ;
    wire \tok.n9_adj_725 ;
    wire \tok.n5531 ;
    wire \tok.n2 ;
    wire \tok.n14_adj_722 ;
    wire \tok.n20_adj_740 ;
    wire \tok.n5527_cascade_ ;
    wire \tok.n5513 ;
    wire \tok.n5539 ;
    wire \tok.n5348 ;
    wire \tok.n13_adj_746_cascade_ ;
    wire \tok.n12_adj_745 ;
    wire \tok.n5525 ;
    wire \tok.n16_adj_749 ;
    wire \tok.n20_adj_753_cascade_ ;
    wire \tok.n5522 ;
    wire \tok.n8 ;
    wire \tok.n14_adj_744 ;
    wire \tok.n9_adj_748 ;
    wire \tok.n2_adj_743 ;
    wire \tok.n204_cascade_ ;
    wire \tok.n16_adj_741 ;
    wire tail_125;
    wire tail_109;
    wire \tok.A_stk.tail_93 ;
    wire \tok.A_stk.tail_77 ;
    wire \tok.A_stk.tail_61 ;
    wire \tok.A_stk.tail_45 ;
    wire \tok.A_stk.tail_29 ;
    wire \tok.A_stk.tail_13 ;
    wire tail_123;
    wire tail_107;
    wire \tok.A_stk.tail_91 ;
    wire tail_124;
    wire tail_108;
    wire \tok.A_stk.tail_92 ;
    wire \tok.A_stk.tail_76 ;
    wire \tok.A_stk.tail_60 ;
    wire \tok.A_stk.tail_7 ;
    wire \tok.A_stk.tail_2 ;
    wire \tok.A_stk.tail_18 ;
    wire \tok.A_stk.tail_34 ;
    wire \tok.A_stk.tail_66 ;
    wire \tok.A_stk.tail_50 ;
    wire \tok.A_stk.tail_44 ;
    wire \tok.A_stk.tail_28 ;
    wire \tok.A_stk.tail_12 ;
    wire \tok.A_12 ;
    wire \tok.A_stk.tail_8 ;
    wire \tok.A_stk.tail_24 ;
    wire \tok.A_stk.tail_56 ;
    wire \tok.A_stk.tail_40 ;
    wire \tok.n22 ;
    wire \tok.n24 ;
    wire \tok.n21 ;
    wire \tok.n30_cascade_ ;
    wire \tok.n15_adj_671 ;
    wire \tok.A_low_6 ;
    wire \tok.n18 ;
    wire \tok.n17_adj_661_cascade_ ;
    wire \tok.n19 ;
    wire \tok.n29 ;
    wire \tok.A_low_2 ;
    wire \tok.n22_adj_698 ;
    wire \tok.n24_adj_703 ;
    wire \tok.n4_adj_699_cascade_ ;
    wire \tok.n9_adj_705 ;
    wire uart_rx_data_1;
    wire \tok.n14_adj_662 ;
    wire \tok.n6_adj_834 ;
    wire \tok.n23_adj_718 ;
    wire \tok.n5_adj_835_cascade_ ;
    wire \tok.n14_adj_644 ;
    wire \tok.n10_adj_836 ;
    wire A_low_7;
    wire \tok.n6_adj_650 ;
    wire \tok.T_7 ;
    wire \tok.n11_adj_706 ;
    wire uart_rx_data_2;
    wire \tok.n12_adj_832 ;
    wire \tok.n6_adj_839_cascade_ ;
    wire \tok.n11_adj_681 ;
    wire \tok.n32 ;
    wire \tok.n15_adj_655 ;
    wire \tok.A_13 ;
    wire \tok.n211 ;
    wire \tok.n184 ;
    wire capture_5;
    wire capture_8;
    wire n4858;
    wire capture_7;
    wire \tok.n17_adj_711 ;
    wire \tok.S_0 ;
    wire \tok.n11_adj_809 ;
    wire bfn_11_9_0_;
    wire \tok.n301 ;
    wire \tok.S_1 ;
    wire \tok.n20_adj_799 ;
    wire \tok.n4769 ;
    wire \tok.S_2 ;
    wire \tok.n300 ;
    wire \tok.n22_adj_797 ;
    wire \tok.n4770 ;
    wire \tok.n10_adj_791 ;
    wire \tok.n4771 ;
    wire \tok.S_4 ;
    wire \tok.n6_adj_762 ;
    wire \tok.n4772 ;
    wire \tok.n4773 ;
    wire \tok.S_6 ;
    wire \tok.n296 ;
    wire \tok.n6 ;
    wire \tok.n4774 ;
    wire \tok.S_7 ;
    wire \tok.n295 ;
    wire \tok.n6_adj_657 ;
    wire \tok.n4775 ;
    wire \tok.n4776 ;
    wire bfn_11_10_0_;
    wire \tok.n293 ;
    wire \tok.n28 ;
    wire \tok.n4777 ;
    wire \tok.n8_adj_792 ;
    wire \tok.n292 ;
    wire \tok.n27_adj_704 ;
    wire \tok.n4778 ;
    wire \tok.n291 ;
    wire \tok.n6_adj_728 ;
    wire \tok.n4779 ;
    wire \tok.n290 ;
    wire \tok.S_12 ;
    wire \tok.n6_adj_742 ;
    wire \tok.n4780 ;
    wire \tok.n289 ;
    wire \tok.S_13 ;
    wire \tok.n6_adj_752 ;
    wire \tok.n4781 ;
    wire \tok.n4782 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \tok.n4783 ;
    wire \tok.n4783_THRU_CRY_0_THRU_CO ;
    wire \tok.n400 ;
    wire bfn_11_11_0_;
    wire \tok.n6_adj_783 ;
    wire \tok.n287 ;
    wire \tok.A_15 ;
    wire \tok.S_15 ;
    wire \tok.A_stk.tail_15 ;
    wire \tok.A_stk.tail_31 ;
    wire \tok.A_stk.tail_47 ;
    wire \tok.A_stk.tail_95 ;
    wire \tok.A_stk.tail_63 ;
    wire \tok.A_stk.tail_79 ;
    wire \tok.A_stk.tail_74 ;
    wire \tok.A_stk.tail_58 ;
    wire \tok.A_stk.tail_42 ;
    wire \tok.A_stk.tail_26 ;
    wire \tok.A_stk.tail_10 ;
    wire tail_117;
    wire tail_101;
    wire \tok.A_stk.tail_85 ;
    wire \tok.A_stk.tail_69 ;
    wire \tok.A_stk.tail_53 ;
    wire \tok.A_stk.tail_37 ;
    wire \tok.A_stk.tail_21 ;
    wire \tok.A_stk.tail_90 ;
    wire tail_122;
    wire tail_106;
    wire \tok.n23_adj_642 ;
    wire \tok.n288 ;
    wire \tok.A_11 ;
    wire \tok.A_stk.tail_14 ;
    wire \tok.S_11 ;
    wire \tok.A_stk.tail_11 ;
    wire \tok.A_stk.tail_27 ;
    wire \tok.A_stk.tail_43 ;
    wire \tok.A_stk.tail_75 ;
    wire \tok.A_stk.tail_59 ;
    wire \tok.n20_adj_648 ;
    wire \tok.n299 ;
    wire \tok.n238 ;
    wire \tok.A_stk.tail_5 ;
    wire \tok.S_3 ;
    wire \tok.A_stk.tail_3 ;
    wire \tok.A_stk.tail_19 ;
    wire \tok.A_stk.tail_35 ;
    wire \tok.A_stk.tail_67 ;
    wire A_stk_delta_1;
    wire \tok.A_stk.tail_51 ;
    wire rd_15__N_301;
    wire \tok.n175 ;
    wire \tok.n15_adj_770 ;
    wire \tok.n14_adj_769 ;
    wire \tok.n13_adj_772_cascade_ ;
    wire \tok.n5412 ;
    wire \tok.n22_adj_773_cascade_ ;
    wire \tok.A_14 ;
    wire rx_data_7__N_511;
    wire capture_6;
    wire \tok.S_5 ;
    wire uart_rx_data_5;
    wire \tok.n6_adj_717 ;
    wire \tok.table_rd_5 ;
    wire \tok.n16_adj_855 ;
    wire \tok.n5_adj_800 ;
    wire \tok.n10_adj_823 ;
    wire \tok.n20_adj_857_cascade_ ;
    wire \tok.n14_adj_856 ;
    wire \tok.n5559 ;
    wire \tok.n3_adj_859 ;
    wire \tok.n22_adj_861_cascade_ ;
    wire \tok.n18_adj_860 ;
    wire \tok.n5556 ;
    wire \tok.n15 ;
    wire \tok.n5_adj_669 ;
    wire \tok.table_rd_8 ;
    wire \tok.n4908 ;
    wire \tok.n181 ;
    wire \tok.n2735 ;
    wire \tok.n15_adj_670 ;
    wire \tok.n13_adj_674_cascade_ ;
    wire \tok.n5416 ;
    wire \tok.n23 ;
    wire \tok.n22_adj_676_cascade_ ;
    wire clk;
    wire \tok.n995 ;
    wire \tok.reset_N_2 ;
    wire \tok.S_8 ;
    wire \tok.n5544 ;
    wire \tok.n5542 ;
    wire \tok.n10_adj_666 ;
    wire \tok.n15_adj_667 ;
    wire \tok.n14_adj_668 ;
    wire \tok.n880 ;
    wire \tok.A_low_0 ;
    wire \tok.n904 ;
    wire \tok.n5372 ;
    wire \tok.S_9 ;
    wire \tok.n8_adj_689 ;
    wire \tok.S_10 ;
    wire \tok.n8_adj_702 ;
    wire \tok.n298 ;
    wire \tok.A_low_5 ;
    wire \tok.n297 ;
    wire \tok.T_2 ;
    wire \tok.n5366 ;
    wire \tok.A_low_3 ;
    wire \tok.A_low_4 ;
    wire \tok.n5396_cascade_ ;
    wire \tok.n18_adj_677 ;
    wire \tok.A_8 ;
    wire \tok.n294 ;
    wire \tok.n191 ;
    wire \tok.A_10 ;
    wire \tok.n2703 ;
    wire \tok.A_9 ;
    wire \tok.n202_cascade_ ;
    wire \tok.n2743 ;
    wire \tok.n5520 ;
    wire \tok.S_14 ;
    wire \tok.n18_adj_774_cascade_ ;
    wire \tok.n2661 ;
    wire \tok.n5518 ;
    wire _gnd_net_;

    defparam \tok.vals.mem1_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .WRITE_MODE=0;
    defparam \tok.vals.mem1_physical .READ_MODE=0;
    defparam \tok.vals.mem1_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \tok.vals.mem1_physical  (
            .RDATA({\tok.table_rd_15 ,\tok.table_rd_14 ,\tok.table_rd_13 ,\tok.table_rd_12 ,\tok.table_rd_11 ,\tok.table_rd_10 ,\tok.table_rd_9 ,\tok.table_rd_8 ,\tok.table_rd_7 ,\tok.table_rd_6 ,\tok.table_rd_5 ,\tok.table_rd_4 ,\tok.table_rd_3 ,\tok.table_rd_2 ,\tok.table_rd_1 ,\tok.table_rd_0 }),
            .RADDR({dangling_wire_0,dangling_wire_1,dangling_wire_2,N__14563,N__14638,N__14719,N__14794,N__16786,N__16996,N__16654,N__14872}),
            .WADDR({dangling_wire_3,dangling_wire_4,dangling_wire_5,N__14560,N__14635,N__14710,N__14785,N__16795,N__16993,N__16645,N__14863}),
            .MASK({dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .WDATA({N__12224,N__12212,N__12152,N__12143,N__12266,N__12257,N__12251,N__12245,N__12161,N__15290,N__12170,N__12065,N__12206,N__12194,N__12179,N__12239}),
            .RCLKE(),
            .RCLK(N__28504),
            .RE(N__24254),
            .WCLKE(),
            .WCLK(N__28503),
            .WE(N__15164));
    defparam \tok.keys.mem0_physical .WRITE_MODE=0;
    defparam \tok.keys.mem0_physical .READ_MODE=0;
    defparam \tok.keys.mem0_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \tok.keys.mem0_physical  (
            .RDATA({\tok.key_rd_15 ,\tok.key_rd_14 ,\tok.key_rd_13 ,\tok.key_rd_12 ,\tok.key_rd_11 ,\tok.key_rd_10 ,\tok.key_rd_9 ,\tok.key_rd_8 ,\tok.key_rd_7 ,\tok.key_rd_6 ,\tok.key_rd_5 ,\tok.key_rd_4 ,\tok.key_rd_3 ,\tok.key_rd_2 ,\tok.key_rd_1 ,\tok.key_rd_0 }),
            .RADDR({dangling_wire_22,dangling_wire_23,dangling_wire_24,N__14573,N__14648,N__14726,N__14801,N__16798,N__17006,N__16661,N__14879}),
            .WADDR({dangling_wire_25,dangling_wire_26,dangling_wire_27,N__14572,N__14647,N__14722,N__14797,N__16802,N__17005,N__16657,N__14875}),
            .MASK({dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .WDATA({N__24863,N__25766,N__23156,N__21633,N__25160,N__29268,N__29080,N__29471,N__22327,N__21895,N__27326,N__29609,N__29730,N__22766,N__21141,N__27780}),
            .RCLKE(),
            .RCLK(N__28490),
            .RE(N__24260),
            .WCLKE(),
            .WCLK(N__28491),
            .WE(N__15163));
    defparam \tok.ram.mem2_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101000100000100000001000001010101000101;
    defparam \tok.ram.mem2_physical .WRITE_MODE=1;
    defparam \tok.ram.mem2_physical .READ_MODE=1;
    defparam \tok.ram.mem2_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \tok.ram.mem2_physical  (
            .RDATA({dangling_wire_44,\tok.T_7 ,dangling_wire_45,\tok.T_6 ,dangling_wire_46,\tok.T_5 ,dangling_wire_47,\tok.T_4 ,dangling_wire_48,\tok.T_3 ,dangling_wire_49,\tok.T_2 ,dangling_wire_50,\tok.T_1 ,dangling_wire_51,\tok.T_0 }),
            .RADDR({dangling_wire_52,dangling_wire_53,dangling_wire_54,N__11597,N__12524,N__12086,N__16220,N__11366,N__11342,N__15695,N__11390}),
            .WADDR({dangling_wire_55,dangling_wire_56,dangling_wire_57,N__23558,N__23678,N__27221,N__23795,N__25379,N__23939,N__24050,N__22879}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,N__22328,dangling_wire_75,N__21896,dangling_wire_76,N__27352,dangling_wire_77,N__29600,dangling_wire_78,N__29729,dangling_wire_79,N__22765,dangling_wire_80,N__21140,dangling_wire_81,N__27781}),
            .RCLKE(),
            .RCLK(N__28515),
            .RE(N__24247),
            .WCLKE(),
            .WCLK(N__28516),
            .WE(N__20764));
    defparam rx_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_pad_iopad.PULLUP=1'b0;
    IO_PAD rx_pad_iopad (
            .OE(N__30069),
            .DIN(N__30068),
            .DOUT(N__30067),
            .PACKAGEPIN(rx));
    defparam rx_pad_preio.PIN_TYPE=6'b000001;
    defparam rx_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_pad_preio (
            .PADOEN(N__30069),
            .PADOUT(N__30068),
            .PADIN(N__30067),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(rx_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam tx_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_pad_iopad.PULLUP=1'b0;
    IO_PAD tx_pad_iopad (
            .OE(N__30060),
            .DIN(N__30059),
            .DOUT(N__30058),
            .PACKAGEPIN(tx));
    defparam tx_pad_preio.PIN_TYPE=6'b011001;
    defparam tx_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_pad_preio (
            .PADOEN(N__30060),
            .PADOUT(N__30059),
            .PADIN(N__30058),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11621),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam reset_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam reset_pad_iopad.PULLUP=1'b0;
    IO_PAD reset_pad_iopad (
            .OE(N__30051),
            .DIN(N__30050),
            .DOUT(N__30049),
            .PACKAGEPIN(reset));
    defparam reset_pad_preio.PIN_TYPE=6'b000001;
    defparam reset_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO reset_pad_preio (
            .PADOEN(N__30051),
            .PADOUT(N__30050),
            .PADIN(N__30049),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(reset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__7478 (
            .O(N__30032),
            .I(N__30022));
    InMux I__7477 (
            .O(N__30031),
            .I(N__30008));
    InMux I__7476 (
            .O(N__30030),
            .I(N__30008));
    InMux I__7475 (
            .O(N__30029),
            .I(N__30003));
    InMux I__7474 (
            .O(N__30028),
            .I(N__30003));
    InMux I__7473 (
            .O(N__30027),
            .I(N__29998));
    InMux I__7472 (
            .O(N__30026),
            .I(N__29998));
    InMux I__7471 (
            .O(N__30025),
            .I(N__29990));
    LocalMux I__7470 (
            .O(N__30022),
            .I(N__29987));
    InMux I__7469 (
            .O(N__30021),
            .I(N__29981));
    InMux I__7468 (
            .O(N__30020),
            .I(N__29978));
    InMux I__7467 (
            .O(N__30019),
            .I(N__29973));
    InMux I__7466 (
            .O(N__30018),
            .I(N__29973));
    InMux I__7465 (
            .O(N__30017),
            .I(N__29970));
    CascadeMux I__7464 (
            .O(N__30016),
            .I(N__29966));
    CascadeMux I__7463 (
            .O(N__30015),
            .I(N__29963));
    CascadeMux I__7462 (
            .O(N__30014),
            .I(N__29959));
    InMux I__7461 (
            .O(N__30013),
            .I(N__29955));
    LocalMux I__7460 (
            .O(N__30008),
            .I(N__29948));
    LocalMux I__7459 (
            .O(N__30003),
            .I(N__29948));
    LocalMux I__7458 (
            .O(N__29998),
            .I(N__29948));
    InMux I__7457 (
            .O(N__29997),
            .I(N__29931));
    InMux I__7456 (
            .O(N__29996),
            .I(N__29931));
    InMux I__7455 (
            .O(N__29995),
            .I(N__29931));
    InMux I__7454 (
            .O(N__29994),
            .I(N__29931));
    InMux I__7453 (
            .O(N__29993),
            .I(N__29931));
    LocalMux I__7452 (
            .O(N__29990),
            .I(N__29928));
    Span4Mux_v I__7451 (
            .O(N__29987),
            .I(N__29924));
    InMux I__7450 (
            .O(N__29986),
            .I(N__29919));
    InMux I__7449 (
            .O(N__29985),
            .I(N__29919));
    InMux I__7448 (
            .O(N__29984),
            .I(N__29916));
    LocalMux I__7447 (
            .O(N__29981),
            .I(N__29901));
    LocalMux I__7446 (
            .O(N__29978),
            .I(N__29901));
    LocalMux I__7445 (
            .O(N__29973),
            .I(N__29901));
    LocalMux I__7444 (
            .O(N__29970),
            .I(N__29901));
    InMux I__7443 (
            .O(N__29969),
            .I(N__29890));
    InMux I__7442 (
            .O(N__29966),
            .I(N__29890));
    InMux I__7441 (
            .O(N__29963),
            .I(N__29890));
    InMux I__7440 (
            .O(N__29962),
            .I(N__29890));
    InMux I__7439 (
            .O(N__29959),
            .I(N__29890));
    InMux I__7438 (
            .O(N__29958),
            .I(N__29887));
    LocalMux I__7437 (
            .O(N__29955),
            .I(N__29882));
    Span4Mux_v I__7436 (
            .O(N__29948),
            .I(N__29882));
    InMux I__7435 (
            .O(N__29947),
            .I(N__29879));
    InMux I__7434 (
            .O(N__29946),
            .I(N__29873));
    InMux I__7433 (
            .O(N__29945),
            .I(N__29873));
    InMux I__7432 (
            .O(N__29944),
            .I(N__29866));
    InMux I__7431 (
            .O(N__29943),
            .I(N__29866));
    InMux I__7430 (
            .O(N__29942),
            .I(N__29866));
    LocalMux I__7429 (
            .O(N__29931),
            .I(N__29861));
    Span4Mux_h I__7428 (
            .O(N__29928),
            .I(N__29861));
    CascadeMux I__7427 (
            .O(N__29927),
            .I(N__29847));
    Span4Mux_h I__7426 (
            .O(N__29924),
            .I(N__29844));
    LocalMux I__7425 (
            .O(N__29919),
            .I(N__29839));
    LocalMux I__7424 (
            .O(N__29916),
            .I(N__29839));
    InMux I__7423 (
            .O(N__29915),
            .I(N__29826));
    InMux I__7422 (
            .O(N__29914),
            .I(N__29826));
    InMux I__7421 (
            .O(N__29913),
            .I(N__29826));
    InMux I__7420 (
            .O(N__29912),
            .I(N__29826));
    InMux I__7419 (
            .O(N__29911),
            .I(N__29826));
    InMux I__7418 (
            .O(N__29910),
            .I(N__29826));
    Span4Mux_s3_v I__7417 (
            .O(N__29901),
            .I(N__29819));
    LocalMux I__7416 (
            .O(N__29890),
            .I(N__29819));
    LocalMux I__7415 (
            .O(N__29887),
            .I(N__29819));
    Span4Mux_v I__7414 (
            .O(N__29882),
            .I(N__29816));
    LocalMux I__7413 (
            .O(N__29879),
            .I(N__29813));
    InMux I__7412 (
            .O(N__29878),
            .I(N__29810));
    LocalMux I__7411 (
            .O(N__29873),
            .I(N__29803));
    LocalMux I__7410 (
            .O(N__29866),
            .I(N__29803));
    Span4Mux_v I__7409 (
            .O(N__29861),
            .I(N__29803));
    InMux I__7408 (
            .O(N__29860),
            .I(N__29790));
    InMux I__7407 (
            .O(N__29859),
            .I(N__29790));
    InMux I__7406 (
            .O(N__29858),
            .I(N__29790));
    InMux I__7405 (
            .O(N__29857),
            .I(N__29790));
    InMux I__7404 (
            .O(N__29856),
            .I(N__29790));
    InMux I__7403 (
            .O(N__29855),
            .I(N__29790));
    InMux I__7402 (
            .O(N__29854),
            .I(N__29777));
    InMux I__7401 (
            .O(N__29853),
            .I(N__29777));
    InMux I__7400 (
            .O(N__29852),
            .I(N__29777));
    InMux I__7399 (
            .O(N__29851),
            .I(N__29777));
    InMux I__7398 (
            .O(N__29850),
            .I(N__29777));
    InMux I__7397 (
            .O(N__29847),
            .I(N__29777));
    Span4Mux_h I__7396 (
            .O(N__29844),
            .I(N__29770));
    Span4Mux_v I__7395 (
            .O(N__29839),
            .I(N__29770));
    LocalMux I__7394 (
            .O(N__29826),
            .I(N__29770));
    Span4Mux_h I__7393 (
            .O(N__29819),
            .I(N__29767));
    Odrv4 I__7392 (
            .O(N__29816),
            .I(\tok.T_2 ));
    Odrv4 I__7391 (
            .O(N__29813),
            .I(\tok.T_2 ));
    LocalMux I__7390 (
            .O(N__29810),
            .I(\tok.T_2 ));
    Odrv4 I__7389 (
            .O(N__29803),
            .I(\tok.T_2 ));
    LocalMux I__7388 (
            .O(N__29790),
            .I(\tok.T_2 ));
    LocalMux I__7387 (
            .O(N__29777),
            .I(\tok.T_2 ));
    Odrv4 I__7386 (
            .O(N__29770),
            .I(\tok.T_2 ));
    Odrv4 I__7385 (
            .O(N__29767),
            .I(\tok.T_2 ));
    InMux I__7384 (
            .O(N__29750),
            .I(N__29747));
    LocalMux I__7383 (
            .O(N__29747),
            .I(N__29744));
    Span4Mux_v I__7382 (
            .O(N__29744),
            .I(N__29741));
    Odrv4 I__7381 (
            .O(N__29741),
            .I(\tok.n5366 ));
    CascadeMux I__7380 (
            .O(N__29738),
            .I(N__29735));
    InMux I__7379 (
            .O(N__29735),
            .I(N__29725));
    InMux I__7378 (
            .O(N__29734),
            .I(N__29717));
    InMux I__7377 (
            .O(N__29733),
            .I(N__29717));
    InMux I__7376 (
            .O(N__29732),
            .I(N__29717));
    InMux I__7375 (
            .O(N__29731),
            .I(N__29714));
    InMux I__7374 (
            .O(N__29730),
            .I(N__29711));
    InMux I__7373 (
            .O(N__29729),
            .I(N__29708));
    InMux I__7372 (
            .O(N__29728),
            .I(N__29705));
    LocalMux I__7371 (
            .O(N__29725),
            .I(N__29697));
    InMux I__7370 (
            .O(N__29724),
            .I(N__29694));
    LocalMux I__7369 (
            .O(N__29717),
            .I(N__29691));
    LocalMux I__7368 (
            .O(N__29714),
            .I(N__29688));
    LocalMux I__7367 (
            .O(N__29711),
            .I(N__29684));
    LocalMux I__7366 (
            .O(N__29708),
            .I(N__29681));
    LocalMux I__7365 (
            .O(N__29705),
            .I(N__29678));
    InMux I__7364 (
            .O(N__29704),
            .I(N__29675));
    InMux I__7363 (
            .O(N__29703),
            .I(N__29672));
    InMux I__7362 (
            .O(N__29702),
            .I(N__29669));
    InMux I__7361 (
            .O(N__29701),
            .I(N__29666));
    InMux I__7360 (
            .O(N__29700),
            .I(N__29663));
    Span4Mux_v I__7359 (
            .O(N__29697),
            .I(N__29658));
    LocalMux I__7358 (
            .O(N__29694),
            .I(N__29658));
    Span4Mux_s2_h I__7357 (
            .O(N__29691),
            .I(N__29655));
    Span4Mux_v I__7356 (
            .O(N__29688),
            .I(N__29652));
    InMux I__7355 (
            .O(N__29687),
            .I(N__29649));
    Span4Mux_h I__7354 (
            .O(N__29684),
            .I(N__29642));
    Span4Mux_h I__7353 (
            .O(N__29681),
            .I(N__29642));
    Span4Mux_h I__7352 (
            .O(N__29678),
            .I(N__29642));
    LocalMux I__7351 (
            .O(N__29675),
            .I(N__29637));
    LocalMux I__7350 (
            .O(N__29672),
            .I(N__29637));
    LocalMux I__7349 (
            .O(N__29669),
            .I(N__29632));
    LocalMux I__7348 (
            .O(N__29666),
            .I(N__29632));
    LocalMux I__7347 (
            .O(N__29663),
            .I(N__29629));
    Span4Mux_h I__7346 (
            .O(N__29658),
            .I(N__29624));
    Span4Mux_h I__7345 (
            .O(N__29655),
            .I(N__29624));
    Odrv4 I__7344 (
            .O(N__29652),
            .I(\tok.A_low_3 ));
    LocalMux I__7343 (
            .O(N__29649),
            .I(\tok.A_low_3 ));
    Odrv4 I__7342 (
            .O(N__29642),
            .I(\tok.A_low_3 ));
    Odrv12 I__7341 (
            .O(N__29637),
            .I(\tok.A_low_3 ));
    Odrv4 I__7340 (
            .O(N__29632),
            .I(\tok.A_low_3 ));
    Odrv4 I__7339 (
            .O(N__29629),
            .I(\tok.A_low_3 ));
    Odrv4 I__7338 (
            .O(N__29624),
            .I(\tok.A_low_3 ));
    InMux I__7337 (
            .O(N__29609),
            .I(N__29604));
    CascadeMux I__7336 (
            .O(N__29608),
            .I(N__29601));
    InMux I__7335 (
            .O(N__29607),
            .I(N__29593));
    LocalMux I__7334 (
            .O(N__29604),
            .I(N__29590));
    InMux I__7333 (
            .O(N__29601),
            .I(N__29587));
    InMux I__7332 (
            .O(N__29600),
            .I(N__29582));
    InMux I__7331 (
            .O(N__29599),
            .I(N__29579));
    InMux I__7330 (
            .O(N__29598),
            .I(N__29576));
    InMux I__7329 (
            .O(N__29597),
            .I(N__29573));
    InMux I__7328 (
            .O(N__29596),
            .I(N__29570));
    LocalMux I__7327 (
            .O(N__29593),
            .I(N__29567));
    Span4Mux_h I__7326 (
            .O(N__29590),
            .I(N__29559));
    LocalMux I__7325 (
            .O(N__29587),
            .I(N__29559));
    InMux I__7324 (
            .O(N__29586),
            .I(N__29556));
    InMux I__7323 (
            .O(N__29585),
            .I(N__29553));
    LocalMux I__7322 (
            .O(N__29582),
            .I(N__29549));
    LocalMux I__7321 (
            .O(N__29579),
            .I(N__29546));
    LocalMux I__7320 (
            .O(N__29576),
            .I(N__29540));
    LocalMux I__7319 (
            .O(N__29573),
            .I(N__29540));
    LocalMux I__7318 (
            .O(N__29570),
            .I(N__29537));
    Sp12to4 I__7317 (
            .O(N__29567),
            .I(N__29534));
    InMux I__7316 (
            .O(N__29566),
            .I(N__29527));
    InMux I__7315 (
            .O(N__29565),
            .I(N__29527));
    InMux I__7314 (
            .O(N__29564),
            .I(N__29527));
    Span4Mux_h I__7313 (
            .O(N__29559),
            .I(N__29520));
    LocalMux I__7312 (
            .O(N__29556),
            .I(N__29520));
    LocalMux I__7311 (
            .O(N__29553),
            .I(N__29520));
    InMux I__7310 (
            .O(N__29552),
            .I(N__29517));
    Span4Mux_h I__7309 (
            .O(N__29549),
            .I(N__29514));
    Span12Mux_s9_v I__7308 (
            .O(N__29546),
            .I(N__29511));
    InMux I__7307 (
            .O(N__29545),
            .I(N__29508));
    Span4Mux_h I__7306 (
            .O(N__29540),
            .I(N__29505));
    Span12Mux_s4_v I__7305 (
            .O(N__29537),
            .I(N__29498));
    Span12Mux_s9_v I__7304 (
            .O(N__29534),
            .I(N__29498));
    LocalMux I__7303 (
            .O(N__29527),
            .I(N__29498));
    Span4Mux_v I__7302 (
            .O(N__29520),
            .I(N__29493));
    LocalMux I__7301 (
            .O(N__29517),
            .I(N__29493));
    Odrv4 I__7300 (
            .O(N__29514),
            .I(\tok.A_low_4 ));
    Odrv12 I__7299 (
            .O(N__29511),
            .I(\tok.A_low_4 ));
    LocalMux I__7298 (
            .O(N__29508),
            .I(\tok.A_low_4 ));
    Odrv4 I__7297 (
            .O(N__29505),
            .I(\tok.A_low_4 ));
    Odrv12 I__7296 (
            .O(N__29498),
            .I(\tok.A_low_4 ));
    Odrv4 I__7295 (
            .O(N__29493),
            .I(\tok.A_low_4 ));
    CascadeMux I__7294 (
            .O(N__29480),
            .I(\tok.n5396_cascade_ ));
    InMux I__7293 (
            .O(N__29477),
            .I(N__29474));
    LocalMux I__7292 (
            .O(N__29474),
            .I(\tok.n18_adj_677 ));
    InMux I__7291 (
            .O(N__29471),
            .I(N__29465));
    CascadeMux I__7290 (
            .O(N__29470),
            .I(N__29461));
    InMux I__7289 (
            .O(N__29469),
            .I(N__29456));
    InMux I__7288 (
            .O(N__29468),
            .I(N__29453));
    LocalMux I__7287 (
            .O(N__29465),
            .I(N__29449));
    InMux I__7286 (
            .O(N__29464),
            .I(N__29442));
    InMux I__7285 (
            .O(N__29461),
            .I(N__29442));
    InMux I__7284 (
            .O(N__29460),
            .I(N__29438));
    InMux I__7283 (
            .O(N__29459),
            .I(N__29435));
    LocalMux I__7282 (
            .O(N__29456),
            .I(N__29430));
    LocalMux I__7281 (
            .O(N__29453),
            .I(N__29430));
    InMux I__7280 (
            .O(N__29452),
            .I(N__29427));
    Span4Mux_v I__7279 (
            .O(N__29449),
            .I(N__29424));
    InMux I__7278 (
            .O(N__29448),
            .I(N__29421));
    InMux I__7277 (
            .O(N__29447),
            .I(N__29418));
    LocalMux I__7276 (
            .O(N__29442),
            .I(N__29415));
    CascadeMux I__7275 (
            .O(N__29441),
            .I(N__29412));
    LocalMux I__7274 (
            .O(N__29438),
            .I(N__29408));
    LocalMux I__7273 (
            .O(N__29435),
            .I(N__29402));
    Span4Mux_h I__7272 (
            .O(N__29430),
            .I(N__29402));
    LocalMux I__7271 (
            .O(N__29427),
            .I(N__29399));
    Span4Mux_h I__7270 (
            .O(N__29424),
            .I(N__29390));
    LocalMux I__7269 (
            .O(N__29421),
            .I(N__29390));
    LocalMux I__7268 (
            .O(N__29418),
            .I(N__29390));
    Span4Mux_v I__7267 (
            .O(N__29415),
            .I(N__29390));
    InMux I__7266 (
            .O(N__29412),
            .I(N__29385));
    InMux I__7265 (
            .O(N__29411),
            .I(N__29385));
    Span4Mux_v I__7264 (
            .O(N__29408),
            .I(N__29382));
    InMux I__7263 (
            .O(N__29407),
            .I(N__29379));
    Span4Mux_h I__7262 (
            .O(N__29402),
            .I(N__29376));
    Span4Mux_v I__7261 (
            .O(N__29399),
            .I(N__29371));
    Span4Mux_h I__7260 (
            .O(N__29390),
            .I(N__29371));
    LocalMux I__7259 (
            .O(N__29385),
            .I(\tok.A_8 ));
    Odrv4 I__7258 (
            .O(N__29382),
            .I(\tok.A_8 ));
    LocalMux I__7257 (
            .O(N__29379),
            .I(\tok.A_8 ));
    Odrv4 I__7256 (
            .O(N__29376),
            .I(\tok.A_8 ));
    Odrv4 I__7255 (
            .O(N__29371),
            .I(\tok.A_8 ));
    InMux I__7254 (
            .O(N__29360),
            .I(N__29357));
    LocalMux I__7253 (
            .O(N__29357),
            .I(\tok.n294 ));
    InMux I__7252 (
            .O(N__29354),
            .I(N__29350));
    InMux I__7251 (
            .O(N__29353),
            .I(N__29346));
    LocalMux I__7250 (
            .O(N__29350),
            .I(N__29340));
    InMux I__7249 (
            .O(N__29349),
            .I(N__29337));
    LocalMux I__7248 (
            .O(N__29346),
            .I(N__29334));
    InMux I__7247 (
            .O(N__29345),
            .I(N__29329));
    InMux I__7246 (
            .O(N__29344),
            .I(N__29329));
    InMux I__7245 (
            .O(N__29343),
            .I(N__29326));
    Span4Mux_v I__7244 (
            .O(N__29340),
            .I(N__29323));
    LocalMux I__7243 (
            .O(N__29337),
            .I(N__29320));
    Span4Mux_s2_h I__7242 (
            .O(N__29334),
            .I(N__29314));
    LocalMux I__7241 (
            .O(N__29329),
            .I(N__29314));
    LocalMux I__7240 (
            .O(N__29326),
            .I(N__29311));
    Span4Mux_h I__7239 (
            .O(N__29323),
            .I(N__29305));
    Span4Mux_v I__7238 (
            .O(N__29320),
            .I(N__29305));
    InMux I__7237 (
            .O(N__29319),
            .I(N__29302));
    Span4Mux_h I__7236 (
            .O(N__29314),
            .I(N__29299));
    Span4Mux_h I__7235 (
            .O(N__29311),
            .I(N__29296));
    InMux I__7234 (
            .O(N__29310),
            .I(N__29293));
    Odrv4 I__7233 (
            .O(N__29305),
            .I(\tok.n191 ));
    LocalMux I__7232 (
            .O(N__29302),
            .I(\tok.n191 ));
    Odrv4 I__7231 (
            .O(N__29299),
            .I(\tok.n191 ));
    Odrv4 I__7230 (
            .O(N__29296),
            .I(\tok.n191 ));
    LocalMux I__7229 (
            .O(N__29293),
            .I(\tok.n191 ));
    InMux I__7228 (
            .O(N__29282),
            .I(N__29279));
    LocalMux I__7227 (
            .O(N__29279),
            .I(N__29275));
    InMux I__7226 (
            .O(N__29278),
            .I(N__29272));
    Span4Mux_s3_v I__7225 (
            .O(N__29275),
            .I(N__29263));
    LocalMux I__7224 (
            .O(N__29272),
            .I(N__29260));
    InMux I__7223 (
            .O(N__29271),
            .I(N__29257));
    InMux I__7222 (
            .O(N__29270),
            .I(N__29254));
    InMux I__7221 (
            .O(N__29269),
            .I(N__29250));
    InMux I__7220 (
            .O(N__29268),
            .I(N__29246));
    InMux I__7219 (
            .O(N__29267),
            .I(N__29241));
    InMux I__7218 (
            .O(N__29266),
            .I(N__29241));
    Span4Mux_v I__7217 (
            .O(N__29263),
            .I(N__29233));
    Span4Mux_v I__7216 (
            .O(N__29260),
            .I(N__29233));
    LocalMux I__7215 (
            .O(N__29257),
            .I(N__29233));
    LocalMux I__7214 (
            .O(N__29254),
            .I(N__29230));
    InMux I__7213 (
            .O(N__29253),
            .I(N__29227));
    LocalMux I__7212 (
            .O(N__29250),
            .I(N__29224));
    InMux I__7211 (
            .O(N__29249),
            .I(N__29221));
    LocalMux I__7210 (
            .O(N__29246),
            .I(N__29216));
    LocalMux I__7209 (
            .O(N__29241),
            .I(N__29216));
    InMux I__7208 (
            .O(N__29240),
            .I(N__29212));
    Span4Mux_h I__7207 (
            .O(N__29233),
            .I(N__29209));
    Span4Mux_v I__7206 (
            .O(N__29230),
            .I(N__29204));
    LocalMux I__7205 (
            .O(N__29227),
            .I(N__29204));
    Span4Mux_h I__7204 (
            .O(N__29224),
            .I(N__29199));
    LocalMux I__7203 (
            .O(N__29221),
            .I(N__29199));
    Span4Mux_h I__7202 (
            .O(N__29216),
            .I(N__29196));
    InMux I__7201 (
            .O(N__29215),
            .I(N__29193));
    LocalMux I__7200 (
            .O(N__29212),
            .I(\tok.A_10 ));
    Odrv4 I__7199 (
            .O(N__29209),
            .I(\tok.A_10 ));
    Odrv4 I__7198 (
            .O(N__29204),
            .I(\tok.A_10 ));
    Odrv4 I__7197 (
            .O(N__29199),
            .I(\tok.A_10 ));
    Odrv4 I__7196 (
            .O(N__29196),
            .I(\tok.A_10 ));
    LocalMux I__7195 (
            .O(N__29193),
            .I(\tok.A_10 ));
    InMux I__7194 (
            .O(N__29180),
            .I(N__29175));
    InMux I__7193 (
            .O(N__29179),
            .I(N__29172));
    InMux I__7192 (
            .O(N__29178),
            .I(N__29168));
    LocalMux I__7191 (
            .O(N__29175),
            .I(N__29164));
    LocalMux I__7190 (
            .O(N__29172),
            .I(N__29161));
    InMux I__7189 (
            .O(N__29171),
            .I(N__29157));
    LocalMux I__7188 (
            .O(N__29168),
            .I(N__29154));
    InMux I__7187 (
            .O(N__29167),
            .I(N__29150));
    Span4Mux_s1_h I__7186 (
            .O(N__29164),
            .I(N__29143));
    Span4Mux_v I__7185 (
            .O(N__29161),
            .I(N__29143));
    InMux I__7184 (
            .O(N__29160),
            .I(N__29140));
    LocalMux I__7183 (
            .O(N__29157),
            .I(N__29135));
    Span4Mux_s3_h I__7182 (
            .O(N__29154),
            .I(N__29132));
    InMux I__7181 (
            .O(N__29153),
            .I(N__29129));
    LocalMux I__7180 (
            .O(N__29150),
            .I(N__29126));
    InMux I__7179 (
            .O(N__29149),
            .I(N__29123));
    InMux I__7178 (
            .O(N__29148),
            .I(N__29120));
    Span4Mux_h I__7177 (
            .O(N__29143),
            .I(N__29114));
    LocalMux I__7176 (
            .O(N__29140),
            .I(N__29114));
    InMux I__7175 (
            .O(N__29139),
            .I(N__29109));
    InMux I__7174 (
            .O(N__29138),
            .I(N__29109));
    Span4Mux_s2_v I__7173 (
            .O(N__29135),
            .I(N__29102));
    Span4Mux_v I__7172 (
            .O(N__29132),
            .I(N__29102));
    LocalMux I__7171 (
            .O(N__29129),
            .I(N__29102));
    Sp12to4 I__7170 (
            .O(N__29126),
            .I(N__29095));
    LocalMux I__7169 (
            .O(N__29123),
            .I(N__29095));
    LocalMux I__7168 (
            .O(N__29120),
            .I(N__29095));
    InMux I__7167 (
            .O(N__29119),
            .I(N__29092));
    Odrv4 I__7166 (
            .O(N__29114),
            .I(\tok.n2703 ));
    LocalMux I__7165 (
            .O(N__29109),
            .I(\tok.n2703 ));
    Odrv4 I__7164 (
            .O(N__29102),
            .I(\tok.n2703 ));
    Odrv12 I__7163 (
            .O(N__29095),
            .I(\tok.n2703 ));
    LocalMux I__7162 (
            .O(N__29092),
            .I(\tok.n2703 ));
    InMux I__7161 (
            .O(N__29081),
            .I(N__29076));
    InMux I__7160 (
            .O(N__29080),
            .I(N__29071));
    InMux I__7159 (
            .O(N__29079),
            .I(N__29067));
    LocalMux I__7158 (
            .O(N__29076),
            .I(N__29062));
    InMux I__7157 (
            .O(N__29075),
            .I(N__29056));
    InMux I__7156 (
            .O(N__29074),
            .I(N__29056));
    LocalMux I__7155 (
            .O(N__29071),
            .I(N__29053));
    InMux I__7154 (
            .O(N__29070),
            .I(N__29050));
    LocalMux I__7153 (
            .O(N__29067),
            .I(N__29047));
    InMux I__7152 (
            .O(N__29066),
            .I(N__29044));
    CascadeMux I__7151 (
            .O(N__29065),
            .I(N__29041));
    Span4Mux_s2_v I__7150 (
            .O(N__29062),
            .I(N__29035));
    InMux I__7149 (
            .O(N__29061),
            .I(N__29032));
    LocalMux I__7148 (
            .O(N__29056),
            .I(N__29029));
    Span4Mux_h I__7147 (
            .O(N__29053),
            .I(N__29024));
    LocalMux I__7146 (
            .O(N__29050),
            .I(N__29024));
    Sp12to4 I__7145 (
            .O(N__29047),
            .I(N__29021));
    LocalMux I__7144 (
            .O(N__29044),
            .I(N__29018));
    InMux I__7143 (
            .O(N__29041),
            .I(N__29015));
    InMux I__7142 (
            .O(N__29040),
            .I(N__29012));
    InMux I__7141 (
            .O(N__29039),
            .I(N__29009));
    InMux I__7140 (
            .O(N__29038),
            .I(N__29006));
    Span4Mux_v I__7139 (
            .O(N__29035),
            .I(N__28997));
    LocalMux I__7138 (
            .O(N__29032),
            .I(N__28997));
    Span4Mux_h I__7137 (
            .O(N__29029),
            .I(N__28997));
    Span4Mux_h I__7136 (
            .O(N__29024),
            .I(N__28997));
    Odrv12 I__7135 (
            .O(N__29021),
            .I(\tok.A_9 ));
    Odrv4 I__7134 (
            .O(N__29018),
            .I(\tok.A_9 ));
    LocalMux I__7133 (
            .O(N__29015),
            .I(\tok.A_9 ));
    LocalMux I__7132 (
            .O(N__29012),
            .I(\tok.A_9 ));
    LocalMux I__7131 (
            .O(N__29009),
            .I(\tok.A_9 ));
    LocalMux I__7130 (
            .O(N__29006),
            .I(\tok.A_9 ));
    Odrv4 I__7129 (
            .O(N__28997),
            .I(\tok.A_9 ));
    CascadeMux I__7128 (
            .O(N__28982),
            .I(\tok.n202_cascade_ ));
    CascadeMux I__7127 (
            .O(N__28979),
            .I(N__28974));
    InMux I__7126 (
            .O(N__28978),
            .I(N__28967));
    InMux I__7125 (
            .O(N__28977),
            .I(N__28964));
    InMux I__7124 (
            .O(N__28974),
            .I(N__28957));
    InMux I__7123 (
            .O(N__28973),
            .I(N__28957));
    InMux I__7122 (
            .O(N__28972),
            .I(N__28957));
    InMux I__7121 (
            .O(N__28971),
            .I(N__28954));
    InMux I__7120 (
            .O(N__28970),
            .I(N__28951));
    LocalMux I__7119 (
            .O(N__28967),
            .I(N__28946));
    LocalMux I__7118 (
            .O(N__28964),
            .I(N__28943));
    LocalMux I__7117 (
            .O(N__28957),
            .I(N__28940));
    LocalMux I__7116 (
            .O(N__28954),
            .I(N__28930));
    LocalMux I__7115 (
            .O(N__28951),
            .I(N__28930));
    InMux I__7114 (
            .O(N__28950),
            .I(N__28925));
    InMux I__7113 (
            .O(N__28949),
            .I(N__28925));
    Span4Mux_v I__7112 (
            .O(N__28946),
            .I(N__28922));
    Span4Mux_v I__7111 (
            .O(N__28943),
            .I(N__28917));
    Span4Mux_v I__7110 (
            .O(N__28940),
            .I(N__28917));
    InMux I__7109 (
            .O(N__28939),
            .I(N__28914));
    InMux I__7108 (
            .O(N__28938),
            .I(N__28905));
    InMux I__7107 (
            .O(N__28937),
            .I(N__28905));
    InMux I__7106 (
            .O(N__28936),
            .I(N__28905));
    InMux I__7105 (
            .O(N__28935),
            .I(N__28905));
    Span4Mux_h I__7104 (
            .O(N__28930),
            .I(N__28901));
    LocalMux I__7103 (
            .O(N__28925),
            .I(N__28898));
    Span4Mux_v I__7102 (
            .O(N__28922),
            .I(N__28893));
    Span4Mux_h I__7101 (
            .O(N__28917),
            .I(N__28893));
    LocalMux I__7100 (
            .O(N__28914),
            .I(N__28888));
    LocalMux I__7099 (
            .O(N__28905),
            .I(N__28888));
    InMux I__7098 (
            .O(N__28904),
            .I(N__28885));
    Odrv4 I__7097 (
            .O(N__28901),
            .I(\tok.n2743 ));
    Odrv4 I__7096 (
            .O(N__28898),
            .I(\tok.n2743 ));
    Odrv4 I__7095 (
            .O(N__28893),
            .I(\tok.n2743 ));
    Odrv12 I__7094 (
            .O(N__28888),
            .I(\tok.n2743 ));
    LocalMux I__7093 (
            .O(N__28885),
            .I(\tok.n2743 ));
    InMux I__7092 (
            .O(N__28874),
            .I(N__28871));
    LocalMux I__7091 (
            .O(N__28871),
            .I(\tok.n5520 ));
    InMux I__7090 (
            .O(N__28868),
            .I(N__28863));
    InMux I__7089 (
            .O(N__28867),
            .I(N__28860));
    InMux I__7088 (
            .O(N__28866),
            .I(N__28854));
    LocalMux I__7087 (
            .O(N__28863),
            .I(N__28851));
    LocalMux I__7086 (
            .O(N__28860),
            .I(N__28847));
    InMux I__7085 (
            .O(N__28859),
            .I(N__28844));
    InMux I__7084 (
            .O(N__28858),
            .I(N__28841));
    InMux I__7083 (
            .O(N__28857),
            .I(N__28838));
    LocalMux I__7082 (
            .O(N__28854),
            .I(N__28834));
    Span4Mux_s3_v I__7081 (
            .O(N__28851),
            .I(N__28831));
    InMux I__7080 (
            .O(N__28850),
            .I(N__28828));
    Span4Mux_h I__7079 (
            .O(N__28847),
            .I(N__28823));
    LocalMux I__7078 (
            .O(N__28844),
            .I(N__28823));
    LocalMux I__7077 (
            .O(N__28841),
            .I(N__28818));
    LocalMux I__7076 (
            .O(N__28838),
            .I(N__28818));
    CascadeMux I__7075 (
            .O(N__28837),
            .I(N__28815));
    Span4Mux_v I__7074 (
            .O(N__28834),
            .I(N__28812));
    Span4Mux_h I__7073 (
            .O(N__28831),
            .I(N__28803));
    LocalMux I__7072 (
            .O(N__28828),
            .I(N__28803));
    Span4Mux_h I__7071 (
            .O(N__28823),
            .I(N__28803));
    Span4Mux_v I__7070 (
            .O(N__28818),
            .I(N__28803));
    InMux I__7069 (
            .O(N__28815),
            .I(N__28800));
    Odrv4 I__7068 (
            .O(N__28812),
            .I(\tok.S_14 ));
    Odrv4 I__7067 (
            .O(N__28803),
            .I(\tok.S_14 ));
    LocalMux I__7066 (
            .O(N__28800),
            .I(\tok.S_14 ));
    CascadeMux I__7065 (
            .O(N__28793),
            .I(\tok.n18_adj_774_cascade_ ));
    InMux I__7064 (
            .O(N__28790),
            .I(N__28778));
    CascadeMux I__7063 (
            .O(N__28789),
            .I(N__28774));
    InMux I__7062 (
            .O(N__28788),
            .I(N__28771));
    InMux I__7061 (
            .O(N__28787),
            .I(N__28768));
    InMux I__7060 (
            .O(N__28786),
            .I(N__28763));
    InMux I__7059 (
            .O(N__28785),
            .I(N__28763));
    InMux I__7058 (
            .O(N__28784),
            .I(N__28759));
    InMux I__7057 (
            .O(N__28783),
            .I(N__28755));
    InMux I__7056 (
            .O(N__28782),
            .I(N__28752));
    InMux I__7055 (
            .O(N__28781),
            .I(N__28748));
    LocalMux I__7054 (
            .O(N__28778),
            .I(N__28745));
    InMux I__7053 (
            .O(N__28777),
            .I(N__28742));
    InMux I__7052 (
            .O(N__28774),
            .I(N__28739));
    LocalMux I__7051 (
            .O(N__28771),
            .I(N__28736));
    LocalMux I__7050 (
            .O(N__28768),
            .I(N__28731));
    LocalMux I__7049 (
            .O(N__28763),
            .I(N__28731));
    CascadeMux I__7048 (
            .O(N__28762),
            .I(N__28727));
    LocalMux I__7047 (
            .O(N__28759),
            .I(N__28724));
    InMux I__7046 (
            .O(N__28758),
            .I(N__28721));
    LocalMux I__7045 (
            .O(N__28755),
            .I(N__28716));
    LocalMux I__7044 (
            .O(N__28752),
            .I(N__28716));
    InMux I__7043 (
            .O(N__28751),
            .I(N__28713));
    LocalMux I__7042 (
            .O(N__28748),
            .I(N__28704));
    Span4Mux_h I__7041 (
            .O(N__28745),
            .I(N__28704));
    LocalMux I__7040 (
            .O(N__28742),
            .I(N__28704));
    LocalMux I__7039 (
            .O(N__28739),
            .I(N__28704));
    Span4Mux_v I__7038 (
            .O(N__28736),
            .I(N__28699));
    Span4Mux_v I__7037 (
            .O(N__28731),
            .I(N__28699));
    InMux I__7036 (
            .O(N__28730),
            .I(N__28696));
    InMux I__7035 (
            .O(N__28727),
            .I(N__28693));
    Span4Mux_s3_h I__7034 (
            .O(N__28724),
            .I(N__28686));
    LocalMux I__7033 (
            .O(N__28721),
            .I(N__28686));
    Span4Mux_v I__7032 (
            .O(N__28716),
            .I(N__28686));
    LocalMux I__7031 (
            .O(N__28713),
            .I(N__28683));
    Span4Mux_v I__7030 (
            .O(N__28704),
            .I(N__28678));
    Span4Mux_h I__7029 (
            .O(N__28699),
            .I(N__28678));
    LocalMux I__7028 (
            .O(N__28696),
            .I(\tok.n2661 ));
    LocalMux I__7027 (
            .O(N__28693),
            .I(\tok.n2661 ));
    Odrv4 I__7026 (
            .O(N__28686),
            .I(\tok.n2661 ));
    Odrv12 I__7025 (
            .O(N__28683),
            .I(\tok.n2661 ));
    Odrv4 I__7024 (
            .O(N__28678),
            .I(\tok.n2661 ));
    InMux I__7023 (
            .O(N__28667),
            .I(N__28664));
    LocalMux I__7022 (
            .O(N__28664),
            .I(N__28661));
    Odrv12 I__7021 (
            .O(N__28661),
            .I(\tok.n5518 ));
    CascadeMux I__7020 (
            .O(N__28658),
            .I(N__28654));
    CascadeMux I__7019 (
            .O(N__28657),
            .I(N__28649));
    InMux I__7018 (
            .O(N__28654),
            .I(N__28639));
    InMux I__7017 (
            .O(N__28653),
            .I(N__28639));
    InMux I__7016 (
            .O(N__28652),
            .I(N__28639));
    InMux I__7015 (
            .O(N__28649),
            .I(N__28639));
    InMux I__7014 (
            .O(N__28648),
            .I(N__28633));
    LocalMux I__7013 (
            .O(N__28639),
            .I(N__28630));
    CascadeMux I__7012 (
            .O(N__28638),
            .I(N__28627));
    CascadeMux I__7011 (
            .O(N__28637),
            .I(N__28621));
    CascadeMux I__7010 (
            .O(N__28636),
            .I(N__28615));
    LocalMux I__7009 (
            .O(N__28633),
            .I(N__28610));
    Span4Mux_h I__7008 (
            .O(N__28630),
            .I(N__28610));
    InMux I__7007 (
            .O(N__28627),
            .I(N__28605));
    InMux I__7006 (
            .O(N__28626),
            .I(N__28605));
    InMux I__7005 (
            .O(N__28625),
            .I(N__28590));
    InMux I__7004 (
            .O(N__28624),
            .I(N__28590));
    InMux I__7003 (
            .O(N__28621),
            .I(N__28590));
    InMux I__7002 (
            .O(N__28620),
            .I(N__28590));
    InMux I__7001 (
            .O(N__28619),
            .I(N__28590));
    InMux I__7000 (
            .O(N__28618),
            .I(N__28590));
    InMux I__6999 (
            .O(N__28615),
            .I(N__28590));
    Span4Mux_v I__6998 (
            .O(N__28610),
            .I(N__28583));
    LocalMux I__6997 (
            .O(N__28605),
            .I(N__28583));
    LocalMux I__6996 (
            .O(N__28590),
            .I(N__28579));
    InMux I__6995 (
            .O(N__28589),
            .I(N__28574));
    InMux I__6994 (
            .O(N__28588),
            .I(N__28574));
    Span4Mux_v I__6993 (
            .O(N__28583),
            .I(N__28571));
    InMux I__6992 (
            .O(N__28582),
            .I(N__28568));
    Span4Mux_v I__6991 (
            .O(N__28579),
            .I(N__28563));
    LocalMux I__6990 (
            .O(N__28574),
            .I(N__28563));
    Span4Mux_h I__6989 (
            .O(N__28571),
            .I(N__28558));
    LocalMux I__6988 (
            .O(N__28568),
            .I(N__28558));
    Span4Mux_v I__6987 (
            .O(N__28563),
            .I(N__28555));
    Span4Mux_h I__6986 (
            .O(N__28558),
            .I(N__28552));
    Odrv4 I__6985 (
            .O(N__28555),
            .I(\tok.n23 ));
    Odrv4 I__6984 (
            .O(N__28552),
            .I(\tok.n23 ));
    CascadeMux I__6983 (
            .O(N__28547),
            .I(\tok.n22_adj_676_cascade_ ));
    ClkMux I__6982 (
            .O(N__28544),
            .I(N__28307));
    ClkMux I__6981 (
            .O(N__28543),
            .I(N__28307));
    ClkMux I__6980 (
            .O(N__28542),
            .I(N__28307));
    ClkMux I__6979 (
            .O(N__28541),
            .I(N__28307));
    ClkMux I__6978 (
            .O(N__28540),
            .I(N__28307));
    ClkMux I__6977 (
            .O(N__28539),
            .I(N__28307));
    ClkMux I__6976 (
            .O(N__28538),
            .I(N__28307));
    ClkMux I__6975 (
            .O(N__28537),
            .I(N__28307));
    ClkMux I__6974 (
            .O(N__28536),
            .I(N__28307));
    ClkMux I__6973 (
            .O(N__28535),
            .I(N__28307));
    ClkMux I__6972 (
            .O(N__28534),
            .I(N__28307));
    ClkMux I__6971 (
            .O(N__28533),
            .I(N__28307));
    ClkMux I__6970 (
            .O(N__28532),
            .I(N__28307));
    ClkMux I__6969 (
            .O(N__28531),
            .I(N__28307));
    ClkMux I__6968 (
            .O(N__28530),
            .I(N__28307));
    ClkMux I__6967 (
            .O(N__28529),
            .I(N__28307));
    ClkMux I__6966 (
            .O(N__28528),
            .I(N__28307));
    ClkMux I__6965 (
            .O(N__28527),
            .I(N__28307));
    ClkMux I__6964 (
            .O(N__28526),
            .I(N__28307));
    ClkMux I__6963 (
            .O(N__28525),
            .I(N__28307));
    ClkMux I__6962 (
            .O(N__28524),
            .I(N__28307));
    ClkMux I__6961 (
            .O(N__28523),
            .I(N__28307));
    ClkMux I__6960 (
            .O(N__28522),
            .I(N__28307));
    ClkMux I__6959 (
            .O(N__28521),
            .I(N__28307));
    ClkMux I__6958 (
            .O(N__28520),
            .I(N__28307));
    ClkMux I__6957 (
            .O(N__28519),
            .I(N__28307));
    ClkMux I__6956 (
            .O(N__28518),
            .I(N__28307));
    ClkMux I__6955 (
            .O(N__28517),
            .I(N__28307));
    ClkMux I__6954 (
            .O(N__28516),
            .I(N__28307));
    ClkMux I__6953 (
            .O(N__28515),
            .I(N__28307));
    ClkMux I__6952 (
            .O(N__28514),
            .I(N__28307));
    ClkMux I__6951 (
            .O(N__28513),
            .I(N__28307));
    ClkMux I__6950 (
            .O(N__28512),
            .I(N__28307));
    ClkMux I__6949 (
            .O(N__28511),
            .I(N__28307));
    ClkMux I__6948 (
            .O(N__28510),
            .I(N__28307));
    ClkMux I__6947 (
            .O(N__28509),
            .I(N__28307));
    ClkMux I__6946 (
            .O(N__28508),
            .I(N__28307));
    ClkMux I__6945 (
            .O(N__28507),
            .I(N__28307));
    ClkMux I__6944 (
            .O(N__28506),
            .I(N__28307));
    ClkMux I__6943 (
            .O(N__28505),
            .I(N__28307));
    ClkMux I__6942 (
            .O(N__28504),
            .I(N__28307));
    ClkMux I__6941 (
            .O(N__28503),
            .I(N__28307));
    ClkMux I__6940 (
            .O(N__28502),
            .I(N__28307));
    ClkMux I__6939 (
            .O(N__28501),
            .I(N__28307));
    ClkMux I__6938 (
            .O(N__28500),
            .I(N__28307));
    ClkMux I__6937 (
            .O(N__28499),
            .I(N__28307));
    ClkMux I__6936 (
            .O(N__28498),
            .I(N__28307));
    ClkMux I__6935 (
            .O(N__28497),
            .I(N__28307));
    ClkMux I__6934 (
            .O(N__28496),
            .I(N__28307));
    ClkMux I__6933 (
            .O(N__28495),
            .I(N__28307));
    ClkMux I__6932 (
            .O(N__28494),
            .I(N__28307));
    ClkMux I__6931 (
            .O(N__28493),
            .I(N__28307));
    ClkMux I__6930 (
            .O(N__28492),
            .I(N__28307));
    ClkMux I__6929 (
            .O(N__28491),
            .I(N__28307));
    ClkMux I__6928 (
            .O(N__28490),
            .I(N__28307));
    ClkMux I__6927 (
            .O(N__28489),
            .I(N__28307));
    ClkMux I__6926 (
            .O(N__28488),
            .I(N__28307));
    ClkMux I__6925 (
            .O(N__28487),
            .I(N__28307));
    ClkMux I__6924 (
            .O(N__28486),
            .I(N__28307));
    ClkMux I__6923 (
            .O(N__28485),
            .I(N__28307));
    ClkMux I__6922 (
            .O(N__28484),
            .I(N__28307));
    ClkMux I__6921 (
            .O(N__28483),
            .I(N__28307));
    ClkMux I__6920 (
            .O(N__28482),
            .I(N__28307));
    ClkMux I__6919 (
            .O(N__28481),
            .I(N__28307));
    ClkMux I__6918 (
            .O(N__28480),
            .I(N__28307));
    ClkMux I__6917 (
            .O(N__28479),
            .I(N__28307));
    ClkMux I__6916 (
            .O(N__28478),
            .I(N__28307));
    ClkMux I__6915 (
            .O(N__28477),
            .I(N__28307));
    ClkMux I__6914 (
            .O(N__28476),
            .I(N__28307));
    ClkMux I__6913 (
            .O(N__28475),
            .I(N__28307));
    ClkMux I__6912 (
            .O(N__28474),
            .I(N__28307));
    ClkMux I__6911 (
            .O(N__28473),
            .I(N__28307));
    ClkMux I__6910 (
            .O(N__28472),
            .I(N__28307));
    ClkMux I__6909 (
            .O(N__28471),
            .I(N__28307));
    ClkMux I__6908 (
            .O(N__28470),
            .I(N__28307));
    ClkMux I__6907 (
            .O(N__28469),
            .I(N__28307));
    ClkMux I__6906 (
            .O(N__28468),
            .I(N__28307));
    ClkMux I__6905 (
            .O(N__28467),
            .I(N__28307));
    ClkMux I__6904 (
            .O(N__28466),
            .I(N__28307));
    GlobalMux I__6903 (
            .O(N__28307),
            .I(N__28304));
    DummyBuf I__6902 (
            .O(N__28304),
            .I(clk));
    CEMux I__6901 (
            .O(N__28301),
            .I(N__28297));
    CEMux I__6900 (
            .O(N__28300),
            .I(N__28293));
    LocalMux I__6899 (
            .O(N__28297),
            .I(N__28289));
    CEMux I__6898 (
            .O(N__28296),
            .I(N__28286));
    LocalMux I__6897 (
            .O(N__28293),
            .I(N__28282));
    CEMux I__6896 (
            .O(N__28292),
            .I(N__28279));
    Span4Mux_s3_h I__6895 (
            .O(N__28289),
            .I(N__28274));
    LocalMux I__6894 (
            .O(N__28286),
            .I(N__28274));
    CEMux I__6893 (
            .O(N__28285),
            .I(N__28271));
    Span4Mux_h I__6892 (
            .O(N__28282),
            .I(N__28268));
    LocalMux I__6891 (
            .O(N__28279),
            .I(N__28265));
    Span4Mux_v I__6890 (
            .O(N__28274),
            .I(N__28262));
    LocalMux I__6889 (
            .O(N__28271),
            .I(N__28259));
    Span4Mux_s1_h I__6888 (
            .O(N__28268),
            .I(N__28254));
    Span4Mux_v I__6887 (
            .O(N__28265),
            .I(N__28254));
    Span4Mux_v I__6886 (
            .O(N__28262),
            .I(N__28251));
    Span4Mux_v I__6885 (
            .O(N__28259),
            .I(N__28246));
    Span4Mux_h I__6884 (
            .O(N__28254),
            .I(N__28246));
    Sp12to4 I__6883 (
            .O(N__28251),
            .I(N__28243));
    Odrv4 I__6882 (
            .O(N__28246),
            .I(\tok.n995 ));
    Odrv12 I__6881 (
            .O(N__28243),
            .I(\tok.n995 ));
    SRMux I__6880 (
            .O(N__28238),
            .I(N__28227));
    SRMux I__6879 (
            .O(N__28237),
            .I(N__28223));
    SRMux I__6878 (
            .O(N__28236),
            .I(N__28220));
    SRMux I__6877 (
            .O(N__28235),
            .I(N__28217));
    SRMux I__6876 (
            .O(N__28234),
            .I(N__28214));
    SRMux I__6875 (
            .O(N__28233),
            .I(N__28209));
    SRMux I__6874 (
            .O(N__28232),
            .I(N__28206));
    SRMux I__6873 (
            .O(N__28231),
            .I(N__28202));
    SRMux I__6872 (
            .O(N__28230),
            .I(N__28199));
    LocalMux I__6871 (
            .O(N__28227),
            .I(N__28196));
    SRMux I__6870 (
            .O(N__28226),
            .I(N__28193));
    LocalMux I__6869 (
            .O(N__28223),
            .I(N__28189));
    LocalMux I__6868 (
            .O(N__28220),
            .I(N__28186));
    LocalMux I__6867 (
            .O(N__28217),
            .I(N__28181));
    LocalMux I__6866 (
            .O(N__28214),
            .I(N__28181));
    SRMux I__6865 (
            .O(N__28213),
            .I(N__28178));
    SRMux I__6864 (
            .O(N__28212),
            .I(N__28175));
    LocalMux I__6863 (
            .O(N__28209),
            .I(N__28171));
    LocalMux I__6862 (
            .O(N__28206),
            .I(N__28168));
    SRMux I__6861 (
            .O(N__28205),
            .I(N__28165));
    LocalMux I__6860 (
            .O(N__28202),
            .I(N__28162));
    LocalMux I__6859 (
            .O(N__28199),
            .I(N__28159));
    Span4Mux_v I__6858 (
            .O(N__28196),
            .I(N__28154));
    LocalMux I__6857 (
            .O(N__28193),
            .I(N__28154));
    SRMux I__6856 (
            .O(N__28192),
            .I(N__28151));
    Span4Mux_h I__6855 (
            .O(N__28189),
            .I(N__28140));
    Span4Mux_h I__6854 (
            .O(N__28186),
            .I(N__28140));
    Span4Mux_s3_v I__6853 (
            .O(N__28181),
            .I(N__28140));
    LocalMux I__6852 (
            .O(N__28178),
            .I(N__28140));
    LocalMux I__6851 (
            .O(N__28175),
            .I(N__28140));
    SRMux I__6850 (
            .O(N__28174),
            .I(N__28137));
    Span4Mux_v I__6849 (
            .O(N__28171),
            .I(N__28134));
    Span4Mux_v I__6848 (
            .O(N__28168),
            .I(N__28129));
    LocalMux I__6847 (
            .O(N__28165),
            .I(N__28129));
    Span4Mux_s3_h I__6846 (
            .O(N__28162),
            .I(N__28125));
    Span4Mux_v I__6845 (
            .O(N__28159),
            .I(N__28122));
    Span4Mux_h I__6844 (
            .O(N__28154),
            .I(N__28117));
    LocalMux I__6843 (
            .O(N__28151),
            .I(N__28117));
    Span4Mux_v I__6842 (
            .O(N__28140),
            .I(N__28114));
    LocalMux I__6841 (
            .O(N__28137),
            .I(N__28111));
    Span4Mux_v I__6840 (
            .O(N__28134),
            .I(N__28108));
    Span4Mux_v I__6839 (
            .O(N__28129),
            .I(N__28105));
    SRMux I__6838 (
            .O(N__28128),
            .I(N__28102));
    Span4Mux_h I__6837 (
            .O(N__28125),
            .I(N__28099));
    Span4Mux_h I__6836 (
            .O(N__28122),
            .I(N__28094));
    Span4Mux_h I__6835 (
            .O(N__28117),
            .I(N__28094));
    Span4Mux_v I__6834 (
            .O(N__28114),
            .I(N__28089));
    Span4Mux_h I__6833 (
            .O(N__28111),
            .I(N__28089));
    Span4Mux_h I__6832 (
            .O(N__28108),
            .I(N__28082));
    Span4Mux_v I__6831 (
            .O(N__28105),
            .I(N__28082));
    LocalMux I__6830 (
            .O(N__28102),
            .I(N__28082));
    Odrv4 I__6829 (
            .O(N__28099),
            .I(\tok.reset_N_2 ));
    Odrv4 I__6828 (
            .O(N__28094),
            .I(\tok.reset_N_2 ));
    Odrv4 I__6827 (
            .O(N__28089),
            .I(\tok.reset_N_2 ));
    Odrv4 I__6826 (
            .O(N__28082),
            .I(\tok.reset_N_2 ));
    CascadeMux I__6825 (
            .O(N__28073),
            .I(N__28068));
    InMux I__6824 (
            .O(N__28072),
            .I(N__28061));
    InMux I__6823 (
            .O(N__28071),
            .I(N__28061));
    InMux I__6822 (
            .O(N__28068),
            .I(N__28058));
    CascadeMux I__6821 (
            .O(N__28067),
            .I(N__28054));
    CascadeMux I__6820 (
            .O(N__28066),
            .I(N__28051));
    LocalMux I__6819 (
            .O(N__28061),
            .I(N__28048));
    LocalMux I__6818 (
            .O(N__28058),
            .I(N__28045));
    InMux I__6817 (
            .O(N__28057),
            .I(N__28042));
    InMux I__6816 (
            .O(N__28054),
            .I(N__28039));
    InMux I__6815 (
            .O(N__28051),
            .I(N__28036));
    Span4Mux_v I__6814 (
            .O(N__28048),
            .I(N__28032));
    Span4Mux_v I__6813 (
            .O(N__28045),
            .I(N__28029));
    LocalMux I__6812 (
            .O(N__28042),
            .I(N__28025));
    LocalMux I__6811 (
            .O(N__28039),
            .I(N__28022));
    LocalMux I__6810 (
            .O(N__28036),
            .I(N__28019));
    InMux I__6809 (
            .O(N__28035),
            .I(N__28016));
    Span4Mux_s1_h I__6808 (
            .O(N__28032),
            .I(N__28013));
    Span4Mux_h I__6807 (
            .O(N__28029),
            .I(N__28010));
    InMux I__6806 (
            .O(N__28028),
            .I(N__28007));
    Span4Mux_h I__6805 (
            .O(N__28025),
            .I(N__28004));
    Span4Mux_v I__6804 (
            .O(N__28022),
            .I(N__27999));
    Span4Mux_h I__6803 (
            .O(N__28019),
            .I(N__27999));
    LocalMux I__6802 (
            .O(N__28016),
            .I(\tok.S_8 ));
    Odrv4 I__6801 (
            .O(N__28013),
            .I(\tok.S_8 ));
    Odrv4 I__6800 (
            .O(N__28010),
            .I(\tok.S_8 ));
    LocalMux I__6799 (
            .O(N__28007),
            .I(\tok.S_8 ));
    Odrv4 I__6798 (
            .O(N__28004),
            .I(\tok.S_8 ));
    Odrv4 I__6797 (
            .O(N__27999),
            .I(\tok.S_8 ));
    CascadeMux I__6796 (
            .O(N__27986),
            .I(N__27983));
    InMux I__6795 (
            .O(N__27983),
            .I(N__27980));
    LocalMux I__6794 (
            .O(N__27980),
            .I(\tok.n5544 ));
    InMux I__6793 (
            .O(N__27977),
            .I(N__27974));
    LocalMux I__6792 (
            .O(N__27974),
            .I(\tok.n5542 ));
    InMux I__6791 (
            .O(N__27971),
            .I(N__27968));
    LocalMux I__6790 (
            .O(N__27968),
            .I(N__27965));
    Span4Mux_v I__6789 (
            .O(N__27965),
            .I(N__27962));
    Odrv4 I__6788 (
            .O(N__27962),
            .I(\tok.n10_adj_666 ));
    CascadeMux I__6787 (
            .O(N__27959),
            .I(N__27954));
    InMux I__6786 (
            .O(N__27958),
            .I(N__27950));
    InMux I__6785 (
            .O(N__27957),
            .I(N__27947));
    InMux I__6784 (
            .O(N__27954),
            .I(N__27944));
    CascadeMux I__6783 (
            .O(N__27953),
            .I(N__27941));
    LocalMux I__6782 (
            .O(N__27950),
            .I(N__27935));
    LocalMux I__6781 (
            .O(N__27947),
            .I(N__27935));
    LocalMux I__6780 (
            .O(N__27944),
            .I(N__27932));
    InMux I__6779 (
            .O(N__27941),
            .I(N__27929));
    InMux I__6778 (
            .O(N__27940),
            .I(N__27926));
    Span4Mux_v I__6777 (
            .O(N__27935),
            .I(N__27923));
    Span4Mux_s3_v I__6776 (
            .O(N__27932),
            .I(N__27918));
    LocalMux I__6775 (
            .O(N__27929),
            .I(N__27918));
    LocalMux I__6774 (
            .O(N__27926),
            .I(N__27915));
    Span4Mux_h I__6773 (
            .O(N__27923),
            .I(N__27908));
    Span4Mux_v I__6772 (
            .O(N__27918),
            .I(N__27908));
    Span4Mux_v I__6771 (
            .O(N__27915),
            .I(N__27905));
    InMux I__6770 (
            .O(N__27914),
            .I(N__27900));
    InMux I__6769 (
            .O(N__27913),
            .I(N__27900));
    Odrv4 I__6768 (
            .O(N__27908),
            .I(\tok.n15_adj_667 ));
    Odrv4 I__6767 (
            .O(N__27905),
            .I(\tok.n15_adj_667 ));
    LocalMux I__6766 (
            .O(N__27900),
            .I(\tok.n15_adj_667 ));
    InMux I__6765 (
            .O(N__27893),
            .I(N__27890));
    LocalMux I__6764 (
            .O(N__27890),
            .I(\tok.n14_adj_668 ));
    CascadeMux I__6763 (
            .O(N__27887),
            .I(N__27879));
    InMux I__6762 (
            .O(N__27886),
            .I(N__27869));
    InMux I__6761 (
            .O(N__27885),
            .I(N__27869));
    InMux I__6760 (
            .O(N__27884),
            .I(N__27864));
    InMux I__6759 (
            .O(N__27883),
            .I(N__27864));
    InMux I__6758 (
            .O(N__27882),
            .I(N__27859));
    InMux I__6757 (
            .O(N__27879),
            .I(N__27859));
    CascadeMux I__6756 (
            .O(N__27878),
            .I(N__27851));
    InMux I__6755 (
            .O(N__27877),
            .I(N__27847));
    InMux I__6754 (
            .O(N__27876),
            .I(N__27840));
    InMux I__6753 (
            .O(N__27875),
            .I(N__27840));
    InMux I__6752 (
            .O(N__27874),
            .I(N__27840));
    LocalMux I__6751 (
            .O(N__27869),
            .I(N__27835));
    LocalMux I__6750 (
            .O(N__27864),
            .I(N__27835));
    LocalMux I__6749 (
            .O(N__27859),
            .I(N__27832));
    InMux I__6748 (
            .O(N__27858),
            .I(N__27825));
    InMux I__6747 (
            .O(N__27857),
            .I(N__27825));
    InMux I__6746 (
            .O(N__27856),
            .I(N__27825));
    InMux I__6745 (
            .O(N__27855),
            .I(N__27818));
    InMux I__6744 (
            .O(N__27854),
            .I(N__27818));
    InMux I__6743 (
            .O(N__27851),
            .I(N__27818));
    InMux I__6742 (
            .O(N__27850),
            .I(N__27815));
    LocalMux I__6741 (
            .O(N__27847),
            .I(N__27810));
    LocalMux I__6740 (
            .O(N__27840),
            .I(N__27810));
    Span4Mux_v I__6739 (
            .O(N__27835),
            .I(N__27807));
    Span4Mux_h I__6738 (
            .O(N__27832),
            .I(N__27800));
    LocalMux I__6737 (
            .O(N__27825),
            .I(N__27800));
    LocalMux I__6736 (
            .O(N__27818),
            .I(N__27800));
    LocalMux I__6735 (
            .O(N__27815),
            .I(N__27797));
    Span4Mux_v I__6734 (
            .O(N__27810),
            .I(N__27790));
    Span4Mux_h I__6733 (
            .O(N__27807),
            .I(N__27790));
    Span4Mux_v I__6732 (
            .O(N__27800),
            .I(N__27790));
    Odrv4 I__6731 (
            .O(N__27797),
            .I(\tok.n880 ));
    Odrv4 I__6730 (
            .O(N__27790),
            .I(\tok.n880 ));
    InMux I__6729 (
            .O(N__27785),
            .I(N__27775));
    InMux I__6728 (
            .O(N__27784),
            .I(N__27775));
    InMux I__6727 (
            .O(N__27783),
            .I(N__27771));
    CascadeMux I__6726 (
            .O(N__27782),
            .I(N__27767));
    InMux I__6725 (
            .O(N__27781),
            .I(N__27763));
    InMux I__6724 (
            .O(N__27780),
            .I(N__27760));
    LocalMux I__6723 (
            .O(N__27775),
            .I(N__27757));
    InMux I__6722 (
            .O(N__27774),
            .I(N__27751));
    LocalMux I__6721 (
            .O(N__27771),
            .I(N__27748));
    InMux I__6720 (
            .O(N__27770),
            .I(N__27745));
    InMux I__6719 (
            .O(N__27767),
            .I(N__27742));
    InMux I__6718 (
            .O(N__27766),
            .I(N__27739));
    LocalMux I__6717 (
            .O(N__27763),
            .I(N__27735));
    LocalMux I__6716 (
            .O(N__27760),
            .I(N__27732));
    Span4Mux_s2_h I__6715 (
            .O(N__27757),
            .I(N__27729));
    InMux I__6714 (
            .O(N__27756),
            .I(N__27726));
    InMux I__6713 (
            .O(N__27755),
            .I(N__27722));
    InMux I__6712 (
            .O(N__27754),
            .I(N__27719));
    LocalMux I__6711 (
            .O(N__27751),
            .I(N__27716));
    Span4Mux_s2_v I__6710 (
            .O(N__27748),
            .I(N__27709));
    LocalMux I__6709 (
            .O(N__27745),
            .I(N__27709));
    LocalMux I__6708 (
            .O(N__27742),
            .I(N__27709));
    LocalMux I__6707 (
            .O(N__27739),
            .I(N__27706));
    InMux I__6706 (
            .O(N__27738),
            .I(N__27703));
    Span4Mux_v I__6705 (
            .O(N__27735),
            .I(N__27694));
    Span4Mux_v I__6704 (
            .O(N__27732),
            .I(N__27694));
    Span4Mux_h I__6703 (
            .O(N__27729),
            .I(N__27694));
    LocalMux I__6702 (
            .O(N__27726),
            .I(N__27694));
    InMux I__6701 (
            .O(N__27725),
            .I(N__27691));
    LocalMux I__6700 (
            .O(N__27722),
            .I(N__27687));
    LocalMux I__6699 (
            .O(N__27719),
            .I(N__27676));
    Span4Mux_v I__6698 (
            .O(N__27716),
            .I(N__27676));
    Span4Mux_v I__6697 (
            .O(N__27709),
            .I(N__27676));
    Span4Mux_v I__6696 (
            .O(N__27706),
            .I(N__27676));
    LocalMux I__6695 (
            .O(N__27703),
            .I(N__27676));
    Span4Mux_h I__6694 (
            .O(N__27694),
            .I(N__27671));
    LocalMux I__6693 (
            .O(N__27691),
            .I(N__27671));
    InMux I__6692 (
            .O(N__27690),
            .I(N__27668));
    Span4Mux_h I__6691 (
            .O(N__27687),
            .I(N__27663));
    Span4Mux_h I__6690 (
            .O(N__27676),
            .I(N__27663));
    Odrv4 I__6689 (
            .O(N__27671),
            .I(\tok.A_low_0 ));
    LocalMux I__6688 (
            .O(N__27668),
            .I(\tok.A_low_0 ));
    Odrv4 I__6687 (
            .O(N__27663),
            .I(\tok.A_low_0 ));
    InMux I__6686 (
            .O(N__27656),
            .I(N__27644));
    InMux I__6685 (
            .O(N__27655),
            .I(N__27644));
    InMux I__6684 (
            .O(N__27654),
            .I(N__27639));
    InMux I__6683 (
            .O(N__27653),
            .I(N__27639));
    InMux I__6682 (
            .O(N__27652),
            .I(N__27634));
    InMux I__6681 (
            .O(N__27651),
            .I(N__27634));
    InMux I__6680 (
            .O(N__27650),
            .I(N__27626));
    InMux I__6679 (
            .O(N__27649),
            .I(N__27621));
    LocalMux I__6678 (
            .O(N__27644),
            .I(N__27618));
    LocalMux I__6677 (
            .O(N__27639),
            .I(N__27615));
    LocalMux I__6676 (
            .O(N__27634),
            .I(N__27612));
    InMux I__6675 (
            .O(N__27633),
            .I(N__27609));
    InMux I__6674 (
            .O(N__27632),
            .I(N__27602));
    InMux I__6673 (
            .O(N__27631),
            .I(N__27602));
    InMux I__6672 (
            .O(N__27630),
            .I(N__27602));
    InMux I__6671 (
            .O(N__27629),
            .I(N__27599));
    LocalMux I__6670 (
            .O(N__27626),
            .I(N__27596));
    InMux I__6669 (
            .O(N__27625),
            .I(N__27593));
    InMux I__6668 (
            .O(N__27624),
            .I(N__27590));
    LocalMux I__6667 (
            .O(N__27621),
            .I(N__27587));
    Span4Mux_s1_h I__6666 (
            .O(N__27618),
            .I(N__27582));
    Span4Mux_v I__6665 (
            .O(N__27615),
            .I(N__27582));
    Odrv4 I__6664 (
            .O(N__27612),
            .I(\tok.n904 ));
    LocalMux I__6663 (
            .O(N__27609),
            .I(\tok.n904 ));
    LocalMux I__6662 (
            .O(N__27602),
            .I(\tok.n904 ));
    LocalMux I__6661 (
            .O(N__27599),
            .I(\tok.n904 ));
    Odrv4 I__6660 (
            .O(N__27596),
            .I(\tok.n904 ));
    LocalMux I__6659 (
            .O(N__27593),
            .I(\tok.n904 ));
    LocalMux I__6658 (
            .O(N__27590),
            .I(\tok.n904 ));
    Odrv4 I__6657 (
            .O(N__27587),
            .I(\tok.n904 ));
    Odrv4 I__6656 (
            .O(N__27582),
            .I(\tok.n904 ));
    InMux I__6655 (
            .O(N__27563),
            .I(N__27560));
    LocalMux I__6654 (
            .O(N__27560),
            .I(N__27557));
    Odrv12 I__6653 (
            .O(N__27557),
            .I(\tok.n5372 ));
    CascadeMux I__6652 (
            .O(N__27554),
            .I(N__27551));
    InMux I__6651 (
            .O(N__27551),
            .I(N__27546));
    InMux I__6650 (
            .O(N__27550),
            .I(N__27540));
    InMux I__6649 (
            .O(N__27549),
            .I(N__27540));
    LocalMux I__6648 (
            .O(N__27546),
            .I(N__27535));
    InMux I__6647 (
            .O(N__27545),
            .I(N__27532));
    LocalMux I__6646 (
            .O(N__27540),
            .I(N__27528));
    InMux I__6645 (
            .O(N__27539),
            .I(N__27525));
    InMux I__6644 (
            .O(N__27538),
            .I(N__27522));
    Span4Mux_s1_h I__6643 (
            .O(N__27535),
            .I(N__27517));
    LocalMux I__6642 (
            .O(N__27532),
            .I(N__27517));
    CascadeMux I__6641 (
            .O(N__27531),
            .I(N__27514));
    Span4Mux_v I__6640 (
            .O(N__27528),
            .I(N__27510));
    LocalMux I__6639 (
            .O(N__27525),
            .I(N__27507));
    LocalMux I__6638 (
            .O(N__27522),
            .I(N__27504));
    Span4Mux_h I__6637 (
            .O(N__27517),
            .I(N__27501));
    InMux I__6636 (
            .O(N__27514),
            .I(N__27498));
    InMux I__6635 (
            .O(N__27513),
            .I(N__27495));
    Span4Mux_v I__6634 (
            .O(N__27510),
            .I(N__27490));
    Span4Mux_v I__6633 (
            .O(N__27507),
            .I(N__27490));
    Span12Mux_s8_h I__6632 (
            .O(N__27504),
            .I(N__27483));
    Sp12to4 I__6631 (
            .O(N__27501),
            .I(N__27483));
    LocalMux I__6630 (
            .O(N__27498),
            .I(N__27483));
    LocalMux I__6629 (
            .O(N__27495),
            .I(\tok.S_9 ));
    Odrv4 I__6628 (
            .O(N__27490),
            .I(\tok.S_9 ));
    Odrv12 I__6627 (
            .O(N__27483),
            .I(\tok.S_9 ));
    InMux I__6626 (
            .O(N__27476),
            .I(N__27473));
    LocalMux I__6625 (
            .O(N__27473),
            .I(N__27470));
    Span4Mux_v I__6624 (
            .O(N__27470),
            .I(N__27467));
    Odrv4 I__6623 (
            .O(N__27467),
            .I(\tok.n8_adj_689 ));
    CascadeMux I__6622 (
            .O(N__27464),
            .I(N__27461));
    InMux I__6621 (
            .O(N__27461),
            .I(N__27456));
    CascadeMux I__6620 (
            .O(N__27460),
            .I(N__27453));
    CascadeMux I__6619 (
            .O(N__27459),
            .I(N__27449));
    LocalMux I__6618 (
            .O(N__27456),
            .I(N__27445));
    InMux I__6617 (
            .O(N__27453),
            .I(N__27442));
    InMux I__6616 (
            .O(N__27452),
            .I(N__27437));
    InMux I__6615 (
            .O(N__27449),
            .I(N__27434));
    CascadeMux I__6614 (
            .O(N__27448),
            .I(N__27431));
    Span4Mux_v I__6613 (
            .O(N__27445),
            .I(N__27426));
    LocalMux I__6612 (
            .O(N__27442),
            .I(N__27426));
    InMux I__6611 (
            .O(N__27441),
            .I(N__27423));
    InMux I__6610 (
            .O(N__27440),
            .I(N__27420));
    LocalMux I__6609 (
            .O(N__27437),
            .I(N__27415));
    LocalMux I__6608 (
            .O(N__27434),
            .I(N__27415));
    InMux I__6607 (
            .O(N__27431),
            .I(N__27411));
    Span4Mux_v I__6606 (
            .O(N__27426),
            .I(N__27408));
    LocalMux I__6605 (
            .O(N__27423),
            .I(N__27405));
    LocalMux I__6604 (
            .O(N__27420),
            .I(N__27402));
    Span4Mux_v I__6603 (
            .O(N__27415),
            .I(N__27399));
    InMux I__6602 (
            .O(N__27414),
            .I(N__27396));
    LocalMux I__6601 (
            .O(N__27411),
            .I(N__27393));
    Span4Mux_h I__6600 (
            .O(N__27408),
            .I(N__27390));
    Span4Mux_v I__6599 (
            .O(N__27405),
            .I(N__27387));
    Span4Mux_v I__6598 (
            .O(N__27402),
            .I(N__27382));
    Span4Mux_h I__6597 (
            .O(N__27399),
            .I(N__27382));
    LocalMux I__6596 (
            .O(N__27396),
            .I(\tok.S_10 ));
    Odrv12 I__6595 (
            .O(N__27393),
            .I(\tok.S_10 ));
    Odrv4 I__6594 (
            .O(N__27390),
            .I(\tok.S_10 ));
    Odrv4 I__6593 (
            .O(N__27387),
            .I(\tok.S_10 ));
    Odrv4 I__6592 (
            .O(N__27382),
            .I(\tok.S_10 ));
    InMux I__6591 (
            .O(N__27371),
            .I(N__27368));
    LocalMux I__6590 (
            .O(N__27368),
            .I(N__27365));
    Odrv12 I__6589 (
            .O(N__27365),
            .I(\tok.n8_adj_702 ));
    CascadeMux I__6588 (
            .O(N__27362),
            .I(N__27359));
    InMux I__6587 (
            .O(N__27359),
            .I(N__27356));
    LocalMux I__6586 (
            .O(N__27356),
            .I(\tok.n298 ));
    CascadeMux I__6585 (
            .O(N__27353),
            .I(N__27348));
    InMux I__6584 (
            .O(N__27352),
            .I(N__27344));
    CascadeMux I__6583 (
            .O(N__27351),
            .I(N__27340));
    InMux I__6582 (
            .O(N__27348),
            .I(N__27337));
    InMux I__6581 (
            .O(N__27347),
            .I(N__27334));
    LocalMux I__6580 (
            .O(N__27344),
            .I(N__27331));
    InMux I__6579 (
            .O(N__27343),
            .I(N__27328));
    InMux I__6578 (
            .O(N__27340),
            .I(N__27321));
    LocalMux I__6577 (
            .O(N__27337),
            .I(N__27318));
    LocalMux I__6576 (
            .O(N__27334),
            .I(N__27313));
    Span4Mux_h I__6575 (
            .O(N__27331),
            .I(N__27313));
    LocalMux I__6574 (
            .O(N__27328),
            .I(N__27310));
    InMux I__6573 (
            .O(N__27327),
            .I(N__27307));
    InMux I__6572 (
            .O(N__27326),
            .I(N__27304));
    InMux I__6571 (
            .O(N__27325),
            .I(N__27298));
    InMux I__6570 (
            .O(N__27324),
            .I(N__27298));
    LocalMux I__6569 (
            .O(N__27321),
            .I(N__27293));
    Span4Mux_h I__6568 (
            .O(N__27318),
            .I(N__27287));
    Span4Mux_h I__6567 (
            .O(N__27313),
            .I(N__27280));
    Span4Mux_s3_v I__6566 (
            .O(N__27310),
            .I(N__27280));
    LocalMux I__6565 (
            .O(N__27307),
            .I(N__27280));
    LocalMux I__6564 (
            .O(N__27304),
            .I(N__27277));
    InMux I__6563 (
            .O(N__27303),
            .I(N__27274));
    LocalMux I__6562 (
            .O(N__27298),
            .I(N__27271));
    InMux I__6561 (
            .O(N__27297),
            .I(N__27266));
    InMux I__6560 (
            .O(N__27296),
            .I(N__27266));
    Span4Mux_h I__6559 (
            .O(N__27293),
            .I(N__27263));
    InMux I__6558 (
            .O(N__27292),
            .I(N__27260));
    InMux I__6557 (
            .O(N__27291),
            .I(N__27255));
    InMux I__6556 (
            .O(N__27290),
            .I(N__27255));
    Span4Mux_v I__6555 (
            .O(N__27287),
            .I(N__27250));
    Span4Mux_v I__6554 (
            .O(N__27280),
            .I(N__27250));
    Span12Mux_s7_v I__6553 (
            .O(N__27277),
            .I(N__27245));
    LocalMux I__6552 (
            .O(N__27274),
            .I(N__27245));
    Span4Mux_h I__6551 (
            .O(N__27271),
            .I(N__27238));
    LocalMux I__6550 (
            .O(N__27266),
            .I(N__27238));
    Span4Mux_h I__6549 (
            .O(N__27263),
            .I(N__27238));
    LocalMux I__6548 (
            .O(N__27260),
            .I(\tok.A_low_5 ));
    LocalMux I__6547 (
            .O(N__27255),
            .I(\tok.A_low_5 ));
    Odrv4 I__6546 (
            .O(N__27250),
            .I(\tok.A_low_5 ));
    Odrv12 I__6545 (
            .O(N__27245),
            .I(\tok.A_low_5 ));
    Odrv4 I__6544 (
            .O(N__27238),
            .I(\tok.A_low_5 ));
    InMux I__6543 (
            .O(N__27227),
            .I(N__27224));
    LocalMux I__6542 (
            .O(N__27224),
            .I(\tok.n297 ));
    CascadeMux I__6541 (
            .O(N__27221),
            .I(N__27218));
    InMux I__6540 (
            .O(N__27218),
            .I(N__27215));
    LocalMux I__6539 (
            .O(N__27215),
            .I(N__27210));
    CascadeMux I__6538 (
            .O(N__27214),
            .I(N__27206));
    InMux I__6537 (
            .O(N__27213),
            .I(N__27203));
    Span4Mux_s3_v I__6536 (
            .O(N__27210),
            .I(N__27200));
    CascadeMux I__6535 (
            .O(N__27209),
            .I(N__27197));
    InMux I__6534 (
            .O(N__27206),
            .I(N__27192));
    LocalMux I__6533 (
            .O(N__27203),
            .I(N__27189));
    Span4Mux_v I__6532 (
            .O(N__27200),
            .I(N__27184));
    InMux I__6531 (
            .O(N__27197),
            .I(N__27181));
    CascadeMux I__6530 (
            .O(N__27196),
            .I(N__27177));
    InMux I__6529 (
            .O(N__27195),
            .I(N__27174));
    LocalMux I__6528 (
            .O(N__27192),
            .I(N__27171));
    Span4Mux_v I__6527 (
            .O(N__27189),
            .I(N__27168));
    InMux I__6526 (
            .O(N__27188),
            .I(N__27165));
    InMux I__6525 (
            .O(N__27187),
            .I(N__27162));
    Span4Mux_h I__6524 (
            .O(N__27184),
            .I(N__27157));
    LocalMux I__6523 (
            .O(N__27181),
            .I(N__27157));
    InMux I__6522 (
            .O(N__27180),
            .I(N__27154));
    InMux I__6521 (
            .O(N__27177),
            .I(N__27151));
    LocalMux I__6520 (
            .O(N__27174),
            .I(N__27146));
    Span4Mux_h I__6519 (
            .O(N__27171),
            .I(N__27146));
    Span4Mux_h I__6518 (
            .O(N__27168),
            .I(N__27141));
    LocalMux I__6517 (
            .O(N__27165),
            .I(N__27141));
    LocalMux I__6516 (
            .O(N__27162),
            .I(N__27136));
    Span4Mux_h I__6515 (
            .O(N__27157),
            .I(N__27136));
    LocalMux I__6514 (
            .O(N__27154),
            .I(\tok.S_5 ));
    LocalMux I__6513 (
            .O(N__27151),
            .I(\tok.S_5 ));
    Odrv4 I__6512 (
            .O(N__27146),
            .I(\tok.S_5 ));
    Odrv4 I__6511 (
            .O(N__27141),
            .I(\tok.S_5 ));
    Odrv4 I__6510 (
            .O(N__27136),
            .I(\tok.S_5 ));
    CascadeMux I__6509 (
            .O(N__27125),
            .I(N__27121));
    InMux I__6508 (
            .O(N__27124),
            .I(N__27116));
    InMux I__6507 (
            .O(N__27121),
            .I(N__27116));
    LocalMux I__6506 (
            .O(N__27116),
            .I(uart_rx_data_5));
    InMux I__6505 (
            .O(N__27113),
            .I(N__27110));
    LocalMux I__6504 (
            .O(N__27110),
            .I(\tok.n6_adj_717 ));
    CascadeMux I__6503 (
            .O(N__27107),
            .I(N__27103));
    CascadeMux I__6502 (
            .O(N__27106),
            .I(N__27100));
    InMux I__6501 (
            .O(N__27103),
            .I(N__27097));
    InMux I__6500 (
            .O(N__27100),
            .I(N__27094));
    LocalMux I__6499 (
            .O(N__27097),
            .I(N__27091));
    LocalMux I__6498 (
            .O(N__27094),
            .I(N__27088));
    Span12Mux_s10_h I__6497 (
            .O(N__27091),
            .I(N__27085));
    Span4Mux_v I__6496 (
            .O(N__27088),
            .I(N__27082));
    Odrv12 I__6495 (
            .O(N__27085),
            .I(\tok.table_rd_5 ));
    Odrv4 I__6494 (
            .O(N__27082),
            .I(\tok.table_rd_5 ));
    InMux I__6493 (
            .O(N__27077),
            .I(N__27074));
    LocalMux I__6492 (
            .O(N__27074),
            .I(\tok.n16_adj_855 ));
    InMux I__6491 (
            .O(N__27071),
            .I(N__27068));
    LocalMux I__6490 (
            .O(N__27068),
            .I(N__27065));
    Span4Mux_v I__6489 (
            .O(N__27065),
            .I(N__27062));
    Span4Mux_h I__6488 (
            .O(N__27062),
            .I(N__27059));
    Odrv4 I__6487 (
            .O(N__27059),
            .I(\tok.n5_adj_800 ));
    InMux I__6486 (
            .O(N__27056),
            .I(N__27053));
    LocalMux I__6485 (
            .O(N__27053),
            .I(N__27050));
    Span4Mux_h I__6484 (
            .O(N__27050),
            .I(N__27047));
    Odrv4 I__6483 (
            .O(N__27047),
            .I(\tok.n10_adj_823 ));
    CascadeMux I__6482 (
            .O(N__27044),
            .I(\tok.n20_adj_857_cascade_ ));
    InMux I__6481 (
            .O(N__27041),
            .I(N__27038));
    LocalMux I__6480 (
            .O(N__27038),
            .I(\tok.n14_adj_856 ));
    InMux I__6479 (
            .O(N__27035),
            .I(N__27032));
    LocalMux I__6478 (
            .O(N__27032),
            .I(N__27029));
    Odrv4 I__6477 (
            .O(N__27029),
            .I(\tok.n5559 ));
    InMux I__6476 (
            .O(N__27026),
            .I(N__27023));
    LocalMux I__6475 (
            .O(N__27023),
            .I(N__27020));
    Span4Mux_s1_h I__6474 (
            .O(N__27020),
            .I(N__27017));
    Span4Mux_h I__6473 (
            .O(N__27017),
            .I(N__27014));
    Odrv4 I__6472 (
            .O(N__27014),
            .I(\tok.n3_adj_859 ));
    CascadeMux I__6471 (
            .O(N__27011),
            .I(\tok.n22_adj_861_cascade_ ));
    InMux I__6470 (
            .O(N__27008),
            .I(N__27005));
    LocalMux I__6469 (
            .O(N__27005),
            .I(\tok.n18_adj_860 ));
    InMux I__6468 (
            .O(N__27002),
            .I(N__26999));
    LocalMux I__6467 (
            .O(N__26999),
            .I(\tok.n5556 ));
    InMux I__6466 (
            .O(N__26996),
            .I(N__26988));
    InMux I__6465 (
            .O(N__26995),
            .I(N__26988));
    InMux I__6464 (
            .O(N__26994),
            .I(N__26985));
    InMux I__6463 (
            .O(N__26993),
            .I(N__26980));
    LocalMux I__6462 (
            .O(N__26988),
            .I(N__26976));
    LocalMux I__6461 (
            .O(N__26985),
            .I(N__26969));
    InMux I__6460 (
            .O(N__26984),
            .I(N__26964));
    InMux I__6459 (
            .O(N__26983),
            .I(N__26964));
    LocalMux I__6458 (
            .O(N__26980),
            .I(N__26961));
    CascadeMux I__6457 (
            .O(N__26979),
            .I(N__26955));
    Span4Mux_s2_h I__6456 (
            .O(N__26976),
            .I(N__26951));
    InMux I__6455 (
            .O(N__26975),
            .I(N__26948));
    InMux I__6454 (
            .O(N__26974),
            .I(N__26941));
    InMux I__6453 (
            .O(N__26973),
            .I(N__26941));
    InMux I__6452 (
            .O(N__26972),
            .I(N__26941));
    Span4Mux_v I__6451 (
            .O(N__26969),
            .I(N__26935));
    LocalMux I__6450 (
            .O(N__26964),
            .I(N__26935));
    Span4Mux_h I__6449 (
            .O(N__26961),
            .I(N__26932));
    InMux I__6448 (
            .O(N__26960),
            .I(N__26927));
    InMux I__6447 (
            .O(N__26959),
            .I(N__26927));
    InMux I__6446 (
            .O(N__26958),
            .I(N__26922));
    InMux I__6445 (
            .O(N__26955),
            .I(N__26922));
    InMux I__6444 (
            .O(N__26954),
            .I(N__26919));
    Span4Mux_h I__6443 (
            .O(N__26951),
            .I(N__26914));
    LocalMux I__6442 (
            .O(N__26948),
            .I(N__26914));
    LocalMux I__6441 (
            .O(N__26941),
            .I(N__26911));
    InMux I__6440 (
            .O(N__26940),
            .I(N__26908));
    Odrv4 I__6439 (
            .O(N__26935),
            .I(\tok.n15 ));
    Odrv4 I__6438 (
            .O(N__26932),
            .I(\tok.n15 ));
    LocalMux I__6437 (
            .O(N__26927),
            .I(\tok.n15 ));
    LocalMux I__6436 (
            .O(N__26922),
            .I(\tok.n15 ));
    LocalMux I__6435 (
            .O(N__26919),
            .I(\tok.n15 ));
    Odrv4 I__6434 (
            .O(N__26914),
            .I(\tok.n15 ));
    Odrv4 I__6433 (
            .O(N__26911),
            .I(\tok.n15 ));
    LocalMux I__6432 (
            .O(N__26908),
            .I(\tok.n15 ));
    InMux I__6431 (
            .O(N__26891),
            .I(N__26888));
    LocalMux I__6430 (
            .O(N__26888),
            .I(N__26885));
    Odrv12 I__6429 (
            .O(N__26885),
            .I(\tok.n5_adj_669 ));
    InMux I__6428 (
            .O(N__26882),
            .I(N__26879));
    LocalMux I__6427 (
            .O(N__26879),
            .I(N__26876));
    Span12Mux_s8_v I__6426 (
            .O(N__26876),
            .I(N__26873));
    Odrv12 I__6425 (
            .O(N__26873),
            .I(\tok.table_rd_8 ));
    CascadeMux I__6424 (
            .O(N__26870),
            .I(N__26865));
    CascadeMux I__6423 (
            .O(N__26869),
            .I(N__26861));
    InMux I__6422 (
            .O(N__26868),
            .I(N__26839));
    InMux I__6421 (
            .O(N__26865),
            .I(N__26839));
    InMux I__6420 (
            .O(N__26864),
            .I(N__26839));
    InMux I__6419 (
            .O(N__26861),
            .I(N__26839));
    InMux I__6418 (
            .O(N__26860),
            .I(N__26839));
    InMux I__6417 (
            .O(N__26859),
            .I(N__26839));
    InMux I__6416 (
            .O(N__26858),
            .I(N__26839));
    InMux I__6415 (
            .O(N__26857),
            .I(N__26830));
    InMux I__6414 (
            .O(N__26856),
            .I(N__26830));
    InMux I__6413 (
            .O(N__26855),
            .I(N__26830));
    InMux I__6412 (
            .O(N__26854),
            .I(N__26830));
    LocalMux I__6411 (
            .O(N__26839),
            .I(N__26824));
    LocalMux I__6410 (
            .O(N__26830),
            .I(N__26821));
    CascadeMux I__6409 (
            .O(N__26829),
            .I(N__26818));
    InMux I__6408 (
            .O(N__26828),
            .I(N__26813));
    InMux I__6407 (
            .O(N__26827),
            .I(N__26813));
    Span4Mux_h I__6406 (
            .O(N__26824),
            .I(N__26808));
    Span4Mux_v I__6405 (
            .O(N__26821),
            .I(N__26808));
    InMux I__6404 (
            .O(N__26818),
            .I(N__26805));
    LocalMux I__6403 (
            .O(N__26813),
            .I(N__26802));
    Span4Mux_h I__6402 (
            .O(N__26808),
            .I(N__26797));
    LocalMux I__6401 (
            .O(N__26805),
            .I(N__26797));
    Span4Mux_h I__6400 (
            .O(N__26802),
            .I(N__26790));
    Span4Mux_v I__6399 (
            .O(N__26797),
            .I(N__26790));
    InMux I__6398 (
            .O(N__26796),
            .I(N__26785));
    InMux I__6397 (
            .O(N__26795),
            .I(N__26785));
    Odrv4 I__6396 (
            .O(N__26790),
            .I(\tok.n4908 ));
    LocalMux I__6395 (
            .O(N__26785),
            .I(\tok.n4908 ));
    InMux I__6394 (
            .O(N__26780),
            .I(N__26777));
    LocalMux I__6393 (
            .O(N__26777),
            .I(N__26774));
    Span4Mux_s2_h I__6392 (
            .O(N__26774),
            .I(N__26771));
    Span4Mux_v I__6391 (
            .O(N__26771),
            .I(N__26768));
    Odrv4 I__6390 (
            .O(N__26768),
            .I(\tok.n181 ));
    InMux I__6389 (
            .O(N__26765),
            .I(N__26757));
    InMux I__6388 (
            .O(N__26764),
            .I(N__26754));
    InMux I__6387 (
            .O(N__26763),
            .I(N__26744));
    InMux I__6386 (
            .O(N__26762),
            .I(N__26741));
    InMux I__6385 (
            .O(N__26761),
            .I(N__26736));
    InMux I__6384 (
            .O(N__26760),
            .I(N__26736));
    LocalMux I__6383 (
            .O(N__26757),
            .I(N__26733));
    LocalMux I__6382 (
            .O(N__26754),
            .I(N__26730));
    InMux I__6381 (
            .O(N__26753),
            .I(N__26727));
    InMux I__6380 (
            .O(N__26752),
            .I(N__26722));
    InMux I__6379 (
            .O(N__26751),
            .I(N__26722));
    InMux I__6378 (
            .O(N__26750),
            .I(N__26719));
    InMux I__6377 (
            .O(N__26749),
            .I(N__26716));
    InMux I__6376 (
            .O(N__26748),
            .I(N__26711));
    InMux I__6375 (
            .O(N__26747),
            .I(N__26711));
    LocalMux I__6374 (
            .O(N__26744),
            .I(N__26707));
    LocalMux I__6373 (
            .O(N__26741),
            .I(N__26704));
    LocalMux I__6372 (
            .O(N__26736),
            .I(N__26699));
    Span4Mux_s3_h I__6371 (
            .O(N__26733),
            .I(N__26699));
    Span4Mux_v I__6370 (
            .O(N__26730),
            .I(N__26694));
    LocalMux I__6369 (
            .O(N__26727),
            .I(N__26694));
    LocalMux I__6368 (
            .O(N__26722),
            .I(N__26685));
    LocalMux I__6367 (
            .O(N__26719),
            .I(N__26685));
    LocalMux I__6366 (
            .O(N__26716),
            .I(N__26685));
    LocalMux I__6365 (
            .O(N__26711),
            .I(N__26685));
    InMux I__6364 (
            .O(N__26710),
            .I(N__26682));
    Span4Mux_h I__6363 (
            .O(N__26707),
            .I(N__26679));
    Span4Mux_h I__6362 (
            .O(N__26704),
            .I(N__26674));
    Span4Mux_h I__6361 (
            .O(N__26699),
            .I(N__26674));
    Span4Mux_h I__6360 (
            .O(N__26694),
            .I(N__26667));
    Span4Mux_v I__6359 (
            .O(N__26685),
            .I(N__26667));
    LocalMux I__6358 (
            .O(N__26682),
            .I(N__26667));
    Odrv4 I__6357 (
            .O(N__26679),
            .I(\tok.n2735 ));
    Odrv4 I__6356 (
            .O(N__26674),
            .I(\tok.n2735 ));
    Odrv4 I__6355 (
            .O(N__26667),
            .I(\tok.n2735 ));
    InMux I__6354 (
            .O(N__26660),
            .I(N__26657));
    LocalMux I__6353 (
            .O(N__26657),
            .I(\tok.n15_adj_670 ));
    CascadeMux I__6352 (
            .O(N__26654),
            .I(\tok.n13_adj_674_cascade_ ));
    InMux I__6351 (
            .O(N__26651),
            .I(N__26648));
    LocalMux I__6350 (
            .O(N__26648),
            .I(\tok.n5416 ));
    InMux I__6349 (
            .O(N__26645),
            .I(N__26639));
    InMux I__6348 (
            .O(N__26644),
            .I(N__26639));
    LocalMux I__6347 (
            .O(N__26639),
            .I(\tok.A_stk.tail_19 ));
    InMux I__6346 (
            .O(N__26636),
            .I(N__26630));
    InMux I__6345 (
            .O(N__26635),
            .I(N__26630));
    LocalMux I__6344 (
            .O(N__26630),
            .I(\tok.A_stk.tail_35 ));
    InMux I__6343 (
            .O(N__26627),
            .I(N__26624));
    LocalMux I__6342 (
            .O(N__26624),
            .I(N__26620));
    InMux I__6341 (
            .O(N__26623),
            .I(N__26617));
    Span4Mux_s3_h I__6340 (
            .O(N__26620),
            .I(N__26614));
    LocalMux I__6339 (
            .O(N__26617),
            .I(N__26611));
    Odrv4 I__6338 (
            .O(N__26614),
            .I(\tok.A_stk.tail_67 ));
    Odrv4 I__6337 (
            .O(N__26611),
            .I(\tok.A_stk.tail_67 ));
    InMux I__6336 (
            .O(N__26606),
            .I(N__26591));
    InMux I__6335 (
            .O(N__26605),
            .I(N__26591));
    InMux I__6334 (
            .O(N__26604),
            .I(N__26591));
    InMux I__6333 (
            .O(N__26603),
            .I(N__26591));
    InMux I__6332 (
            .O(N__26602),
            .I(N__26591));
    LocalMux I__6331 (
            .O(N__26591),
            .I(N__26550));
    InMux I__6330 (
            .O(N__26590),
            .I(N__26541));
    InMux I__6329 (
            .O(N__26589),
            .I(N__26541));
    InMux I__6328 (
            .O(N__26588),
            .I(N__26541));
    InMux I__6327 (
            .O(N__26587),
            .I(N__26541));
    InMux I__6326 (
            .O(N__26586),
            .I(N__26532));
    InMux I__6325 (
            .O(N__26585),
            .I(N__26532));
    InMux I__6324 (
            .O(N__26584),
            .I(N__26532));
    InMux I__6323 (
            .O(N__26583),
            .I(N__26532));
    CascadeMux I__6322 (
            .O(N__26582),
            .I(N__26513));
    InMux I__6321 (
            .O(N__26581),
            .I(N__26503));
    InMux I__6320 (
            .O(N__26580),
            .I(N__26486));
    InMux I__6319 (
            .O(N__26579),
            .I(N__26486));
    InMux I__6318 (
            .O(N__26578),
            .I(N__26486));
    InMux I__6317 (
            .O(N__26577),
            .I(N__26486));
    InMux I__6316 (
            .O(N__26576),
            .I(N__26486));
    InMux I__6315 (
            .O(N__26575),
            .I(N__26486));
    InMux I__6314 (
            .O(N__26574),
            .I(N__26486));
    InMux I__6313 (
            .O(N__26573),
            .I(N__26473));
    InMux I__6312 (
            .O(N__26572),
            .I(N__26473));
    InMux I__6311 (
            .O(N__26571),
            .I(N__26473));
    InMux I__6310 (
            .O(N__26570),
            .I(N__26473));
    InMux I__6309 (
            .O(N__26569),
            .I(N__26473));
    InMux I__6308 (
            .O(N__26568),
            .I(N__26473));
    InMux I__6307 (
            .O(N__26567),
            .I(N__26456));
    InMux I__6306 (
            .O(N__26566),
            .I(N__26456));
    InMux I__6305 (
            .O(N__26565),
            .I(N__26456));
    InMux I__6304 (
            .O(N__26564),
            .I(N__26456));
    InMux I__6303 (
            .O(N__26563),
            .I(N__26456));
    InMux I__6302 (
            .O(N__26562),
            .I(N__26456));
    InMux I__6301 (
            .O(N__26561),
            .I(N__26456));
    InMux I__6300 (
            .O(N__26560),
            .I(N__26456));
    InMux I__6299 (
            .O(N__26559),
            .I(N__26434));
    InMux I__6298 (
            .O(N__26558),
            .I(N__26434));
    InMux I__6297 (
            .O(N__26557),
            .I(N__26434));
    InMux I__6296 (
            .O(N__26556),
            .I(N__26434));
    InMux I__6295 (
            .O(N__26555),
            .I(N__26434));
    InMux I__6294 (
            .O(N__26554),
            .I(N__26434));
    InMux I__6293 (
            .O(N__26553),
            .I(N__26434));
    Span4Mux_v I__6292 (
            .O(N__26550),
            .I(N__26429));
    LocalMux I__6291 (
            .O(N__26541),
            .I(N__26429));
    LocalMux I__6290 (
            .O(N__26532),
            .I(N__26426));
    InMux I__6289 (
            .O(N__26531),
            .I(N__26415));
    InMux I__6288 (
            .O(N__26530),
            .I(N__26415));
    InMux I__6287 (
            .O(N__26529),
            .I(N__26415));
    InMux I__6286 (
            .O(N__26528),
            .I(N__26415));
    InMux I__6285 (
            .O(N__26527),
            .I(N__26415));
    InMux I__6284 (
            .O(N__26526),
            .I(N__26390));
    InMux I__6283 (
            .O(N__26525),
            .I(N__26373));
    InMux I__6282 (
            .O(N__26524),
            .I(N__26373));
    InMux I__6281 (
            .O(N__26523),
            .I(N__26373));
    InMux I__6280 (
            .O(N__26522),
            .I(N__26373));
    InMux I__6279 (
            .O(N__26521),
            .I(N__26373));
    InMux I__6278 (
            .O(N__26520),
            .I(N__26373));
    InMux I__6277 (
            .O(N__26519),
            .I(N__26373));
    InMux I__6276 (
            .O(N__26518),
            .I(N__26373));
    InMux I__6275 (
            .O(N__26517),
            .I(N__26364));
    InMux I__6274 (
            .O(N__26516),
            .I(N__26364));
    InMux I__6273 (
            .O(N__26513),
            .I(N__26364));
    InMux I__6272 (
            .O(N__26512),
            .I(N__26364));
    InMux I__6271 (
            .O(N__26511),
            .I(N__26351));
    InMux I__6270 (
            .O(N__26510),
            .I(N__26351));
    InMux I__6269 (
            .O(N__26509),
            .I(N__26351));
    InMux I__6268 (
            .O(N__26508),
            .I(N__26351));
    InMux I__6267 (
            .O(N__26507),
            .I(N__26351));
    InMux I__6266 (
            .O(N__26506),
            .I(N__26351));
    LocalMux I__6265 (
            .O(N__26503),
            .I(N__26340));
    InMux I__6264 (
            .O(N__26502),
            .I(N__26335));
    InMux I__6263 (
            .O(N__26501),
            .I(N__26335));
    LocalMux I__6262 (
            .O(N__26486),
            .I(N__26332));
    LocalMux I__6261 (
            .O(N__26473),
            .I(N__26327));
    LocalMux I__6260 (
            .O(N__26456),
            .I(N__26327));
    InMux I__6259 (
            .O(N__26455),
            .I(N__26312));
    InMux I__6258 (
            .O(N__26454),
            .I(N__26312));
    InMux I__6257 (
            .O(N__26453),
            .I(N__26312));
    InMux I__6256 (
            .O(N__26452),
            .I(N__26312));
    InMux I__6255 (
            .O(N__26451),
            .I(N__26312));
    InMux I__6254 (
            .O(N__26450),
            .I(N__26312));
    InMux I__6253 (
            .O(N__26449),
            .I(N__26312));
    LocalMux I__6252 (
            .O(N__26434),
            .I(N__26309));
    Span4Mux_v I__6251 (
            .O(N__26429),
            .I(N__26302));
    Span4Mux_s1_h I__6250 (
            .O(N__26426),
            .I(N__26302));
    LocalMux I__6249 (
            .O(N__26415),
            .I(N__26302));
    InMux I__6248 (
            .O(N__26414),
            .I(N__26287));
    InMux I__6247 (
            .O(N__26413),
            .I(N__26287));
    InMux I__6246 (
            .O(N__26412),
            .I(N__26287));
    InMux I__6245 (
            .O(N__26411),
            .I(N__26287));
    InMux I__6244 (
            .O(N__26410),
            .I(N__26287));
    InMux I__6243 (
            .O(N__26409),
            .I(N__26287));
    InMux I__6242 (
            .O(N__26408),
            .I(N__26287));
    InMux I__6241 (
            .O(N__26407),
            .I(N__26264));
    InMux I__6240 (
            .O(N__26406),
            .I(N__26264));
    InMux I__6239 (
            .O(N__26405),
            .I(N__26264));
    InMux I__6238 (
            .O(N__26404),
            .I(N__26264));
    InMux I__6237 (
            .O(N__26403),
            .I(N__26264));
    InMux I__6236 (
            .O(N__26402),
            .I(N__26264));
    InMux I__6235 (
            .O(N__26401),
            .I(N__26264));
    InMux I__6234 (
            .O(N__26400),
            .I(N__26247));
    InMux I__6233 (
            .O(N__26399),
            .I(N__26247));
    InMux I__6232 (
            .O(N__26398),
            .I(N__26247));
    InMux I__6231 (
            .O(N__26397),
            .I(N__26247));
    InMux I__6230 (
            .O(N__26396),
            .I(N__26247));
    InMux I__6229 (
            .O(N__26395),
            .I(N__26247));
    InMux I__6228 (
            .O(N__26394),
            .I(N__26247));
    InMux I__6227 (
            .O(N__26393),
            .I(N__26247));
    LocalMux I__6226 (
            .O(N__26390),
            .I(N__26235));
    LocalMux I__6225 (
            .O(N__26373),
            .I(N__26230));
    LocalMux I__6224 (
            .O(N__26364),
            .I(N__26230));
    LocalMux I__6223 (
            .O(N__26351),
            .I(N__26227));
    InMux I__6222 (
            .O(N__26350),
            .I(N__26210));
    InMux I__6221 (
            .O(N__26349),
            .I(N__26210));
    InMux I__6220 (
            .O(N__26348),
            .I(N__26210));
    InMux I__6219 (
            .O(N__26347),
            .I(N__26210));
    InMux I__6218 (
            .O(N__26346),
            .I(N__26210));
    InMux I__6217 (
            .O(N__26345),
            .I(N__26210));
    InMux I__6216 (
            .O(N__26344),
            .I(N__26210));
    InMux I__6215 (
            .O(N__26343),
            .I(N__26210));
    Span4Mux_s3_v I__6214 (
            .O(N__26340),
            .I(N__26207));
    LocalMux I__6213 (
            .O(N__26335),
            .I(N__26204));
    Span4Mux_s2_v I__6212 (
            .O(N__26332),
            .I(N__26197));
    Span4Mux_s2_h I__6211 (
            .O(N__26327),
            .I(N__26197));
    LocalMux I__6210 (
            .O(N__26312),
            .I(N__26197));
    Span4Mux_s3_v I__6209 (
            .O(N__26309),
            .I(N__26189));
    Span4Mux_h I__6208 (
            .O(N__26302),
            .I(N__26184));
    LocalMux I__6207 (
            .O(N__26287),
            .I(N__26184));
    InMux I__6206 (
            .O(N__26286),
            .I(N__26167));
    InMux I__6205 (
            .O(N__26285),
            .I(N__26167));
    InMux I__6204 (
            .O(N__26284),
            .I(N__26167));
    InMux I__6203 (
            .O(N__26283),
            .I(N__26167));
    InMux I__6202 (
            .O(N__26282),
            .I(N__26167));
    InMux I__6201 (
            .O(N__26281),
            .I(N__26167));
    InMux I__6200 (
            .O(N__26280),
            .I(N__26167));
    InMux I__6199 (
            .O(N__26279),
            .I(N__26167));
    LocalMux I__6198 (
            .O(N__26264),
            .I(N__26162));
    LocalMux I__6197 (
            .O(N__26247),
            .I(N__26162));
    InMux I__6196 (
            .O(N__26246),
            .I(N__26159));
    InMux I__6195 (
            .O(N__26245),
            .I(N__26142));
    InMux I__6194 (
            .O(N__26244),
            .I(N__26142));
    InMux I__6193 (
            .O(N__26243),
            .I(N__26142));
    InMux I__6192 (
            .O(N__26242),
            .I(N__26142));
    InMux I__6191 (
            .O(N__26241),
            .I(N__26142));
    InMux I__6190 (
            .O(N__26240),
            .I(N__26142));
    InMux I__6189 (
            .O(N__26239),
            .I(N__26142));
    InMux I__6188 (
            .O(N__26238),
            .I(N__26142));
    Span4Mux_s3_v I__6187 (
            .O(N__26235),
            .I(N__26129));
    Span4Mux_s3_h I__6186 (
            .O(N__26230),
            .I(N__26129));
    Span4Mux_v I__6185 (
            .O(N__26227),
            .I(N__26129));
    LocalMux I__6184 (
            .O(N__26210),
            .I(N__26129));
    Span4Mux_h I__6183 (
            .O(N__26207),
            .I(N__26129));
    Span4Mux_s3_v I__6182 (
            .O(N__26204),
            .I(N__26129));
    Span4Mux_h I__6181 (
            .O(N__26197),
            .I(N__26126));
    InMux I__6180 (
            .O(N__26196),
            .I(N__26115));
    InMux I__6179 (
            .O(N__26195),
            .I(N__26115));
    InMux I__6178 (
            .O(N__26194),
            .I(N__26115));
    InMux I__6177 (
            .O(N__26193),
            .I(N__26115));
    InMux I__6176 (
            .O(N__26192),
            .I(N__26115));
    Odrv4 I__6175 (
            .O(N__26189),
            .I(A_stk_delta_1));
    Odrv4 I__6174 (
            .O(N__26184),
            .I(A_stk_delta_1));
    LocalMux I__6173 (
            .O(N__26167),
            .I(A_stk_delta_1));
    Odrv4 I__6172 (
            .O(N__26162),
            .I(A_stk_delta_1));
    LocalMux I__6171 (
            .O(N__26159),
            .I(A_stk_delta_1));
    LocalMux I__6170 (
            .O(N__26142),
            .I(A_stk_delta_1));
    Odrv4 I__6169 (
            .O(N__26129),
            .I(A_stk_delta_1));
    Odrv4 I__6168 (
            .O(N__26126),
            .I(A_stk_delta_1));
    LocalMux I__6167 (
            .O(N__26115),
            .I(A_stk_delta_1));
    InMux I__6166 (
            .O(N__26096),
            .I(N__26093));
    LocalMux I__6165 (
            .O(N__26093),
            .I(N__26089));
    InMux I__6164 (
            .O(N__26092),
            .I(N__26086));
    Span12Mux_s5_v I__6163 (
            .O(N__26089),
            .I(N__26083));
    LocalMux I__6162 (
            .O(N__26086),
            .I(\tok.A_stk.tail_51 ));
    Odrv12 I__6161 (
            .O(N__26083),
            .I(\tok.A_stk.tail_51 ));
    CEMux I__6160 (
            .O(N__26078),
            .I(N__26075));
    LocalMux I__6159 (
            .O(N__26075),
            .I(N__26068));
    CEMux I__6158 (
            .O(N__26074),
            .I(N__26065));
    CEMux I__6157 (
            .O(N__26073),
            .I(N__26062));
    CEMux I__6156 (
            .O(N__26072),
            .I(N__26050));
    CEMux I__6155 (
            .O(N__26071),
            .I(N__26044));
    Span4Mux_v I__6154 (
            .O(N__26068),
            .I(N__26039));
    LocalMux I__6153 (
            .O(N__26065),
            .I(N__26039));
    LocalMux I__6152 (
            .O(N__26062),
            .I(N__26036));
    CEMux I__6151 (
            .O(N__26061),
            .I(N__26032));
    CEMux I__6150 (
            .O(N__26060),
            .I(N__26028));
    CEMux I__6149 (
            .O(N__26059),
            .I(N__26025));
    CEMux I__6148 (
            .O(N__26058),
            .I(N__26022));
    InMux I__6147 (
            .O(N__26057),
            .I(N__26016));
    CascadeMux I__6146 (
            .O(N__26056),
            .I(N__26013));
    CascadeMux I__6145 (
            .O(N__26055),
            .I(N__26007));
    CascadeMux I__6144 (
            .O(N__26054),
            .I(N__26003));
    CascadeMux I__6143 (
            .O(N__26053),
            .I(N__26000));
    LocalMux I__6142 (
            .O(N__26050),
            .I(N__25996));
    CEMux I__6141 (
            .O(N__26049),
            .I(N__25993));
    CEMux I__6140 (
            .O(N__26048),
            .I(N__25990));
    CEMux I__6139 (
            .O(N__26047),
            .I(N__25987));
    LocalMux I__6138 (
            .O(N__26044),
            .I(N__25983));
    Span4Mux_v I__6137 (
            .O(N__26039),
            .I(N__25978));
    Span4Mux_s3_v I__6136 (
            .O(N__26036),
            .I(N__25978));
    CEMux I__6135 (
            .O(N__26035),
            .I(N__25975));
    LocalMux I__6134 (
            .O(N__26032),
            .I(N__25972));
    CEMux I__6133 (
            .O(N__26031),
            .I(N__25969));
    LocalMux I__6132 (
            .O(N__26028),
            .I(N__25965));
    LocalMux I__6131 (
            .O(N__26025),
            .I(N__25960));
    LocalMux I__6130 (
            .O(N__26022),
            .I(N__25960));
    CEMux I__6129 (
            .O(N__26021),
            .I(N__25957));
    CEMux I__6128 (
            .O(N__26020),
            .I(N__25954));
    CEMux I__6127 (
            .O(N__26019),
            .I(N__25951));
    LocalMux I__6126 (
            .O(N__26016),
            .I(N__25948));
    InMux I__6125 (
            .O(N__26013),
            .I(N__25943));
    InMux I__6124 (
            .O(N__26012),
            .I(N__25943));
    InMux I__6123 (
            .O(N__26011),
            .I(N__25928));
    InMux I__6122 (
            .O(N__26010),
            .I(N__25928));
    InMux I__6121 (
            .O(N__26007),
            .I(N__25928));
    InMux I__6120 (
            .O(N__26006),
            .I(N__25928));
    InMux I__6119 (
            .O(N__26003),
            .I(N__25928));
    InMux I__6118 (
            .O(N__26000),
            .I(N__25928));
    InMux I__6117 (
            .O(N__25999),
            .I(N__25928));
    Span4Mux_s3_v I__6116 (
            .O(N__25996),
            .I(N__25923));
    LocalMux I__6115 (
            .O(N__25993),
            .I(N__25918));
    LocalMux I__6114 (
            .O(N__25990),
            .I(N__25918));
    LocalMux I__6113 (
            .O(N__25987),
            .I(N__25915));
    CEMux I__6112 (
            .O(N__25986),
            .I(N__25912));
    Span4Mux_s3_v I__6111 (
            .O(N__25983),
            .I(N__25901));
    Span4Mux_s1_h I__6110 (
            .O(N__25978),
            .I(N__25901));
    LocalMux I__6109 (
            .O(N__25975),
            .I(N__25901));
    Span4Mux_s3_v I__6108 (
            .O(N__25972),
            .I(N__25901));
    LocalMux I__6107 (
            .O(N__25969),
            .I(N__25901));
    CEMux I__6106 (
            .O(N__25968),
            .I(N__25898));
    Span4Mux_s2_h I__6105 (
            .O(N__25965),
            .I(N__25889));
    Span4Mux_v I__6104 (
            .O(N__25960),
            .I(N__25889));
    LocalMux I__6103 (
            .O(N__25957),
            .I(N__25889));
    LocalMux I__6102 (
            .O(N__25954),
            .I(N__25889));
    LocalMux I__6101 (
            .O(N__25951),
            .I(N__25886));
    Span4Mux_s3_v I__6100 (
            .O(N__25948),
            .I(N__25883));
    LocalMux I__6099 (
            .O(N__25943),
            .I(N__25880));
    LocalMux I__6098 (
            .O(N__25928),
            .I(N__25877));
    CascadeMux I__6097 (
            .O(N__25927),
            .I(N__25874));
    CascadeMux I__6096 (
            .O(N__25926),
            .I(N__25871));
    Span4Mux_h I__6095 (
            .O(N__25923),
            .I(N__25863));
    Span4Mux_s3_v I__6094 (
            .O(N__25918),
            .I(N__25863));
    Span4Mux_s1_v I__6093 (
            .O(N__25915),
            .I(N__25860));
    LocalMux I__6092 (
            .O(N__25912),
            .I(N__25853));
    Sp12to4 I__6091 (
            .O(N__25901),
            .I(N__25853));
    LocalMux I__6090 (
            .O(N__25898),
            .I(N__25853));
    Span4Mux_h I__6089 (
            .O(N__25889),
            .I(N__25850));
    Span4Mux_s3_v I__6088 (
            .O(N__25886),
            .I(N__25841));
    Span4Mux_h I__6087 (
            .O(N__25883),
            .I(N__25841));
    Span4Mux_s3_v I__6086 (
            .O(N__25880),
            .I(N__25841));
    Span4Mux_s3_v I__6085 (
            .O(N__25877),
            .I(N__25841));
    InMux I__6084 (
            .O(N__25874),
            .I(N__25830));
    InMux I__6083 (
            .O(N__25871),
            .I(N__25830));
    InMux I__6082 (
            .O(N__25870),
            .I(N__25830));
    InMux I__6081 (
            .O(N__25869),
            .I(N__25830));
    InMux I__6080 (
            .O(N__25868),
            .I(N__25830));
    Odrv4 I__6079 (
            .O(N__25863),
            .I(rd_15__N_301));
    Odrv4 I__6078 (
            .O(N__25860),
            .I(rd_15__N_301));
    Odrv12 I__6077 (
            .O(N__25853),
            .I(rd_15__N_301));
    Odrv4 I__6076 (
            .O(N__25850),
            .I(rd_15__N_301));
    Odrv4 I__6075 (
            .O(N__25841),
            .I(rd_15__N_301));
    LocalMux I__6074 (
            .O(N__25830),
            .I(rd_15__N_301));
    InMux I__6073 (
            .O(N__25817),
            .I(N__25814));
    LocalMux I__6072 (
            .O(N__25814),
            .I(\tok.n175 ));
    InMux I__6071 (
            .O(N__25811),
            .I(N__25808));
    LocalMux I__6070 (
            .O(N__25808),
            .I(N__25805));
    Span4Mux_s3_h I__6069 (
            .O(N__25805),
            .I(N__25802));
    Odrv4 I__6068 (
            .O(N__25802),
            .I(\tok.n15_adj_770 ));
    InMux I__6067 (
            .O(N__25799),
            .I(N__25796));
    LocalMux I__6066 (
            .O(N__25796),
            .I(N__25793));
    Span4Mux_s3_h I__6065 (
            .O(N__25793),
            .I(N__25790));
    Span4Mux_v I__6064 (
            .O(N__25790),
            .I(N__25787));
    Odrv4 I__6063 (
            .O(N__25787),
            .I(\tok.n14_adj_769 ));
    CascadeMux I__6062 (
            .O(N__25784),
            .I(\tok.n13_adj_772_cascade_ ));
    InMux I__6061 (
            .O(N__25781),
            .I(N__25778));
    LocalMux I__6060 (
            .O(N__25778),
            .I(\tok.n5412 ));
    CascadeMux I__6059 (
            .O(N__25775),
            .I(\tok.n22_adj_773_cascade_ ));
    CascadeMux I__6058 (
            .O(N__25772),
            .I(N__25768));
    InMux I__6057 (
            .O(N__25771),
            .I(N__25758));
    InMux I__6056 (
            .O(N__25768),
            .I(N__25755));
    InMux I__6055 (
            .O(N__25767),
            .I(N__25752));
    InMux I__6054 (
            .O(N__25766),
            .I(N__25749));
    CascadeMux I__6053 (
            .O(N__25765),
            .I(N__25746));
    CascadeMux I__6052 (
            .O(N__25764),
            .I(N__25743));
    InMux I__6051 (
            .O(N__25763),
            .I(N__25735));
    InMux I__6050 (
            .O(N__25762),
            .I(N__25735));
    InMux I__6049 (
            .O(N__25761),
            .I(N__25735));
    LocalMux I__6048 (
            .O(N__25758),
            .I(N__25732));
    LocalMux I__6047 (
            .O(N__25755),
            .I(N__25727));
    LocalMux I__6046 (
            .O(N__25752),
            .I(N__25727));
    LocalMux I__6045 (
            .O(N__25749),
            .I(N__25724));
    InMux I__6044 (
            .O(N__25746),
            .I(N__25721));
    InMux I__6043 (
            .O(N__25743),
            .I(N__25716));
    InMux I__6042 (
            .O(N__25742),
            .I(N__25716));
    LocalMux I__6041 (
            .O(N__25735),
            .I(N__25713));
    Span4Mux_v I__6040 (
            .O(N__25732),
            .I(N__25708));
    Span4Mux_v I__6039 (
            .O(N__25727),
            .I(N__25708));
    Span12Mux_s5_h I__6038 (
            .O(N__25724),
            .I(N__25703));
    LocalMux I__6037 (
            .O(N__25721),
            .I(N__25703));
    LocalMux I__6036 (
            .O(N__25716),
            .I(\tok.A_14 ));
    Odrv4 I__6035 (
            .O(N__25713),
            .I(\tok.A_14 ));
    Odrv4 I__6034 (
            .O(N__25708),
            .I(\tok.A_14 ));
    Odrv12 I__6033 (
            .O(N__25703),
            .I(\tok.A_14 ));
    InMux I__6032 (
            .O(N__25694),
            .I(N__25689));
    InMux I__6031 (
            .O(N__25693),
            .I(N__25685));
    InMux I__6030 (
            .O(N__25692),
            .I(N__25682));
    LocalMux I__6029 (
            .O(N__25689),
            .I(N__25676));
    InMux I__6028 (
            .O(N__25688),
            .I(N__25673));
    LocalMux I__6027 (
            .O(N__25685),
            .I(N__25668));
    LocalMux I__6026 (
            .O(N__25682),
            .I(N__25668));
    InMux I__6025 (
            .O(N__25681),
            .I(N__25665));
    InMux I__6024 (
            .O(N__25680),
            .I(N__25662));
    InMux I__6023 (
            .O(N__25679),
            .I(N__25657));
    Span4Mux_v I__6022 (
            .O(N__25676),
            .I(N__25652));
    LocalMux I__6021 (
            .O(N__25673),
            .I(N__25652));
    Span4Mux_h I__6020 (
            .O(N__25668),
            .I(N__25645));
    LocalMux I__6019 (
            .O(N__25665),
            .I(N__25645));
    LocalMux I__6018 (
            .O(N__25662),
            .I(N__25645));
    InMux I__6017 (
            .O(N__25661),
            .I(N__25642));
    InMux I__6016 (
            .O(N__25660),
            .I(N__25639));
    LocalMux I__6015 (
            .O(N__25657),
            .I(N__25634));
    Span4Mux_h I__6014 (
            .O(N__25652),
            .I(N__25634));
    Span4Mux_h I__6013 (
            .O(N__25645),
            .I(N__25631));
    LocalMux I__6012 (
            .O(N__25642),
            .I(N__25628));
    LocalMux I__6011 (
            .O(N__25639),
            .I(N__25623));
    Span4Mux_v I__6010 (
            .O(N__25634),
            .I(N__25623));
    Odrv4 I__6009 (
            .O(N__25631),
            .I(rx_data_7__N_511));
    Odrv12 I__6008 (
            .O(N__25628),
            .I(rx_data_7__N_511));
    Odrv4 I__6007 (
            .O(N__25623),
            .I(rx_data_7__N_511));
    InMux I__6006 (
            .O(N__25616),
            .I(N__25612));
    CascadeMux I__6005 (
            .O(N__25615),
            .I(N__25608));
    LocalMux I__6004 (
            .O(N__25612),
            .I(N__25605));
    InMux I__6003 (
            .O(N__25611),
            .I(N__25600));
    InMux I__6002 (
            .O(N__25608),
            .I(N__25600));
    Odrv4 I__6001 (
            .O(N__25605),
            .I(capture_6));
    LocalMux I__6000 (
            .O(N__25600),
            .I(capture_6));
    InMux I__5999 (
            .O(N__25595),
            .I(N__25589));
    InMux I__5998 (
            .O(N__25594),
            .I(N__25589));
    LocalMux I__5997 (
            .O(N__25589),
            .I(\tok.A_stk.tail_11 ));
    InMux I__5996 (
            .O(N__25586),
            .I(N__25580));
    InMux I__5995 (
            .O(N__25585),
            .I(N__25580));
    LocalMux I__5994 (
            .O(N__25580),
            .I(\tok.A_stk.tail_27 ));
    InMux I__5993 (
            .O(N__25577),
            .I(N__25571));
    InMux I__5992 (
            .O(N__25576),
            .I(N__25571));
    LocalMux I__5991 (
            .O(N__25571),
            .I(\tok.A_stk.tail_43 ));
    InMux I__5990 (
            .O(N__25568),
            .I(N__25565));
    LocalMux I__5989 (
            .O(N__25565),
            .I(N__25561));
    InMux I__5988 (
            .O(N__25564),
            .I(N__25558));
    Odrv4 I__5987 (
            .O(N__25561),
            .I(\tok.A_stk.tail_75 ));
    LocalMux I__5986 (
            .O(N__25558),
            .I(\tok.A_stk.tail_75 ));
    InMux I__5985 (
            .O(N__25553),
            .I(N__25550));
    LocalMux I__5984 (
            .O(N__25550),
            .I(N__25546));
    InMux I__5983 (
            .O(N__25549),
            .I(N__25543));
    Span4Mux_h I__5982 (
            .O(N__25546),
            .I(N__25540));
    LocalMux I__5981 (
            .O(N__25543),
            .I(\tok.A_stk.tail_59 ));
    Odrv4 I__5980 (
            .O(N__25540),
            .I(\tok.A_stk.tail_59 ));
    InMux I__5979 (
            .O(N__25535),
            .I(N__25532));
    LocalMux I__5978 (
            .O(N__25532),
            .I(\tok.n20_adj_648 ));
    CascadeMux I__5977 (
            .O(N__25529),
            .I(N__25526));
    InMux I__5976 (
            .O(N__25526),
            .I(N__25523));
    LocalMux I__5975 (
            .O(N__25523),
            .I(N__25520));
    Span4Mux_v I__5974 (
            .O(N__25520),
            .I(N__25517));
    Odrv4 I__5973 (
            .O(N__25517),
            .I(\tok.n299 ));
    InMux I__5972 (
            .O(N__25514),
            .I(N__25508));
    CascadeMux I__5971 (
            .O(N__25513),
            .I(N__25505));
    InMux I__5970 (
            .O(N__25512),
            .I(N__25495));
    InMux I__5969 (
            .O(N__25511),
            .I(N__25492));
    LocalMux I__5968 (
            .O(N__25508),
            .I(N__25489));
    InMux I__5967 (
            .O(N__25505),
            .I(N__25484));
    InMux I__5966 (
            .O(N__25504),
            .I(N__25484));
    InMux I__5965 (
            .O(N__25503),
            .I(N__25479));
    InMux I__5964 (
            .O(N__25502),
            .I(N__25479));
    InMux I__5963 (
            .O(N__25501),
            .I(N__25474));
    InMux I__5962 (
            .O(N__25500),
            .I(N__25474));
    InMux I__5961 (
            .O(N__25499),
            .I(N__25468));
    InMux I__5960 (
            .O(N__25498),
            .I(N__25468));
    LocalMux I__5959 (
            .O(N__25495),
            .I(N__25461));
    LocalMux I__5958 (
            .O(N__25492),
            .I(N__25461));
    Span4Mux_v I__5957 (
            .O(N__25489),
            .I(N__25452));
    LocalMux I__5956 (
            .O(N__25484),
            .I(N__25452));
    LocalMux I__5955 (
            .O(N__25479),
            .I(N__25452));
    LocalMux I__5954 (
            .O(N__25474),
            .I(N__25452));
    InMux I__5953 (
            .O(N__25473),
            .I(N__25447));
    LocalMux I__5952 (
            .O(N__25468),
            .I(N__25444));
    InMux I__5951 (
            .O(N__25467),
            .I(N__25441));
    InMux I__5950 (
            .O(N__25466),
            .I(N__25438));
    Span4Mux_s3_v I__5949 (
            .O(N__25461),
            .I(N__25433));
    Span4Mux_v I__5948 (
            .O(N__25452),
            .I(N__25433));
    InMux I__5947 (
            .O(N__25451),
            .I(N__25430));
    InMux I__5946 (
            .O(N__25450),
            .I(N__25427));
    LocalMux I__5945 (
            .O(N__25447),
            .I(N__25424));
    Span4Mux_v I__5944 (
            .O(N__25444),
            .I(N__25421));
    LocalMux I__5943 (
            .O(N__25441),
            .I(N__25418));
    LocalMux I__5942 (
            .O(N__25438),
            .I(N__25415));
    Sp12to4 I__5941 (
            .O(N__25433),
            .I(N__25408));
    LocalMux I__5940 (
            .O(N__25430),
            .I(N__25408));
    LocalMux I__5939 (
            .O(N__25427),
            .I(N__25408));
    Span4Mux_h I__5938 (
            .O(N__25424),
            .I(N__25399));
    Span4Mux_h I__5937 (
            .O(N__25421),
            .I(N__25399));
    Span4Mux_h I__5936 (
            .O(N__25418),
            .I(N__25399));
    Span4Mux_s1_v I__5935 (
            .O(N__25415),
            .I(N__25399));
    Odrv12 I__5934 (
            .O(N__25408),
            .I(\tok.n238 ));
    Odrv4 I__5933 (
            .O(N__25399),
            .I(\tok.n238 ));
    InMux I__5932 (
            .O(N__25394),
            .I(N__25391));
    LocalMux I__5931 (
            .O(N__25391),
            .I(N__25387));
    InMux I__5930 (
            .O(N__25390),
            .I(N__25384));
    Odrv4 I__5929 (
            .O(N__25387),
            .I(\tok.A_stk.tail_5 ));
    LocalMux I__5928 (
            .O(N__25384),
            .I(\tok.A_stk.tail_5 ));
    CascadeMux I__5927 (
            .O(N__25379),
            .I(N__25376));
    InMux I__5926 (
            .O(N__25376),
            .I(N__25370));
    CascadeMux I__5925 (
            .O(N__25375),
            .I(N__25366));
    InMux I__5924 (
            .O(N__25374),
            .I(N__25363));
    CascadeMux I__5923 (
            .O(N__25373),
            .I(N__25360));
    LocalMux I__5922 (
            .O(N__25370),
            .I(N__25357));
    InMux I__5921 (
            .O(N__25369),
            .I(N__25354));
    InMux I__5920 (
            .O(N__25366),
            .I(N__25351));
    LocalMux I__5919 (
            .O(N__25363),
            .I(N__25348));
    InMux I__5918 (
            .O(N__25360),
            .I(N__25345));
    Span4Mux_v I__5917 (
            .O(N__25357),
            .I(N__25340));
    LocalMux I__5916 (
            .O(N__25354),
            .I(N__25340));
    LocalMux I__5915 (
            .O(N__25351),
            .I(N__25336));
    Span4Mux_v I__5914 (
            .O(N__25348),
            .I(N__25330));
    LocalMux I__5913 (
            .O(N__25345),
            .I(N__25330));
    Span4Mux_h I__5912 (
            .O(N__25340),
            .I(N__25325));
    InMux I__5911 (
            .O(N__25339),
            .I(N__25322));
    Span4Mux_v I__5910 (
            .O(N__25336),
            .I(N__25319));
    InMux I__5909 (
            .O(N__25335),
            .I(N__25316));
    Span4Mux_h I__5908 (
            .O(N__25330),
            .I(N__25313));
    InMux I__5907 (
            .O(N__25329),
            .I(N__25308));
    InMux I__5906 (
            .O(N__25328),
            .I(N__25308));
    Span4Mux_h I__5905 (
            .O(N__25325),
            .I(N__25303));
    LocalMux I__5904 (
            .O(N__25322),
            .I(N__25303));
    Span4Mux_h I__5903 (
            .O(N__25319),
            .I(N__25298));
    LocalMux I__5902 (
            .O(N__25316),
            .I(N__25298));
    Span4Mux_s1_h I__5901 (
            .O(N__25313),
            .I(N__25295));
    LocalMux I__5900 (
            .O(N__25308),
            .I(\tok.S_3 ));
    Odrv4 I__5899 (
            .O(N__25303),
            .I(\tok.S_3 ));
    Odrv4 I__5898 (
            .O(N__25298),
            .I(\tok.S_3 ));
    Odrv4 I__5897 (
            .O(N__25295),
            .I(\tok.S_3 ));
    CascadeMux I__5896 (
            .O(N__25286),
            .I(N__25283));
    InMux I__5895 (
            .O(N__25283),
            .I(N__25277));
    InMux I__5894 (
            .O(N__25282),
            .I(N__25277));
    LocalMux I__5893 (
            .O(N__25277),
            .I(\tok.A_stk.tail_3 ));
    InMux I__5892 (
            .O(N__25274),
            .I(N__25268));
    InMux I__5891 (
            .O(N__25273),
            .I(N__25268));
    LocalMux I__5890 (
            .O(N__25268),
            .I(\tok.A_stk.tail_53 ));
    InMux I__5889 (
            .O(N__25265),
            .I(N__25259));
    InMux I__5888 (
            .O(N__25264),
            .I(N__25259));
    LocalMux I__5887 (
            .O(N__25259),
            .I(\tok.A_stk.tail_37 ));
    InMux I__5886 (
            .O(N__25256),
            .I(N__25250));
    InMux I__5885 (
            .O(N__25255),
            .I(N__25250));
    LocalMux I__5884 (
            .O(N__25250),
            .I(\tok.A_stk.tail_21 ));
    InMux I__5883 (
            .O(N__25247),
            .I(N__25243));
    InMux I__5882 (
            .O(N__25246),
            .I(N__25240));
    LocalMux I__5881 (
            .O(N__25243),
            .I(\tok.A_stk.tail_90 ));
    LocalMux I__5880 (
            .O(N__25240),
            .I(\tok.A_stk.tail_90 ));
    InMux I__5879 (
            .O(N__25235),
            .I(N__25232));
    LocalMux I__5878 (
            .O(N__25232),
            .I(N__25229));
    IoSpan4Mux I__5877 (
            .O(N__25229),
            .I(N__25225));
    CascadeMux I__5876 (
            .O(N__25228),
            .I(N__25222));
    Span4Mux_s1_v I__5875 (
            .O(N__25225),
            .I(N__25219));
    InMux I__5874 (
            .O(N__25222),
            .I(N__25216));
    Odrv4 I__5873 (
            .O(N__25219),
            .I(tail_122));
    LocalMux I__5872 (
            .O(N__25216),
            .I(tail_122));
    InMux I__5871 (
            .O(N__25211),
            .I(N__25208));
    LocalMux I__5870 (
            .O(N__25208),
            .I(N__25204));
    InMux I__5869 (
            .O(N__25207),
            .I(N__25201));
    Span4Mux_h I__5868 (
            .O(N__25204),
            .I(N__25198));
    LocalMux I__5867 (
            .O(N__25201),
            .I(N__25195));
    Odrv4 I__5866 (
            .O(N__25198),
            .I(tail_106));
    Odrv4 I__5865 (
            .O(N__25195),
            .I(tail_106));
    InMux I__5864 (
            .O(N__25190),
            .I(N__25187));
    LocalMux I__5863 (
            .O(N__25187),
            .I(\tok.n23_adj_642 ));
    CascadeMux I__5862 (
            .O(N__25184),
            .I(N__25181));
    InMux I__5861 (
            .O(N__25181),
            .I(N__25178));
    LocalMux I__5860 (
            .O(N__25178),
            .I(N__25175));
    Span4Mux_v I__5859 (
            .O(N__25175),
            .I(N__25172));
    Odrv4 I__5858 (
            .O(N__25172),
            .I(\tok.n288 ));
    InMux I__5857 (
            .O(N__25169),
            .I(N__25161));
    InMux I__5856 (
            .O(N__25168),
            .I(N__25161));
    InMux I__5855 (
            .O(N__25167),
            .I(N__25153));
    InMux I__5854 (
            .O(N__25166),
            .I(N__25150));
    LocalMux I__5853 (
            .O(N__25161),
            .I(N__25147));
    InMux I__5852 (
            .O(N__25160),
            .I(N__25142));
    InMux I__5851 (
            .O(N__25159),
            .I(N__25139));
    InMux I__5850 (
            .O(N__25158),
            .I(N__25136));
    InMux I__5849 (
            .O(N__25157),
            .I(N__25131));
    InMux I__5848 (
            .O(N__25156),
            .I(N__25131));
    LocalMux I__5847 (
            .O(N__25153),
            .I(N__25126));
    LocalMux I__5846 (
            .O(N__25150),
            .I(N__25126));
    Span4Mux_v I__5845 (
            .O(N__25147),
            .I(N__25123));
    InMux I__5844 (
            .O(N__25146),
            .I(N__25120));
    CascadeMux I__5843 (
            .O(N__25145),
            .I(N__25117));
    LocalMux I__5842 (
            .O(N__25142),
            .I(N__25109));
    LocalMux I__5841 (
            .O(N__25139),
            .I(N__25109));
    LocalMux I__5840 (
            .O(N__25136),
            .I(N__25109));
    LocalMux I__5839 (
            .O(N__25131),
            .I(N__25106));
    Span4Mux_s3_v I__5838 (
            .O(N__25126),
            .I(N__25099));
    Span4Mux_h I__5837 (
            .O(N__25123),
            .I(N__25099));
    LocalMux I__5836 (
            .O(N__25120),
            .I(N__25099));
    InMux I__5835 (
            .O(N__25117),
            .I(N__25094));
    InMux I__5834 (
            .O(N__25116),
            .I(N__25094));
    Span4Mux_h I__5833 (
            .O(N__25109),
            .I(N__25091));
    Odrv4 I__5832 (
            .O(N__25106),
            .I(\tok.A_11 ));
    Odrv4 I__5831 (
            .O(N__25099),
            .I(\tok.A_11 ));
    LocalMux I__5830 (
            .O(N__25094),
            .I(\tok.A_11 ));
    Odrv4 I__5829 (
            .O(N__25091),
            .I(\tok.A_11 ));
    InMux I__5828 (
            .O(N__25082),
            .I(N__25079));
    LocalMux I__5827 (
            .O(N__25079),
            .I(N__25076));
    Span4Mux_s1_h I__5826 (
            .O(N__25076),
            .I(N__25073));
    Span4Mux_h I__5825 (
            .O(N__25073),
            .I(N__25069));
    InMux I__5824 (
            .O(N__25072),
            .I(N__25066));
    Odrv4 I__5823 (
            .O(N__25069),
            .I(\tok.A_stk.tail_14 ));
    LocalMux I__5822 (
            .O(N__25066),
            .I(\tok.A_stk.tail_14 ));
    InMux I__5821 (
            .O(N__25061),
            .I(N__25056));
    InMux I__5820 (
            .O(N__25060),
            .I(N__25051));
    CascadeMux I__5819 (
            .O(N__25059),
            .I(N__25048));
    LocalMux I__5818 (
            .O(N__25056),
            .I(N__25045));
    InMux I__5817 (
            .O(N__25055),
            .I(N__25042));
    InMux I__5816 (
            .O(N__25054),
            .I(N__25038));
    LocalMux I__5815 (
            .O(N__25051),
            .I(N__25035));
    InMux I__5814 (
            .O(N__25048),
            .I(N__25032));
    Span4Mux_h I__5813 (
            .O(N__25045),
            .I(N__25027));
    LocalMux I__5812 (
            .O(N__25042),
            .I(N__25027));
    InMux I__5811 (
            .O(N__25041),
            .I(N__25024));
    LocalMux I__5810 (
            .O(N__25038),
            .I(N__25021));
    Span4Mux_v I__5809 (
            .O(N__25035),
            .I(N__25016));
    LocalMux I__5808 (
            .O(N__25032),
            .I(N__25016));
    Span4Mux_h I__5807 (
            .O(N__25027),
            .I(N__25011));
    LocalMux I__5806 (
            .O(N__25024),
            .I(N__25011));
    Span4Mux_v I__5805 (
            .O(N__25021),
            .I(N__25004));
    Span4Mux_h I__5804 (
            .O(N__25016),
            .I(N__25004));
    Span4Mux_v I__5803 (
            .O(N__25011),
            .I(N__25001));
    InMux I__5802 (
            .O(N__25010),
            .I(N__24996));
    InMux I__5801 (
            .O(N__25009),
            .I(N__24996));
    Span4Mux_h I__5800 (
            .O(N__25004),
            .I(N__24993));
    Odrv4 I__5799 (
            .O(N__25001),
            .I(\tok.S_11 ));
    LocalMux I__5798 (
            .O(N__24996),
            .I(\tok.S_11 ));
    Odrv4 I__5797 (
            .O(N__24993),
            .I(\tok.S_11 ));
    CascadeMux I__5796 (
            .O(N__24986),
            .I(N__24983));
    InMux I__5795 (
            .O(N__24983),
            .I(N__24977));
    InMux I__5794 (
            .O(N__24982),
            .I(N__24977));
    LocalMux I__5793 (
            .O(N__24977),
            .I(\tok.A_stk.tail_74 ));
    CascadeMux I__5792 (
            .O(N__24974),
            .I(N__24971));
    InMux I__5791 (
            .O(N__24971),
            .I(N__24965));
    InMux I__5790 (
            .O(N__24970),
            .I(N__24965));
    LocalMux I__5789 (
            .O(N__24965),
            .I(\tok.A_stk.tail_58 ));
    InMux I__5788 (
            .O(N__24962),
            .I(N__24956));
    InMux I__5787 (
            .O(N__24961),
            .I(N__24956));
    LocalMux I__5786 (
            .O(N__24956),
            .I(\tok.A_stk.tail_42 ));
    InMux I__5785 (
            .O(N__24953),
            .I(N__24947));
    InMux I__5784 (
            .O(N__24952),
            .I(N__24947));
    LocalMux I__5783 (
            .O(N__24947),
            .I(\tok.A_stk.tail_26 ));
    CascadeMux I__5782 (
            .O(N__24944),
            .I(N__24941));
    InMux I__5781 (
            .O(N__24941),
            .I(N__24935));
    InMux I__5780 (
            .O(N__24940),
            .I(N__24935));
    LocalMux I__5779 (
            .O(N__24935),
            .I(\tok.A_stk.tail_10 ));
    InMux I__5778 (
            .O(N__24932),
            .I(N__24929));
    LocalMux I__5777 (
            .O(N__24929),
            .I(N__24926));
    Span4Mux_s2_h I__5776 (
            .O(N__24926),
            .I(N__24922));
    InMux I__5775 (
            .O(N__24925),
            .I(N__24919));
    Odrv4 I__5774 (
            .O(N__24922),
            .I(tail_117));
    LocalMux I__5773 (
            .O(N__24919),
            .I(tail_117));
    InMux I__5772 (
            .O(N__24914),
            .I(N__24911));
    LocalMux I__5771 (
            .O(N__24911),
            .I(N__24908));
    Span4Mux_h I__5770 (
            .O(N__24908),
            .I(N__24905));
    Span4Mux_h I__5769 (
            .O(N__24905),
            .I(N__24901));
    InMux I__5768 (
            .O(N__24904),
            .I(N__24898));
    Odrv4 I__5767 (
            .O(N__24901),
            .I(tail_101));
    LocalMux I__5766 (
            .O(N__24898),
            .I(tail_101));
    InMux I__5765 (
            .O(N__24893),
            .I(N__24889));
    InMux I__5764 (
            .O(N__24892),
            .I(N__24886));
    LocalMux I__5763 (
            .O(N__24889),
            .I(\tok.A_stk.tail_85 ));
    LocalMux I__5762 (
            .O(N__24886),
            .I(\tok.A_stk.tail_85 ));
    InMux I__5761 (
            .O(N__24881),
            .I(N__24875));
    InMux I__5760 (
            .O(N__24880),
            .I(N__24875));
    LocalMux I__5759 (
            .O(N__24875),
            .I(\tok.A_stk.tail_69 ));
    CascadeMux I__5758 (
            .O(N__24872),
            .I(N__24869));
    InMux I__5757 (
            .O(N__24869),
            .I(N__24866));
    LocalMux I__5756 (
            .O(N__24866),
            .I(\tok.n287 ));
    InMux I__5755 (
            .O(N__24863),
            .I(N__24857));
    CascadeMux I__5754 (
            .O(N__24862),
            .I(N__24854));
    InMux I__5753 (
            .O(N__24861),
            .I(N__24851));
    InMux I__5752 (
            .O(N__24860),
            .I(N__24848));
    LocalMux I__5751 (
            .O(N__24857),
            .I(N__24840));
    InMux I__5750 (
            .O(N__24854),
            .I(N__24837));
    LocalMux I__5749 (
            .O(N__24851),
            .I(N__24834));
    LocalMux I__5748 (
            .O(N__24848),
            .I(N__24831));
    InMux I__5747 (
            .O(N__24847),
            .I(N__24826));
    InMux I__5746 (
            .O(N__24846),
            .I(N__24826));
    CascadeMux I__5745 (
            .O(N__24845),
            .I(N__24822));
    CascadeMux I__5744 (
            .O(N__24844),
            .I(N__24819));
    InMux I__5743 (
            .O(N__24843),
            .I(N__24816));
    Span4Mux_h I__5742 (
            .O(N__24840),
            .I(N__24811));
    LocalMux I__5741 (
            .O(N__24837),
            .I(N__24811));
    Span4Mux_h I__5740 (
            .O(N__24834),
            .I(N__24804));
    Span4Mux_v I__5739 (
            .O(N__24831),
            .I(N__24804));
    LocalMux I__5738 (
            .O(N__24826),
            .I(N__24804));
    InMux I__5737 (
            .O(N__24825),
            .I(N__24801));
    InMux I__5736 (
            .O(N__24822),
            .I(N__24796));
    InMux I__5735 (
            .O(N__24819),
            .I(N__24796));
    LocalMux I__5734 (
            .O(N__24816),
            .I(N__24791));
    Span4Mux_h I__5733 (
            .O(N__24811),
            .I(N__24791));
    Odrv4 I__5732 (
            .O(N__24804),
            .I(\tok.A_15 ));
    LocalMux I__5731 (
            .O(N__24801),
            .I(\tok.A_15 ));
    LocalMux I__5730 (
            .O(N__24796),
            .I(\tok.A_15 ));
    Odrv4 I__5729 (
            .O(N__24791),
            .I(\tok.A_15 ));
    CascadeMux I__5728 (
            .O(N__24782),
            .I(N__24779));
    InMux I__5727 (
            .O(N__24779),
            .I(N__24774));
    CascadeMux I__5726 (
            .O(N__24778),
            .I(N__24771));
    InMux I__5725 (
            .O(N__24777),
            .I(N__24768));
    LocalMux I__5724 (
            .O(N__24774),
            .I(N__24764));
    InMux I__5723 (
            .O(N__24771),
            .I(N__24761));
    LocalMux I__5722 (
            .O(N__24768),
            .I(N__24755));
    InMux I__5721 (
            .O(N__24767),
            .I(N__24752));
    Span4Mux_h I__5720 (
            .O(N__24764),
            .I(N__24747));
    LocalMux I__5719 (
            .O(N__24761),
            .I(N__24747));
    CascadeMux I__5718 (
            .O(N__24760),
            .I(N__24743));
    InMux I__5717 (
            .O(N__24759),
            .I(N__24738));
    InMux I__5716 (
            .O(N__24758),
            .I(N__24738));
    Span4Mux_h I__5715 (
            .O(N__24755),
            .I(N__24735));
    LocalMux I__5714 (
            .O(N__24752),
            .I(N__24732));
    Span4Mux_h I__5713 (
            .O(N__24747),
            .I(N__24729));
    InMux I__5712 (
            .O(N__24746),
            .I(N__24724));
    InMux I__5711 (
            .O(N__24743),
            .I(N__24724));
    LocalMux I__5710 (
            .O(N__24738),
            .I(N__24719));
    Span4Mux_v I__5709 (
            .O(N__24735),
            .I(N__24719));
    Span4Mux_h I__5708 (
            .O(N__24732),
            .I(N__24714));
    Span4Mux_s1_h I__5707 (
            .O(N__24729),
            .I(N__24714));
    LocalMux I__5706 (
            .O(N__24724),
            .I(N__24711));
    Odrv4 I__5705 (
            .O(N__24719),
            .I(\tok.S_15 ));
    Odrv4 I__5704 (
            .O(N__24714),
            .I(\tok.S_15 ));
    Odrv12 I__5703 (
            .O(N__24711),
            .I(\tok.S_15 ));
    InMux I__5702 (
            .O(N__24704),
            .I(N__24698));
    InMux I__5701 (
            .O(N__24703),
            .I(N__24698));
    LocalMux I__5700 (
            .O(N__24698),
            .I(\tok.A_stk.tail_15 ));
    InMux I__5699 (
            .O(N__24695),
            .I(N__24689));
    InMux I__5698 (
            .O(N__24694),
            .I(N__24689));
    LocalMux I__5697 (
            .O(N__24689),
            .I(\tok.A_stk.tail_31 ));
    InMux I__5696 (
            .O(N__24686),
            .I(N__24680));
    InMux I__5695 (
            .O(N__24685),
            .I(N__24680));
    LocalMux I__5694 (
            .O(N__24680),
            .I(\tok.A_stk.tail_47 ));
    InMux I__5693 (
            .O(N__24677),
            .I(N__24674));
    LocalMux I__5692 (
            .O(N__24674),
            .I(N__24671));
    Span4Mux_v I__5691 (
            .O(N__24671),
            .I(N__24668));
    Span4Mux_v I__5690 (
            .O(N__24668),
            .I(N__24664));
    InMux I__5689 (
            .O(N__24667),
            .I(N__24661));
    Span4Mux_h I__5688 (
            .O(N__24664),
            .I(N__24658));
    LocalMux I__5687 (
            .O(N__24661),
            .I(N__24655));
    Odrv4 I__5686 (
            .O(N__24658),
            .I(\tok.A_stk.tail_95 ));
    Odrv4 I__5685 (
            .O(N__24655),
            .I(\tok.A_stk.tail_95 ));
    InMux I__5684 (
            .O(N__24650),
            .I(N__24644));
    InMux I__5683 (
            .O(N__24649),
            .I(N__24644));
    LocalMux I__5682 (
            .O(N__24644),
            .I(\tok.A_stk.tail_63 ));
    InMux I__5681 (
            .O(N__24641),
            .I(N__24638));
    LocalMux I__5680 (
            .O(N__24638),
            .I(N__24635));
    Span4Mux_h I__5679 (
            .O(N__24635),
            .I(N__24631));
    InMux I__5678 (
            .O(N__24634),
            .I(N__24628));
    Span4Mux_v I__5677 (
            .O(N__24631),
            .I(N__24625));
    LocalMux I__5676 (
            .O(N__24628),
            .I(\tok.A_stk.tail_79 ));
    Odrv4 I__5675 (
            .O(N__24625),
            .I(\tok.A_stk.tail_79 ));
    CascadeMux I__5674 (
            .O(N__24620),
            .I(N__24617));
    InMux I__5673 (
            .O(N__24617),
            .I(N__24614));
    LocalMux I__5672 (
            .O(N__24614),
            .I(N__24611));
    Odrv4 I__5671 (
            .O(N__24611),
            .I(\tok.n293 ));
    InMux I__5670 (
            .O(N__24608),
            .I(N__24605));
    LocalMux I__5669 (
            .O(N__24605),
            .I(N__24602));
    Span4Mux_v I__5668 (
            .O(N__24602),
            .I(N__24599));
    Odrv4 I__5667 (
            .O(N__24599),
            .I(\tok.n28 ));
    InMux I__5666 (
            .O(N__24596),
            .I(\tok.n4777 ));
    InMux I__5665 (
            .O(N__24593),
            .I(N__24585));
    InMux I__5664 (
            .O(N__24592),
            .I(N__24580));
    InMux I__5663 (
            .O(N__24591),
            .I(N__24580));
    InMux I__5662 (
            .O(N__24590),
            .I(N__24577));
    InMux I__5661 (
            .O(N__24589),
            .I(N__24572));
    InMux I__5660 (
            .O(N__24588),
            .I(N__24572));
    LocalMux I__5659 (
            .O(N__24585),
            .I(N__24567));
    LocalMux I__5658 (
            .O(N__24580),
            .I(N__24567));
    LocalMux I__5657 (
            .O(N__24577),
            .I(N__24562));
    LocalMux I__5656 (
            .O(N__24572),
            .I(N__24562));
    Span4Mux_v I__5655 (
            .O(N__24567),
            .I(N__24559));
    Span4Mux_v I__5654 (
            .O(N__24562),
            .I(N__24556));
    Span4Mux_h I__5653 (
            .O(N__24559),
            .I(N__24551));
    Span4Mux_h I__5652 (
            .O(N__24556),
            .I(N__24551));
    Odrv4 I__5651 (
            .O(N__24551),
            .I(\tok.n8_adj_792 ));
    CascadeMux I__5650 (
            .O(N__24548),
            .I(N__24545));
    InMux I__5649 (
            .O(N__24545),
            .I(N__24542));
    LocalMux I__5648 (
            .O(N__24542),
            .I(N__24539));
    Odrv12 I__5647 (
            .O(N__24539),
            .I(\tok.n292 ));
    InMux I__5646 (
            .O(N__24536),
            .I(N__24533));
    LocalMux I__5645 (
            .O(N__24533),
            .I(N__24530));
    Odrv4 I__5644 (
            .O(N__24530),
            .I(\tok.n27_adj_704 ));
    InMux I__5643 (
            .O(N__24527),
            .I(\tok.n4778 ));
    CascadeMux I__5642 (
            .O(N__24524),
            .I(N__24521));
    InMux I__5641 (
            .O(N__24521),
            .I(N__24518));
    LocalMux I__5640 (
            .O(N__24518),
            .I(N__24515));
    Span4Mux_s2_h I__5639 (
            .O(N__24515),
            .I(N__24512));
    Odrv4 I__5638 (
            .O(N__24512),
            .I(\tok.n291 ));
    InMux I__5637 (
            .O(N__24509),
            .I(N__24506));
    LocalMux I__5636 (
            .O(N__24506),
            .I(N__24503));
    Odrv12 I__5635 (
            .O(N__24503),
            .I(\tok.n6_adj_728 ));
    InMux I__5634 (
            .O(N__24500),
            .I(\tok.n4779 ));
    InMux I__5633 (
            .O(N__24497),
            .I(N__24494));
    LocalMux I__5632 (
            .O(N__24494),
            .I(N__24491));
    Odrv12 I__5631 (
            .O(N__24491),
            .I(\tok.n290 ));
    CascadeMux I__5630 (
            .O(N__24488),
            .I(N__24485));
    InMux I__5629 (
            .O(N__24485),
            .I(N__24482));
    LocalMux I__5628 (
            .O(N__24482),
            .I(N__24474));
    InMux I__5627 (
            .O(N__24481),
            .I(N__24471));
    InMux I__5626 (
            .O(N__24480),
            .I(N__24468));
    InMux I__5625 (
            .O(N__24479),
            .I(N__24465));
    CascadeMux I__5624 (
            .O(N__24478),
            .I(N__24461));
    CascadeMux I__5623 (
            .O(N__24477),
            .I(N__24458));
    Span4Mux_h I__5622 (
            .O(N__24474),
            .I(N__24452));
    LocalMux I__5621 (
            .O(N__24471),
            .I(N__24452));
    LocalMux I__5620 (
            .O(N__24468),
            .I(N__24447));
    LocalMux I__5619 (
            .O(N__24465),
            .I(N__24447));
    InMux I__5618 (
            .O(N__24464),
            .I(N__24444));
    InMux I__5617 (
            .O(N__24461),
            .I(N__24441));
    InMux I__5616 (
            .O(N__24458),
            .I(N__24438));
    InMux I__5615 (
            .O(N__24457),
            .I(N__24435));
    Span4Mux_v I__5614 (
            .O(N__24452),
            .I(N__24432));
    Span4Mux_v I__5613 (
            .O(N__24447),
            .I(N__24427));
    LocalMux I__5612 (
            .O(N__24444),
            .I(N__24427));
    LocalMux I__5611 (
            .O(N__24441),
            .I(N__24424));
    LocalMux I__5610 (
            .O(N__24438),
            .I(N__24421));
    LocalMux I__5609 (
            .O(N__24435),
            .I(N__24414));
    Span4Mux_h I__5608 (
            .O(N__24432),
            .I(N__24414));
    Span4Mux_v I__5607 (
            .O(N__24427),
            .I(N__24414));
    Span4Mux_v I__5606 (
            .O(N__24424),
            .I(N__24409));
    Span4Mux_h I__5605 (
            .O(N__24421),
            .I(N__24409));
    Odrv4 I__5604 (
            .O(N__24414),
            .I(\tok.S_12 ));
    Odrv4 I__5603 (
            .O(N__24409),
            .I(\tok.S_12 ));
    InMux I__5602 (
            .O(N__24404),
            .I(N__24401));
    LocalMux I__5601 (
            .O(N__24401),
            .I(N__24398));
    Span4Mux_v I__5600 (
            .O(N__24398),
            .I(N__24395));
    Odrv4 I__5599 (
            .O(N__24395),
            .I(\tok.n6_adj_742 ));
    InMux I__5598 (
            .O(N__24392),
            .I(\tok.n4780 ));
    InMux I__5597 (
            .O(N__24389),
            .I(N__24386));
    LocalMux I__5596 (
            .O(N__24386),
            .I(N__24383));
    Span4Mux_s3_h I__5595 (
            .O(N__24383),
            .I(N__24380));
    Span4Mux_h I__5594 (
            .O(N__24380),
            .I(N__24377));
    Odrv4 I__5593 (
            .O(N__24377),
            .I(\tok.n289 ));
    CascadeMux I__5592 (
            .O(N__24374),
            .I(N__24371));
    InMux I__5591 (
            .O(N__24371),
            .I(N__24366));
    InMux I__5590 (
            .O(N__24370),
            .I(N__24361));
    CascadeMux I__5589 (
            .O(N__24369),
            .I(N__24358));
    LocalMux I__5588 (
            .O(N__24366),
            .I(N__24355));
    InMux I__5587 (
            .O(N__24365),
            .I(N__24352));
    CascadeMux I__5586 (
            .O(N__24364),
            .I(N__24348));
    LocalMux I__5585 (
            .O(N__24361),
            .I(N__24345));
    InMux I__5584 (
            .O(N__24358),
            .I(N__24342));
    Span4Mux_h I__5583 (
            .O(N__24355),
            .I(N__24338));
    LocalMux I__5582 (
            .O(N__24352),
            .I(N__24335));
    InMux I__5581 (
            .O(N__24351),
            .I(N__24332));
    InMux I__5580 (
            .O(N__24348),
            .I(N__24329));
    Span4Mux_h I__5579 (
            .O(N__24345),
            .I(N__24326));
    LocalMux I__5578 (
            .O(N__24342),
            .I(N__24323));
    CascadeMux I__5577 (
            .O(N__24341),
            .I(N__24320));
    Span4Mux_v I__5576 (
            .O(N__24338),
            .I(N__24314));
    Span4Mux_h I__5575 (
            .O(N__24335),
            .I(N__24314));
    LocalMux I__5574 (
            .O(N__24332),
            .I(N__24311));
    LocalMux I__5573 (
            .O(N__24329),
            .I(N__24308));
    Span4Mux_v I__5572 (
            .O(N__24326),
            .I(N__24303));
    Span4Mux_h I__5571 (
            .O(N__24323),
            .I(N__24303));
    InMux I__5570 (
            .O(N__24320),
            .I(N__24300));
    InMux I__5569 (
            .O(N__24319),
            .I(N__24297));
    Span4Mux_v I__5568 (
            .O(N__24314),
            .I(N__24294));
    Span12Mux_s11_h I__5567 (
            .O(N__24311),
            .I(N__24285));
    Span12Mux_s5_v I__5566 (
            .O(N__24308),
            .I(N__24285));
    Sp12to4 I__5565 (
            .O(N__24303),
            .I(N__24285));
    LocalMux I__5564 (
            .O(N__24300),
            .I(N__24285));
    LocalMux I__5563 (
            .O(N__24297),
            .I(\tok.S_13 ));
    Odrv4 I__5562 (
            .O(N__24294),
            .I(\tok.S_13 ));
    Odrv12 I__5561 (
            .O(N__24285),
            .I(\tok.S_13 ));
    InMux I__5560 (
            .O(N__24278),
            .I(N__24275));
    LocalMux I__5559 (
            .O(N__24275),
            .I(N__24272));
    Span4Mux_h I__5558 (
            .O(N__24272),
            .I(N__24269));
    Odrv4 I__5557 (
            .O(N__24269),
            .I(\tok.n6_adj_752 ));
    InMux I__5556 (
            .O(N__24266),
            .I(\tok.n4781 ));
    InMux I__5555 (
            .O(N__24263),
            .I(\tok.n4782 ));
    SRMux I__5554 (
            .O(N__24260),
            .I(N__24255));
    DummyBuf I__5553 (
            .O(N__24259),
            .I(N__24251));
    DummyBuf I__5552 (
            .O(N__24258),
            .I(N__24248));
    LocalMux I__5551 (
            .O(N__24255),
            .I(N__24244));
    SRMux I__5550 (
            .O(N__24254),
            .I(N__24241));
    InMux I__5549 (
            .O(N__24251),
            .I(N__24238));
    InMux I__5548 (
            .O(N__24248),
            .I(N__24235));
    SRMux I__5547 (
            .O(N__24247),
            .I(N__24232));
    Span4Mux_v I__5546 (
            .O(N__24244),
            .I(N__24227));
    LocalMux I__5545 (
            .O(N__24241),
            .I(N__24227));
    LocalMux I__5544 (
            .O(N__24238),
            .I(N__24221));
    LocalMux I__5543 (
            .O(N__24235),
            .I(N__24221));
    LocalMux I__5542 (
            .O(N__24232),
            .I(N__24216));
    Span4Mux_h I__5541 (
            .O(N__24227),
            .I(N__24213));
    InMux I__5540 (
            .O(N__24226),
            .I(N__24210));
    Span4Mux_h I__5539 (
            .O(N__24221),
            .I(N__24206));
    CascadeMux I__5538 (
            .O(N__24220),
            .I(N__24203));
    CascadeMux I__5537 (
            .O(N__24219),
            .I(N__24200));
    Span4Mux_h I__5536 (
            .O(N__24216),
            .I(N__24197));
    Span4Mux_v I__5535 (
            .O(N__24213),
            .I(N__24194));
    LocalMux I__5534 (
            .O(N__24210),
            .I(N__24191));
    CascadeMux I__5533 (
            .O(N__24209),
            .I(N__24186));
    Sp12to4 I__5532 (
            .O(N__24206),
            .I(N__24183));
    InMux I__5531 (
            .O(N__24203),
            .I(N__24178));
    InMux I__5530 (
            .O(N__24200),
            .I(N__24178));
    Span4Mux_h I__5529 (
            .O(N__24197),
            .I(N__24175));
    Span4Mux_s1_v I__5528 (
            .O(N__24194),
            .I(N__24170));
    Span4Mux_v I__5527 (
            .O(N__24191),
            .I(N__24170));
    InMux I__5526 (
            .O(N__24190),
            .I(N__24167));
    InMux I__5525 (
            .O(N__24189),
            .I(N__24164));
    InMux I__5524 (
            .O(N__24186),
            .I(N__24161));
    Span12Mux_v I__5523 (
            .O(N__24183),
            .I(N__24156));
    LocalMux I__5522 (
            .O(N__24178),
            .I(N__24156));
    Odrv4 I__5521 (
            .O(N__24175),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5520 (
            .O(N__24170),
            .I(CONSTANT_ONE_NET));
    LocalMux I__5519 (
            .O(N__24167),
            .I(CONSTANT_ONE_NET));
    LocalMux I__5518 (
            .O(N__24164),
            .I(CONSTANT_ONE_NET));
    LocalMux I__5517 (
            .O(N__24161),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__5516 (
            .O(N__24156),
            .I(CONSTANT_ONE_NET));
    InMux I__5515 (
            .O(N__24143),
            .I(N__24131));
    InMux I__5514 (
            .O(N__24142),
            .I(N__24126));
    InMux I__5513 (
            .O(N__24141),
            .I(N__24126));
    InMux I__5512 (
            .O(N__24140),
            .I(N__24119));
    InMux I__5511 (
            .O(N__24139),
            .I(N__24119));
    InMux I__5510 (
            .O(N__24138),
            .I(N__24119));
    InMux I__5509 (
            .O(N__24137),
            .I(N__24114));
    InMux I__5508 (
            .O(N__24136),
            .I(N__24114));
    InMux I__5507 (
            .O(N__24135),
            .I(N__24109));
    InMux I__5506 (
            .O(N__24134),
            .I(N__24109));
    LocalMux I__5505 (
            .O(N__24131),
            .I(N__24106));
    LocalMux I__5504 (
            .O(N__24126),
            .I(N__24103));
    LocalMux I__5503 (
            .O(N__24119),
            .I(N__24098));
    LocalMux I__5502 (
            .O(N__24114),
            .I(N__24098));
    LocalMux I__5501 (
            .O(N__24109),
            .I(N__24095));
    Span4Mux_v I__5500 (
            .O(N__24106),
            .I(N__24090));
    Span4Mux_v I__5499 (
            .O(N__24103),
            .I(N__24090));
    Span4Mux_s3_h I__5498 (
            .O(N__24098),
            .I(N__24087));
    Sp12to4 I__5497 (
            .O(N__24095),
            .I(N__24082));
    Sp12to4 I__5496 (
            .O(N__24090),
            .I(N__24082));
    Span4Mux_h I__5495 (
            .O(N__24087),
            .I(N__24079));
    Odrv12 I__5494 (
            .O(N__24082),
            .I(\tok.n400 ));
    Odrv4 I__5493 (
            .O(N__24079),
            .I(\tok.n400 ));
    InMux I__5492 (
            .O(N__24074),
            .I(bfn_11_11_0_));
    InMux I__5491 (
            .O(N__24071),
            .I(N__24068));
    LocalMux I__5490 (
            .O(N__24068),
            .I(N__24065));
    Span4Mux_h I__5489 (
            .O(N__24065),
            .I(N__24062));
    Odrv4 I__5488 (
            .O(N__24062),
            .I(\tok.n6_adj_783 ));
    InMux I__5487 (
            .O(N__24059),
            .I(N__24056));
    LocalMux I__5486 (
            .O(N__24056),
            .I(N__24053));
    Odrv12 I__5485 (
            .O(N__24053),
            .I(\tok.n301 ));
    CascadeMux I__5484 (
            .O(N__24050),
            .I(N__24047));
    InMux I__5483 (
            .O(N__24047),
            .I(N__24044));
    LocalMux I__5482 (
            .O(N__24044),
            .I(N__24040));
    CascadeMux I__5481 (
            .O(N__24043),
            .I(N__24036));
    Span4Mux_v I__5480 (
            .O(N__24040),
            .I(N__24032));
    InMux I__5479 (
            .O(N__24039),
            .I(N__24025));
    InMux I__5478 (
            .O(N__24036),
            .I(N__24022));
    CascadeMux I__5477 (
            .O(N__24035),
            .I(N__24019));
    Span4Mux_s3_h I__5476 (
            .O(N__24032),
            .I(N__24016));
    InMux I__5475 (
            .O(N__24031),
            .I(N__24011));
    InMux I__5474 (
            .O(N__24030),
            .I(N__24011));
    InMux I__5473 (
            .O(N__24029),
            .I(N__24008));
    CascadeMux I__5472 (
            .O(N__24028),
            .I(N__24005));
    LocalMux I__5471 (
            .O(N__24025),
            .I(N__24000));
    LocalMux I__5470 (
            .O(N__24022),
            .I(N__24000));
    InMux I__5469 (
            .O(N__24019),
            .I(N__23997));
    Span4Mux_h I__5468 (
            .O(N__24016),
            .I(N__23992));
    LocalMux I__5467 (
            .O(N__24011),
            .I(N__23992));
    LocalMux I__5466 (
            .O(N__24008),
            .I(N__23989));
    InMux I__5465 (
            .O(N__24005),
            .I(N__23986));
    Span4Mux_h I__5464 (
            .O(N__24000),
            .I(N__23981));
    LocalMux I__5463 (
            .O(N__23997),
            .I(N__23981));
    Span4Mux_v I__5462 (
            .O(N__23992),
            .I(N__23975));
    Span4Mux_h I__5461 (
            .O(N__23989),
            .I(N__23975));
    LocalMux I__5460 (
            .O(N__23986),
            .I(N__23972));
    Span4Mux_v I__5459 (
            .O(N__23981),
            .I(N__23969));
    InMux I__5458 (
            .O(N__23980),
            .I(N__23966));
    Span4Mux_v I__5457 (
            .O(N__23975),
            .I(N__23963));
    Span4Mux_v I__5456 (
            .O(N__23972),
            .I(N__23958));
    Span4Mux_h I__5455 (
            .O(N__23969),
            .I(N__23958));
    LocalMux I__5454 (
            .O(N__23966),
            .I(\tok.S_1 ));
    Odrv4 I__5453 (
            .O(N__23963),
            .I(\tok.S_1 ));
    Odrv4 I__5452 (
            .O(N__23958),
            .I(\tok.S_1 ));
    InMux I__5451 (
            .O(N__23951),
            .I(N__23948));
    LocalMux I__5450 (
            .O(N__23948),
            .I(N__23945));
    Odrv4 I__5449 (
            .O(N__23945),
            .I(\tok.n20_adj_799 ));
    InMux I__5448 (
            .O(N__23942),
            .I(\tok.n4769 ));
    CascadeMux I__5447 (
            .O(N__23939),
            .I(N__23936));
    InMux I__5446 (
            .O(N__23936),
            .I(N__23933));
    LocalMux I__5445 (
            .O(N__23933),
            .I(N__23928));
    InMux I__5444 (
            .O(N__23932),
            .I(N__23925));
    InMux I__5443 (
            .O(N__23931),
            .I(N__23921));
    Span4Mux_h I__5442 (
            .O(N__23928),
            .I(N__23917));
    LocalMux I__5441 (
            .O(N__23925),
            .I(N__23914));
    InMux I__5440 (
            .O(N__23924),
            .I(N__23910));
    LocalMux I__5439 (
            .O(N__23921),
            .I(N__23907));
    CascadeMux I__5438 (
            .O(N__23920),
            .I(N__23903));
    Span4Mux_h I__5437 (
            .O(N__23917),
            .I(N__23900));
    Span4Mux_h I__5436 (
            .O(N__23914),
            .I(N__23897));
    InMux I__5435 (
            .O(N__23913),
            .I(N__23894));
    LocalMux I__5434 (
            .O(N__23910),
            .I(N__23891));
    Span4Mux_s3_v I__5433 (
            .O(N__23907),
            .I(N__23888));
    InMux I__5432 (
            .O(N__23906),
            .I(N__23885));
    InMux I__5431 (
            .O(N__23903),
            .I(N__23882));
    Span4Mux_v I__5430 (
            .O(N__23900),
            .I(N__23873));
    Span4Mux_h I__5429 (
            .O(N__23897),
            .I(N__23873));
    LocalMux I__5428 (
            .O(N__23894),
            .I(N__23873));
    Span4Mux_v I__5427 (
            .O(N__23891),
            .I(N__23870));
    Span4Mux_h I__5426 (
            .O(N__23888),
            .I(N__23865));
    LocalMux I__5425 (
            .O(N__23885),
            .I(N__23865));
    LocalMux I__5424 (
            .O(N__23882),
            .I(N__23862));
    InMux I__5423 (
            .O(N__23881),
            .I(N__23857));
    InMux I__5422 (
            .O(N__23880),
            .I(N__23857));
    Span4Mux_v I__5421 (
            .O(N__23873),
            .I(N__23854));
    Span4Mux_h I__5420 (
            .O(N__23870),
            .I(N__23847));
    Span4Mux_v I__5419 (
            .O(N__23865),
            .I(N__23847));
    Span4Mux_h I__5418 (
            .O(N__23862),
            .I(N__23847));
    LocalMux I__5417 (
            .O(N__23857),
            .I(\tok.S_2 ));
    Odrv4 I__5416 (
            .O(N__23854),
            .I(\tok.S_2 ));
    Odrv4 I__5415 (
            .O(N__23847),
            .I(\tok.S_2 ));
    CascadeMux I__5414 (
            .O(N__23840),
            .I(N__23837));
    InMux I__5413 (
            .O(N__23837),
            .I(N__23834));
    LocalMux I__5412 (
            .O(N__23834),
            .I(N__23831));
    Span4Mux_s3_h I__5411 (
            .O(N__23831),
            .I(N__23828));
    Odrv4 I__5410 (
            .O(N__23828),
            .I(\tok.n300 ));
    InMux I__5409 (
            .O(N__23825),
            .I(N__23822));
    LocalMux I__5408 (
            .O(N__23822),
            .I(N__23819));
    Odrv4 I__5407 (
            .O(N__23819),
            .I(\tok.n22_adj_797 ));
    InMux I__5406 (
            .O(N__23816),
            .I(\tok.n4770 ));
    InMux I__5405 (
            .O(N__23813),
            .I(N__23810));
    LocalMux I__5404 (
            .O(N__23810),
            .I(N__23807));
    Span4Mux_h I__5403 (
            .O(N__23807),
            .I(N__23804));
    Span4Mux_h I__5402 (
            .O(N__23804),
            .I(N__23801));
    Odrv4 I__5401 (
            .O(N__23801),
            .I(\tok.n10_adj_791 ));
    InMux I__5400 (
            .O(N__23798),
            .I(\tok.n4771 ));
    CascadeMux I__5399 (
            .O(N__23795),
            .I(N__23789));
    CascadeMux I__5398 (
            .O(N__23794),
            .I(N__23786));
    InMux I__5397 (
            .O(N__23793),
            .I(N__23783));
    CascadeMux I__5396 (
            .O(N__23792),
            .I(N__23780));
    InMux I__5395 (
            .O(N__23789),
            .I(N__23777));
    InMux I__5394 (
            .O(N__23786),
            .I(N__23772));
    LocalMux I__5393 (
            .O(N__23783),
            .I(N__23769));
    InMux I__5392 (
            .O(N__23780),
            .I(N__23766));
    LocalMux I__5391 (
            .O(N__23777),
            .I(N__23763));
    InMux I__5390 (
            .O(N__23776),
            .I(N__23759));
    InMux I__5389 (
            .O(N__23775),
            .I(N__23756));
    LocalMux I__5388 (
            .O(N__23772),
            .I(N__23749));
    Span4Mux_v I__5387 (
            .O(N__23769),
            .I(N__23749));
    LocalMux I__5386 (
            .O(N__23766),
            .I(N__23749));
    Span4Mux_h I__5385 (
            .O(N__23763),
            .I(N__23746));
    CascadeMux I__5384 (
            .O(N__23762),
            .I(N__23743));
    LocalMux I__5383 (
            .O(N__23759),
            .I(N__23739));
    LocalMux I__5382 (
            .O(N__23756),
            .I(N__23736));
    Span4Mux_h I__5381 (
            .O(N__23749),
            .I(N__23733));
    Span4Mux_h I__5380 (
            .O(N__23746),
            .I(N__23729));
    InMux I__5379 (
            .O(N__23743),
            .I(N__23726));
    InMux I__5378 (
            .O(N__23742),
            .I(N__23723));
    Span4Mux_v I__5377 (
            .O(N__23739),
            .I(N__23718));
    Span4Mux_v I__5376 (
            .O(N__23736),
            .I(N__23718));
    Span4Mux_v I__5375 (
            .O(N__23733),
            .I(N__23715));
    InMux I__5374 (
            .O(N__23732),
            .I(N__23712));
    Span4Mux_v I__5373 (
            .O(N__23729),
            .I(N__23707));
    LocalMux I__5372 (
            .O(N__23726),
            .I(N__23707));
    LocalMux I__5371 (
            .O(N__23723),
            .I(\tok.S_4 ));
    Odrv4 I__5370 (
            .O(N__23718),
            .I(\tok.S_4 ));
    Odrv4 I__5369 (
            .O(N__23715),
            .I(\tok.S_4 ));
    LocalMux I__5368 (
            .O(N__23712),
            .I(\tok.S_4 ));
    Odrv4 I__5367 (
            .O(N__23707),
            .I(\tok.S_4 ));
    InMux I__5366 (
            .O(N__23696),
            .I(N__23693));
    LocalMux I__5365 (
            .O(N__23693),
            .I(N__23690));
    Span4Mux_h I__5364 (
            .O(N__23690),
            .I(N__23687));
    Odrv4 I__5363 (
            .O(N__23687),
            .I(\tok.n6_adj_762 ));
    InMux I__5362 (
            .O(N__23684),
            .I(\tok.n4772 ));
    InMux I__5361 (
            .O(N__23681),
            .I(\tok.n4773 ));
    CascadeMux I__5360 (
            .O(N__23678),
            .I(N__23674));
    CascadeMux I__5359 (
            .O(N__23677),
            .I(N__23671));
    InMux I__5358 (
            .O(N__23674),
            .I(N__23668));
    InMux I__5357 (
            .O(N__23671),
            .I(N__23661));
    LocalMux I__5356 (
            .O(N__23668),
            .I(N__23658));
    InMux I__5355 (
            .O(N__23667),
            .I(N__23655));
    CascadeMux I__5354 (
            .O(N__23666),
            .I(N__23652));
    InMux I__5353 (
            .O(N__23665),
            .I(N__23649));
    InMux I__5352 (
            .O(N__23664),
            .I(N__23645));
    LocalMux I__5351 (
            .O(N__23661),
            .I(N__23642));
    Span4Mux_v I__5350 (
            .O(N__23658),
            .I(N__23637));
    LocalMux I__5349 (
            .O(N__23655),
            .I(N__23637));
    InMux I__5348 (
            .O(N__23652),
            .I(N__23634));
    LocalMux I__5347 (
            .O(N__23649),
            .I(N__23630));
    InMux I__5346 (
            .O(N__23648),
            .I(N__23626));
    LocalMux I__5345 (
            .O(N__23645),
            .I(N__23623));
    Span4Mux_v I__5344 (
            .O(N__23642),
            .I(N__23620));
    Span4Mux_h I__5343 (
            .O(N__23637),
            .I(N__23615));
    LocalMux I__5342 (
            .O(N__23634),
            .I(N__23615));
    InMux I__5341 (
            .O(N__23633),
            .I(N__23612));
    Span4Mux_h I__5340 (
            .O(N__23630),
            .I(N__23609));
    InMux I__5339 (
            .O(N__23629),
            .I(N__23606));
    LocalMux I__5338 (
            .O(N__23626),
            .I(N__23597));
    Span4Mux_v I__5337 (
            .O(N__23623),
            .I(N__23597));
    Span4Mux_s1_h I__5336 (
            .O(N__23620),
            .I(N__23597));
    Span4Mux_v I__5335 (
            .O(N__23615),
            .I(N__23597));
    LocalMux I__5334 (
            .O(N__23612),
            .I(\tok.S_6 ));
    Odrv4 I__5333 (
            .O(N__23609),
            .I(\tok.S_6 ));
    LocalMux I__5332 (
            .O(N__23606),
            .I(\tok.S_6 ));
    Odrv4 I__5331 (
            .O(N__23597),
            .I(\tok.S_6 ));
    CascadeMux I__5330 (
            .O(N__23588),
            .I(N__23585));
    InMux I__5329 (
            .O(N__23585),
            .I(N__23582));
    LocalMux I__5328 (
            .O(N__23582),
            .I(N__23579));
    Span4Mux_v I__5327 (
            .O(N__23579),
            .I(N__23576));
    Odrv4 I__5326 (
            .O(N__23576),
            .I(\tok.n296 ));
    InMux I__5325 (
            .O(N__23573),
            .I(N__23570));
    LocalMux I__5324 (
            .O(N__23570),
            .I(N__23567));
    Span4Mux_h I__5323 (
            .O(N__23567),
            .I(N__23564));
    Odrv4 I__5322 (
            .O(N__23564),
            .I(\tok.n6 ));
    InMux I__5321 (
            .O(N__23561),
            .I(\tok.n4774 ));
    CascadeMux I__5320 (
            .O(N__23558),
            .I(N__23555));
    InMux I__5319 (
            .O(N__23555),
            .I(N__23550));
    CascadeMux I__5318 (
            .O(N__23554),
            .I(N__23547));
    CascadeMux I__5317 (
            .O(N__23553),
            .I(N__23544));
    LocalMux I__5316 (
            .O(N__23550),
            .I(N__23540));
    InMux I__5315 (
            .O(N__23547),
            .I(N__23537));
    InMux I__5314 (
            .O(N__23544),
            .I(N__23534));
    InMux I__5313 (
            .O(N__23543),
            .I(N__23530));
    Span4Mux_s3_v I__5312 (
            .O(N__23540),
            .I(N__23527));
    LocalMux I__5311 (
            .O(N__23537),
            .I(N__23524));
    LocalMux I__5310 (
            .O(N__23534),
            .I(N__23520));
    CascadeMux I__5309 (
            .O(N__23533),
            .I(N__23516));
    LocalMux I__5308 (
            .O(N__23530),
            .I(N__23513));
    Span4Mux_h I__5307 (
            .O(N__23527),
            .I(N__23508));
    Span4Mux_s3_v I__5306 (
            .O(N__23524),
            .I(N__23508));
    InMux I__5305 (
            .O(N__23523),
            .I(N__23503));
    Span4Mux_h I__5304 (
            .O(N__23520),
            .I(N__23500));
    InMux I__5303 (
            .O(N__23519),
            .I(N__23497));
    InMux I__5302 (
            .O(N__23516),
            .I(N__23494));
    Span4Mux_v I__5301 (
            .O(N__23513),
            .I(N__23491));
    Span4Mux_h I__5300 (
            .O(N__23508),
            .I(N__23488));
    CascadeMux I__5299 (
            .O(N__23507),
            .I(N__23485));
    InMux I__5298 (
            .O(N__23506),
            .I(N__23482));
    LocalMux I__5297 (
            .O(N__23503),
            .I(N__23475));
    Span4Mux_h I__5296 (
            .O(N__23500),
            .I(N__23475));
    LocalMux I__5295 (
            .O(N__23497),
            .I(N__23475));
    LocalMux I__5294 (
            .O(N__23494),
            .I(N__23472));
    Span4Mux_h I__5293 (
            .O(N__23491),
            .I(N__23467));
    Span4Mux_v I__5292 (
            .O(N__23488),
            .I(N__23467));
    InMux I__5291 (
            .O(N__23485),
            .I(N__23464));
    LocalMux I__5290 (
            .O(N__23482),
            .I(N__23461));
    Span4Mux_v I__5289 (
            .O(N__23475),
            .I(N__23458));
    Span12Mux_s11_h I__5288 (
            .O(N__23472),
            .I(N__23455));
    Odrv4 I__5287 (
            .O(N__23467),
            .I(\tok.S_7 ));
    LocalMux I__5286 (
            .O(N__23464),
            .I(\tok.S_7 ));
    Odrv12 I__5285 (
            .O(N__23461),
            .I(\tok.S_7 ));
    Odrv4 I__5284 (
            .O(N__23458),
            .I(\tok.S_7 ));
    Odrv12 I__5283 (
            .O(N__23455),
            .I(\tok.S_7 ));
    CascadeMux I__5282 (
            .O(N__23444),
            .I(N__23441));
    InMux I__5281 (
            .O(N__23441),
            .I(N__23438));
    LocalMux I__5280 (
            .O(N__23438),
            .I(N__23435));
    Odrv12 I__5279 (
            .O(N__23435),
            .I(\tok.n295 ));
    InMux I__5278 (
            .O(N__23432),
            .I(N__23429));
    LocalMux I__5277 (
            .O(N__23429),
            .I(N__23426));
    Span4Mux_h I__5276 (
            .O(N__23426),
            .I(N__23423));
    Span4Mux_v I__5275 (
            .O(N__23423),
            .I(N__23420));
    Odrv4 I__5274 (
            .O(N__23420),
            .I(\tok.n6_adj_657 ));
    InMux I__5273 (
            .O(N__23417),
            .I(\tok.n4775 ));
    InMux I__5272 (
            .O(N__23414),
            .I(bfn_11_10_0_));
    InMux I__5271 (
            .O(N__23411),
            .I(N__23407));
    InMux I__5270 (
            .O(N__23410),
            .I(N__23403));
    LocalMux I__5269 (
            .O(N__23407),
            .I(N__23399));
    InMux I__5268 (
            .O(N__23406),
            .I(N__23396));
    LocalMux I__5267 (
            .O(N__23403),
            .I(N__23393));
    InMux I__5266 (
            .O(N__23402),
            .I(N__23390));
    Span4Mux_v I__5265 (
            .O(N__23399),
            .I(N__23385));
    LocalMux I__5264 (
            .O(N__23396),
            .I(N__23385));
    Span4Mux_v I__5263 (
            .O(N__23393),
            .I(N__23378));
    LocalMux I__5262 (
            .O(N__23390),
            .I(N__23378));
    Span4Mux_h I__5261 (
            .O(N__23385),
            .I(N__23378));
    Span4Mux_h I__5260 (
            .O(N__23378),
            .I(N__23374));
    InMux I__5259 (
            .O(N__23377),
            .I(N__23371));
    Odrv4 I__5258 (
            .O(N__23374),
            .I(\tok.n11_adj_706 ));
    LocalMux I__5257 (
            .O(N__23371),
            .I(\tok.n11_adj_706 ));
    InMux I__5256 (
            .O(N__23366),
            .I(N__23362));
    InMux I__5255 (
            .O(N__23365),
            .I(N__23359));
    LocalMux I__5254 (
            .O(N__23362),
            .I(N__23356));
    LocalMux I__5253 (
            .O(N__23359),
            .I(uart_rx_data_2));
    Odrv12 I__5252 (
            .O(N__23356),
            .I(uart_rx_data_2));
    InMux I__5251 (
            .O(N__23351),
            .I(N__23348));
    LocalMux I__5250 (
            .O(N__23348),
            .I(N__23345));
    Span4Mux_v I__5249 (
            .O(N__23345),
            .I(N__23342));
    Odrv4 I__5248 (
            .O(N__23342),
            .I(\tok.n12_adj_832 ));
    CascadeMux I__5247 (
            .O(N__23339),
            .I(\tok.n6_adj_839_cascade_ ));
    InMux I__5246 (
            .O(N__23336),
            .I(N__23327));
    CascadeMux I__5245 (
            .O(N__23335),
            .I(N__23324));
    InMux I__5244 (
            .O(N__23334),
            .I(N__23321));
    InMux I__5243 (
            .O(N__23333),
            .I(N__23318));
    InMux I__5242 (
            .O(N__23332),
            .I(N__23315));
    InMux I__5241 (
            .O(N__23331),
            .I(N__23309));
    InMux I__5240 (
            .O(N__23330),
            .I(N__23309));
    LocalMux I__5239 (
            .O(N__23327),
            .I(N__23303));
    InMux I__5238 (
            .O(N__23324),
            .I(N__23300));
    LocalMux I__5237 (
            .O(N__23321),
            .I(N__23297));
    LocalMux I__5236 (
            .O(N__23318),
            .I(N__23292));
    LocalMux I__5235 (
            .O(N__23315),
            .I(N__23292));
    InMux I__5234 (
            .O(N__23314),
            .I(N__23289));
    LocalMux I__5233 (
            .O(N__23309),
            .I(N__23286));
    InMux I__5232 (
            .O(N__23308),
            .I(N__23279));
    InMux I__5231 (
            .O(N__23307),
            .I(N__23279));
    InMux I__5230 (
            .O(N__23306),
            .I(N__23279));
    Span4Mux_h I__5229 (
            .O(N__23303),
            .I(N__23275));
    LocalMux I__5228 (
            .O(N__23300),
            .I(N__23268));
    Span4Mux_v I__5227 (
            .O(N__23297),
            .I(N__23268));
    Span4Mux_h I__5226 (
            .O(N__23292),
            .I(N__23268));
    LocalMux I__5225 (
            .O(N__23289),
            .I(N__23263));
    Span4Mux_h I__5224 (
            .O(N__23286),
            .I(N__23263));
    LocalMux I__5223 (
            .O(N__23279),
            .I(N__23260));
    CascadeMux I__5222 (
            .O(N__23278),
            .I(N__23255));
    Span4Mux_h I__5221 (
            .O(N__23275),
            .I(N__23252));
    Span4Mux_h I__5220 (
            .O(N__23268),
            .I(N__23249));
    Span4Mux_h I__5219 (
            .O(N__23263),
            .I(N__23244));
    Span4Mux_h I__5218 (
            .O(N__23260),
            .I(N__23244));
    InMux I__5217 (
            .O(N__23259),
            .I(N__23239));
    InMux I__5216 (
            .O(N__23258),
            .I(N__23239));
    InMux I__5215 (
            .O(N__23255),
            .I(N__23236));
    Odrv4 I__5214 (
            .O(N__23252),
            .I(\tok.n11_adj_681 ));
    Odrv4 I__5213 (
            .O(N__23249),
            .I(\tok.n11_adj_681 ));
    Odrv4 I__5212 (
            .O(N__23244),
            .I(\tok.n11_adj_681 ));
    LocalMux I__5211 (
            .O(N__23239),
            .I(\tok.n11_adj_681 ));
    LocalMux I__5210 (
            .O(N__23236),
            .I(\tok.n11_adj_681 ));
    InMux I__5209 (
            .O(N__23225),
            .I(N__23222));
    LocalMux I__5208 (
            .O(N__23222),
            .I(N__23219));
    Span4Mux_h I__5207 (
            .O(N__23219),
            .I(N__23216));
    Odrv4 I__5206 (
            .O(N__23216),
            .I(\tok.n32 ));
    InMux I__5205 (
            .O(N__23213),
            .I(N__23209));
    InMux I__5204 (
            .O(N__23212),
            .I(N__23205));
    LocalMux I__5203 (
            .O(N__23209),
            .I(N__23201));
    InMux I__5202 (
            .O(N__23208),
            .I(N__23198));
    LocalMux I__5201 (
            .O(N__23205),
            .I(N__23195));
    InMux I__5200 (
            .O(N__23204),
            .I(N__23192));
    Span4Mux_v I__5199 (
            .O(N__23201),
            .I(N__23189));
    LocalMux I__5198 (
            .O(N__23198),
            .I(N__23186));
    Span4Mux_v I__5197 (
            .O(N__23195),
            .I(N__23183));
    LocalMux I__5196 (
            .O(N__23192),
            .I(N__23180));
    Span4Mux_v I__5195 (
            .O(N__23189),
            .I(N__23177));
    Span4Mux_v I__5194 (
            .O(N__23186),
            .I(N__23172));
    Span4Mux_s3_v I__5193 (
            .O(N__23183),
            .I(N__23172));
    Span4Mux_v I__5192 (
            .O(N__23180),
            .I(N__23169));
    Odrv4 I__5191 (
            .O(N__23177),
            .I(\tok.n15_adj_655 ));
    Odrv4 I__5190 (
            .O(N__23172),
            .I(\tok.n15_adj_655 ));
    Odrv4 I__5189 (
            .O(N__23169),
            .I(\tok.n15_adj_655 ));
    InMux I__5188 (
            .O(N__23162),
            .I(N__23159));
    LocalMux I__5187 (
            .O(N__23159),
            .I(N__23151));
    InMux I__5186 (
            .O(N__23158),
            .I(N__23147));
    InMux I__5185 (
            .O(N__23157),
            .I(N__23144));
    InMux I__5184 (
            .O(N__23156),
            .I(N__23141));
    InMux I__5183 (
            .O(N__23155),
            .I(N__23138));
    InMux I__5182 (
            .O(N__23154),
            .I(N__23135));
    Span4Mux_h I__5181 (
            .O(N__23151),
            .I(N__23132));
    InMux I__5180 (
            .O(N__23150),
            .I(N__23129));
    LocalMux I__5179 (
            .O(N__23147),
            .I(N__23126));
    LocalMux I__5178 (
            .O(N__23144),
            .I(N__23123));
    LocalMux I__5177 (
            .O(N__23141),
            .I(N__23120));
    LocalMux I__5176 (
            .O(N__23138),
            .I(N__23117));
    LocalMux I__5175 (
            .O(N__23135),
            .I(N__23113));
    Span4Mux_v I__5174 (
            .O(N__23132),
            .I(N__23102));
    LocalMux I__5173 (
            .O(N__23129),
            .I(N__23102));
    Span4Mux_h I__5172 (
            .O(N__23126),
            .I(N__23102));
    Span4Mux_h I__5171 (
            .O(N__23123),
            .I(N__23102));
    Span12Mux_s10_v I__5170 (
            .O(N__23120),
            .I(N__23099));
    Span4Mux_s3_h I__5169 (
            .O(N__23117),
            .I(N__23096));
    InMux I__5168 (
            .O(N__23116),
            .I(N__23093));
    Span4Mux_s3_v I__5167 (
            .O(N__23113),
            .I(N__23090));
    InMux I__5166 (
            .O(N__23112),
            .I(N__23085));
    InMux I__5165 (
            .O(N__23111),
            .I(N__23085));
    Span4Mux_v I__5164 (
            .O(N__23102),
            .I(N__23082));
    Odrv12 I__5163 (
            .O(N__23099),
            .I(\tok.A_13 ));
    Odrv4 I__5162 (
            .O(N__23096),
            .I(\tok.A_13 ));
    LocalMux I__5161 (
            .O(N__23093),
            .I(\tok.A_13 ));
    Odrv4 I__5160 (
            .O(N__23090),
            .I(\tok.A_13 ));
    LocalMux I__5159 (
            .O(N__23085),
            .I(\tok.A_13 ));
    Odrv4 I__5158 (
            .O(N__23082),
            .I(\tok.A_13 ));
    InMux I__5157 (
            .O(N__23069),
            .I(N__23066));
    LocalMux I__5156 (
            .O(N__23066),
            .I(N__23063));
    Span4Mux_v I__5155 (
            .O(N__23063),
            .I(N__23060));
    Span4Mux_h I__5154 (
            .O(N__23060),
            .I(N__23057));
    Odrv4 I__5153 (
            .O(N__23057),
            .I(\tok.n211 ));
    CascadeMux I__5152 (
            .O(N__23054),
            .I(N__23051));
    InMux I__5151 (
            .O(N__23051),
            .I(N__23048));
    LocalMux I__5150 (
            .O(N__23048),
            .I(N__23045));
    Span4Mux_h I__5149 (
            .O(N__23045),
            .I(N__23042));
    Odrv4 I__5148 (
            .O(N__23042),
            .I(\tok.n184 ));
    InMux I__5147 (
            .O(N__23039),
            .I(N__23036));
    LocalMux I__5146 (
            .O(N__23036),
            .I(N__23032));
    InMux I__5145 (
            .O(N__23035),
            .I(N__23029));
    Span4Mux_v I__5144 (
            .O(N__23032),
            .I(N__23024));
    LocalMux I__5143 (
            .O(N__23029),
            .I(N__23024));
    Span4Mux_h I__5142 (
            .O(N__23024),
            .I(N__23020));
    InMux I__5141 (
            .O(N__23023),
            .I(N__23017));
    Odrv4 I__5140 (
            .O(N__23020),
            .I(capture_5));
    LocalMux I__5139 (
            .O(N__23017),
            .I(capture_5));
    InMux I__5138 (
            .O(N__23012),
            .I(N__23009));
    LocalMux I__5137 (
            .O(N__23009),
            .I(N__23005));
    InMux I__5136 (
            .O(N__23008),
            .I(N__23002));
    Span4Mux_s2_h I__5135 (
            .O(N__23005),
            .I(N__22997));
    LocalMux I__5134 (
            .O(N__23002),
            .I(N__22997));
    Span4Mux_h I__5133 (
            .O(N__22997),
            .I(N__22994));
    Span4Mux_h I__5132 (
            .O(N__22994),
            .I(N__22990));
    InMux I__5131 (
            .O(N__22993),
            .I(N__22987));
    Odrv4 I__5130 (
            .O(N__22990),
            .I(capture_8));
    LocalMux I__5129 (
            .O(N__22987),
            .I(capture_8));
    InMux I__5128 (
            .O(N__22982),
            .I(N__22979));
    LocalMux I__5127 (
            .O(N__22979),
            .I(N__22967));
    InMux I__5126 (
            .O(N__22978),
            .I(N__22964));
    InMux I__5125 (
            .O(N__22977),
            .I(N__22957));
    InMux I__5124 (
            .O(N__22976),
            .I(N__22957));
    InMux I__5123 (
            .O(N__22975),
            .I(N__22957));
    InMux I__5122 (
            .O(N__22974),
            .I(N__22952));
    InMux I__5121 (
            .O(N__22973),
            .I(N__22952));
    InMux I__5120 (
            .O(N__22972),
            .I(N__22945));
    InMux I__5119 (
            .O(N__22971),
            .I(N__22945));
    InMux I__5118 (
            .O(N__22970),
            .I(N__22945));
    Span4Mux_v I__5117 (
            .O(N__22967),
            .I(N__22938));
    LocalMux I__5116 (
            .O(N__22964),
            .I(N__22938));
    LocalMux I__5115 (
            .O(N__22957),
            .I(N__22938));
    LocalMux I__5114 (
            .O(N__22952),
            .I(N__22935));
    LocalMux I__5113 (
            .O(N__22945),
            .I(N__22932));
    Span4Mux_v I__5112 (
            .O(N__22938),
            .I(N__22927));
    Span4Mux_h I__5111 (
            .O(N__22935),
            .I(N__22927));
    Span12Mux_s9_v I__5110 (
            .O(N__22932),
            .I(N__22924));
    Span4Mux_h I__5109 (
            .O(N__22927),
            .I(N__22921));
    Odrv12 I__5108 (
            .O(N__22924),
            .I(n4858));
    Odrv4 I__5107 (
            .O(N__22921),
            .I(n4858));
    InMux I__5106 (
            .O(N__22916),
            .I(N__22913));
    LocalMux I__5105 (
            .O(N__22913),
            .I(N__22910));
    Span4Mux_v I__5104 (
            .O(N__22910),
            .I(N__22907));
    Span4Mux_h I__5103 (
            .O(N__22907),
            .I(N__22902));
    InMux I__5102 (
            .O(N__22906),
            .I(N__22897));
    InMux I__5101 (
            .O(N__22905),
            .I(N__22897));
    Odrv4 I__5100 (
            .O(N__22902),
            .I(capture_7));
    LocalMux I__5099 (
            .O(N__22897),
            .I(capture_7));
    InMux I__5098 (
            .O(N__22892),
            .I(N__22889));
    LocalMux I__5097 (
            .O(N__22889),
            .I(\tok.n17_adj_711 ));
    InMux I__5096 (
            .O(N__22886),
            .I(N__22883));
    LocalMux I__5095 (
            .O(N__22883),
            .I(N__22876));
    InMux I__5094 (
            .O(N__22882),
            .I(N__22873));
    InMux I__5093 (
            .O(N__22881),
            .I(N__22868));
    CascadeMux I__5092 (
            .O(N__22880),
            .I(N__22865));
    CascadeMux I__5091 (
            .O(N__22879),
            .I(N__22862));
    Span4Mux_h I__5090 (
            .O(N__22876),
            .I(N__22857));
    LocalMux I__5089 (
            .O(N__22873),
            .I(N__22857));
    InMux I__5088 (
            .O(N__22872),
            .I(N__22854));
    CascadeMux I__5087 (
            .O(N__22871),
            .I(N__22850));
    LocalMux I__5086 (
            .O(N__22868),
            .I(N__22847));
    InMux I__5085 (
            .O(N__22865),
            .I(N__22844));
    InMux I__5084 (
            .O(N__22862),
            .I(N__22841));
    Span4Mux_v I__5083 (
            .O(N__22857),
            .I(N__22835));
    LocalMux I__5082 (
            .O(N__22854),
            .I(N__22835));
    InMux I__5081 (
            .O(N__22853),
            .I(N__22832));
    InMux I__5080 (
            .O(N__22850),
            .I(N__22829));
    Span4Mux_v I__5079 (
            .O(N__22847),
            .I(N__22824));
    LocalMux I__5078 (
            .O(N__22844),
            .I(N__22824));
    LocalMux I__5077 (
            .O(N__22841),
            .I(N__22821));
    InMux I__5076 (
            .O(N__22840),
            .I(N__22818));
    Span4Mux_h I__5075 (
            .O(N__22835),
            .I(N__22815));
    LocalMux I__5074 (
            .O(N__22832),
            .I(N__22812));
    LocalMux I__5073 (
            .O(N__22829),
            .I(N__22809));
    Span4Mux_h I__5072 (
            .O(N__22824),
            .I(N__22806));
    Span12Mux_v I__5071 (
            .O(N__22821),
            .I(N__22803));
    LocalMux I__5070 (
            .O(N__22818),
            .I(N__22798));
    Span4Mux_v I__5069 (
            .O(N__22815),
            .I(N__22798));
    Span12Mux_s6_h I__5068 (
            .O(N__22812),
            .I(N__22793));
    Span12Mux_s7_h I__5067 (
            .O(N__22809),
            .I(N__22793));
    Span4Mux_v I__5066 (
            .O(N__22806),
            .I(N__22790));
    Odrv12 I__5065 (
            .O(N__22803),
            .I(\tok.S_0 ));
    Odrv4 I__5064 (
            .O(N__22798),
            .I(\tok.S_0 ));
    Odrv12 I__5063 (
            .O(N__22793),
            .I(\tok.S_0 ));
    Odrv4 I__5062 (
            .O(N__22790),
            .I(\tok.S_0 ));
    InMux I__5061 (
            .O(N__22781),
            .I(N__22778));
    LocalMux I__5060 (
            .O(N__22778),
            .I(N__22775));
    Span4Mux_h I__5059 (
            .O(N__22775),
            .I(N__22772));
    Odrv4 I__5058 (
            .O(N__22772),
            .I(\tok.n11_adj_809 ));
    InMux I__5057 (
            .O(N__22769),
            .I(bfn_11_9_0_));
    InMux I__5056 (
            .O(N__22766),
            .I(N__22754));
    InMux I__5055 (
            .O(N__22765),
            .I(N__22751));
    InMux I__5054 (
            .O(N__22764),
            .I(N__22747));
    InMux I__5053 (
            .O(N__22763),
            .I(N__22742));
    InMux I__5052 (
            .O(N__22762),
            .I(N__22742));
    InMux I__5051 (
            .O(N__22761),
            .I(N__22739));
    InMux I__5050 (
            .O(N__22760),
            .I(N__22736));
    InMux I__5049 (
            .O(N__22759),
            .I(N__22733));
    InMux I__5048 (
            .O(N__22758),
            .I(N__22728));
    InMux I__5047 (
            .O(N__22757),
            .I(N__22725));
    LocalMux I__5046 (
            .O(N__22754),
            .I(N__22722));
    LocalMux I__5045 (
            .O(N__22751),
            .I(N__22719));
    InMux I__5044 (
            .O(N__22750),
            .I(N__22716));
    LocalMux I__5043 (
            .O(N__22747),
            .I(N__22711));
    LocalMux I__5042 (
            .O(N__22742),
            .I(N__22711));
    LocalMux I__5041 (
            .O(N__22739),
            .I(N__22702));
    LocalMux I__5040 (
            .O(N__22736),
            .I(N__22702));
    LocalMux I__5039 (
            .O(N__22733),
            .I(N__22702));
    InMux I__5038 (
            .O(N__22732),
            .I(N__22699));
    CascadeMux I__5037 (
            .O(N__22731),
            .I(N__22696));
    LocalMux I__5036 (
            .O(N__22728),
            .I(N__22693));
    LocalMux I__5035 (
            .O(N__22725),
            .I(N__22690));
    Span4Mux_h I__5034 (
            .O(N__22722),
            .I(N__22685));
    Span4Mux_h I__5033 (
            .O(N__22719),
            .I(N__22685));
    LocalMux I__5032 (
            .O(N__22716),
            .I(N__22682));
    Span12Mux_s9_v I__5031 (
            .O(N__22711),
            .I(N__22679));
    InMux I__5030 (
            .O(N__22710),
            .I(N__22674));
    InMux I__5029 (
            .O(N__22709),
            .I(N__22674));
    Span4Mux_v I__5028 (
            .O(N__22702),
            .I(N__22669));
    LocalMux I__5027 (
            .O(N__22699),
            .I(N__22669));
    InMux I__5026 (
            .O(N__22696),
            .I(N__22666));
    Span4Mux_v I__5025 (
            .O(N__22693),
            .I(N__22661));
    Span4Mux_v I__5024 (
            .O(N__22690),
            .I(N__22661));
    Odrv4 I__5023 (
            .O(N__22685),
            .I(\tok.A_low_2 ));
    Odrv4 I__5022 (
            .O(N__22682),
            .I(\tok.A_low_2 ));
    Odrv12 I__5021 (
            .O(N__22679),
            .I(\tok.A_low_2 ));
    LocalMux I__5020 (
            .O(N__22674),
            .I(\tok.A_low_2 ));
    Odrv4 I__5019 (
            .O(N__22669),
            .I(\tok.A_low_2 ));
    LocalMux I__5018 (
            .O(N__22666),
            .I(\tok.A_low_2 ));
    Odrv4 I__5017 (
            .O(N__22661),
            .I(\tok.A_low_2 ));
    InMux I__5016 (
            .O(N__22646),
            .I(N__22643));
    LocalMux I__5015 (
            .O(N__22643),
            .I(N__22640));
    Span4Mux_s3_h I__5014 (
            .O(N__22640),
            .I(N__22637));
    Odrv4 I__5013 (
            .O(N__22637),
            .I(\tok.n22_adj_698 ));
    InMux I__5012 (
            .O(N__22634),
            .I(N__22631));
    LocalMux I__5011 (
            .O(N__22631),
            .I(N__22628));
    Span4Mux_h I__5010 (
            .O(N__22628),
            .I(N__22625));
    Span4Mux_v I__5009 (
            .O(N__22625),
            .I(N__22622));
    Odrv4 I__5008 (
            .O(N__22622),
            .I(\tok.n24_adj_703 ));
    CascadeMux I__5007 (
            .O(N__22619),
            .I(\tok.n4_adj_699_cascade_ ));
    InMux I__5006 (
            .O(N__22616),
            .I(N__22613));
    LocalMux I__5005 (
            .O(N__22613),
            .I(N__22610));
    Span4Mux_h I__5004 (
            .O(N__22610),
            .I(N__22607));
    Odrv4 I__5003 (
            .O(N__22607),
            .I(\tok.n9_adj_705 ));
    InMux I__5002 (
            .O(N__22604),
            .I(N__22601));
    LocalMux I__5001 (
            .O(N__22601),
            .I(N__22597));
    InMux I__5000 (
            .O(N__22600),
            .I(N__22594));
    Span4Mux_s3_h I__4999 (
            .O(N__22597),
            .I(N__22591));
    LocalMux I__4998 (
            .O(N__22594),
            .I(uart_rx_data_1));
    Odrv4 I__4997 (
            .O(N__22591),
            .I(uart_rx_data_1));
    InMux I__4996 (
            .O(N__22586),
            .I(N__22583));
    LocalMux I__4995 (
            .O(N__22583),
            .I(N__22580));
    Span12Mux_s4_h I__4994 (
            .O(N__22580),
            .I(N__22577));
    Odrv12 I__4993 (
            .O(N__22577),
            .I(\tok.n14_adj_662 ));
    InMux I__4992 (
            .O(N__22574),
            .I(N__22571));
    LocalMux I__4991 (
            .O(N__22571),
            .I(\tok.n6_adj_834 ));
    InMux I__4990 (
            .O(N__22568),
            .I(N__22565));
    LocalMux I__4989 (
            .O(N__22565),
            .I(N__22562));
    Span4Mux_v I__4988 (
            .O(N__22562),
            .I(N__22559));
    Span4Mux_h I__4987 (
            .O(N__22559),
            .I(N__22556));
    Odrv4 I__4986 (
            .O(N__22556),
            .I(\tok.n23_adj_718 ));
    CascadeMux I__4985 (
            .O(N__22553),
            .I(\tok.n5_adj_835_cascade_ ));
    InMux I__4984 (
            .O(N__22550),
            .I(N__22536));
    InMux I__4983 (
            .O(N__22549),
            .I(N__22533));
    InMux I__4982 (
            .O(N__22548),
            .I(N__22530));
    CascadeMux I__4981 (
            .O(N__22547),
            .I(N__22524));
    CascadeMux I__4980 (
            .O(N__22546),
            .I(N__22520));
    CascadeMux I__4979 (
            .O(N__22545),
            .I(N__22517));
    InMux I__4978 (
            .O(N__22544),
            .I(N__22512));
    InMux I__4977 (
            .O(N__22543),
            .I(N__22512));
    CascadeMux I__4976 (
            .O(N__22542),
            .I(N__22498));
    CascadeMux I__4975 (
            .O(N__22541),
            .I(N__22493));
    CascadeMux I__4974 (
            .O(N__22540),
            .I(N__22489));
    InMux I__4973 (
            .O(N__22539),
            .I(N__22486));
    LocalMux I__4972 (
            .O(N__22536),
            .I(N__22482));
    LocalMux I__4971 (
            .O(N__22533),
            .I(N__22474));
    LocalMux I__4970 (
            .O(N__22530),
            .I(N__22474));
    InMux I__4969 (
            .O(N__22529),
            .I(N__22469));
    InMux I__4968 (
            .O(N__22528),
            .I(N__22469));
    InMux I__4967 (
            .O(N__22527),
            .I(N__22466));
    InMux I__4966 (
            .O(N__22524),
            .I(N__22457));
    InMux I__4965 (
            .O(N__22523),
            .I(N__22457));
    InMux I__4964 (
            .O(N__22520),
            .I(N__22457));
    InMux I__4963 (
            .O(N__22517),
            .I(N__22457));
    LocalMux I__4962 (
            .O(N__22512),
            .I(N__22454));
    InMux I__4961 (
            .O(N__22511),
            .I(N__22451));
    CascadeMux I__4960 (
            .O(N__22510),
            .I(N__22447));
    InMux I__4959 (
            .O(N__22509),
            .I(N__22432));
    InMux I__4958 (
            .O(N__22508),
            .I(N__22432));
    InMux I__4957 (
            .O(N__22507),
            .I(N__22432));
    InMux I__4956 (
            .O(N__22506),
            .I(N__22432));
    InMux I__4955 (
            .O(N__22505),
            .I(N__22432));
    InMux I__4954 (
            .O(N__22504),
            .I(N__22432));
    InMux I__4953 (
            .O(N__22503),
            .I(N__22432));
    InMux I__4952 (
            .O(N__22502),
            .I(N__22415));
    InMux I__4951 (
            .O(N__22501),
            .I(N__22415));
    InMux I__4950 (
            .O(N__22498),
            .I(N__22415));
    InMux I__4949 (
            .O(N__22497),
            .I(N__22415));
    InMux I__4948 (
            .O(N__22496),
            .I(N__22415));
    InMux I__4947 (
            .O(N__22493),
            .I(N__22415));
    InMux I__4946 (
            .O(N__22492),
            .I(N__22415));
    InMux I__4945 (
            .O(N__22489),
            .I(N__22415));
    LocalMux I__4944 (
            .O(N__22486),
            .I(N__22412));
    InMux I__4943 (
            .O(N__22485),
            .I(N__22408));
    Span4Mux_v I__4942 (
            .O(N__22482),
            .I(N__22405));
    InMux I__4941 (
            .O(N__22481),
            .I(N__22398));
    InMux I__4940 (
            .O(N__22480),
            .I(N__22398));
    InMux I__4939 (
            .O(N__22479),
            .I(N__22398));
    Span4Mux_v I__4938 (
            .O(N__22474),
            .I(N__22389));
    LocalMux I__4937 (
            .O(N__22469),
            .I(N__22389));
    LocalMux I__4936 (
            .O(N__22466),
            .I(N__22389));
    LocalMux I__4935 (
            .O(N__22457),
            .I(N__22389));
    Span4Mux_h I__4934 (
            .O(N__22454),
            .I(N__22384));
    LocalMux I__4933 (
            .O(N__22451),
            .I(N__22384));
    InMux I__4932 (
            .O(N__22450),
            .I(N__22379));
    InMux I__4931 (
            .O(N__22447),
            .I(N__22379));
    LocalMux I__4930 (
            .O(N__22432),
            .I(N__22374));
    LocalMux I__4929 (
            .O(N__22415),
            .I(N__22374));
    Span4Mux_v I__4928 (
            .O(N__22412),
            .I(N__22371));
    InMux I__4927 (
            .O(N__22411),
            .I(N__22368));
    LocalMux I__4926 (
            .O(N__22408),
            .I(N__22361));
    Span4Mux_v I__4925 (
            .O(N__22405),
            .I(N__22361));
    LocalMux I__4924 (
            .O(N__22398),
            .I(N__22361));
    Span4Mux_h I__4923 (
            .O(N__22389),
            .I(N__22358));
    Span4Mux_h I__4922 (
            .O(N__22384),
            .I(N__22353));
    LocalMux I__4921 (
            .O(N__22379),
            .I(N__22353));
    Odrv4 I__4920 (
            .O(N__22374),
            .I(\tok.n14_adj_644 ));
    Odrv4 I__4919 (
            .O(N__22371),
            .I(\tok.n14_adj_644 ));
    LocalMux I__4918 (
            .O(N__22368),
            .I(\tok.n14_adj_644 ));
    Odrv4 I__4917 (
            .O(N__22361),
            .I(\tok.n14_adj_644 ));
    Odrv4 I__4916 (
            .O(N__22358),
            .I(\tok.n14_adj_644 ));
    Odrv4 I__4915 (
            .O(N__22353),
            .I(\tok.n14_adj_644 ));
    InMux I__4914 (
            .O(N__22340),
            .I(N__22337));
    LocalMux I__4913 (
            .O(N__22337),
            .I(N__22334));
    Span4Mux_h I__4912 (
            .O(N__22334),
            .I(N__22331));
    Odrv4 I__4911 (
            .O(N__22331),
            .I(\tok.n10_adj_836 ));
    InMux I__4910 (
            .O(N__22328),
            .I(N__22323));
    InMux I__4909 (
            .O(N__22327),
            .I(N__22317));
    InMux I__4908 (
            .O(N__22326),
            .I(N__22314));
    LocalMux I__4907 (
            .O(N__22323),
            .I(N__22307));
    InMux I__4906 (
            .O(N__22322),
            .I(N__22304));
    CascadeMux I__4905 (
            .O(N__22321),
            .I(N__22300));
    CascadeMux I__4904 (
            .O(N__22320),
            .I(N__22296));
    LocalMux I__4903 (
            .O(N__22317),
            .I(N__22293));
    LocalMux I__4902 (
            .O(N__22314),
            .I(N__22290));
    CascadeMux I__4901 (
            .O(N__22313),
            .I(N__22287));
    InMux I__4900 (
            .O(N__22312),
            .I(N__22282));
    InMux I__4899 (
            .O(N__22311),
            .I(N__22282));
    InMux I__4898 (
            .O(N__22310),
            .I(N__22279));
    Span4Mux_v I__4897 (
            .O(N__22307),
            .I(N__22276));
    LocalMux I__4896 (
            .O(N__22304),
            .I(N__22273));
    InMux I__4895 (
            .O(N__22303),
            .I(N__22270));
    InMux I__4894 (
            .O(N__22300),
            .I(N__22265));
    InMux I__4893 (
            .O(N__22299),
            .I(N__22262));
    InMux I__4892 (
            .O(N__22296),
            .I(N__22259));
    Span4Mux_v I__4891 (
            .O(N__22293),
            .I(N__22253));
    Span4Mux_v I__4890 (
            .O(N__22290),
            .I(N__22253));
    InMux I__4889 (
            .O(N__22287),
            .I(N__22250));
    LocalMux I__4888 (
            .O(N__22282),
            .I(N__22247));
    LocalMux I__4887 (
            .O(N__22279),
            .I(N__22244));
    Span4Mux_h I__4886 (
            .O(N__22276),
            .I(N__22237));
    Span4Mux_h I__4885 (
            .O(N__22273),
            .I(N__22237));
    LocalMux I__4884 (
            .O(N__22270),
            .I(N__22237));
    InMux I__4883 (
            .O(N__22269),
            .I(N__22234));
    InMux I__4882 (
            .O(N__22268),
            .I(N__22231));
    LocalMux I__4881 (
            .O(N__22265),
            .I(N__22228));
    LocalMux I__4880 (
            .O(N__22262),
            .I(N__22225));
    LocalMux I__4879 (
            .O(N__22259),
            .I(N__22222));
    InMux I__4878 (
            .O(N__22258),
            .I(N__22219));
    Span4Mux_h I__4877 (
            .O(N__22253),
            .I(N__22210));
    LocalMux I__4876 (
            .O(N__22250),
            .I(N__22210));
    Span4Mux_v I__4875 (
            .O(N__22247),
            .I(N__22210));
    Span4Mux_v I__4874 (
            .O(N__22244),
            .I(N__22210));
    Sp12to4 I__4873 (
            .O(N__22237),
            .I(N__22203));
    LocalMux I__4872 (
            .O(N__22234),
            .I(N__22203));
    LocalMux I__4871 (
            .O(N__22231),
            .I(N__22203));
    Span4Mux_v I__4870 (
            .O(N__22228),
            .I(N__22196));
    Span4Mux_v I__4869 (
            .O(N__22225),
            .I(N__22196));
    Span4Mux_v I__4868 (
            .O(N__22222),
            .I(N__22196));
    LocalMux I__4867 (
            .O(N__22219),
            .I(A_low_7));
    Odrv4 I__4866 (
            .O(N__22210),
            .I(A_low_7));
    Odrv12 I__4865 (
            .O(N__22203),
            .I(A_low_7));
    Odrv4 I__4864 (
            .O(N__22196),
            .I(A_low_7));
    CascadeMux I__4863 (
            .O(N__22187),
            .I(N__22183));
    InMux I__4862 (
            .O(N__22186),
            .I(N__22179));
    InMux I__4861 (
            .O(N__22183),
            .I(N__22174));
    InMux I__4860 (
            .O(N__22182),
            .I(N__22174));
    LocalMux I__4859 (
            .O(N__22179),
            .I(N__22171));
    LocalMux I__4858 (
            .O(N__22174),
            .I(N__22167));
    Span4Mux_h I__4857 (
            .O(N__22171),
            .I(N__22164));
    InMux I__4856 (
            .O(N__22170),
            .I(N__22161));
    Span4Mux_v I__4855 (
            .O(N__22167),
            .I(N__22158));
    Odrv4 I__4854 (
            .O(N__22164),
            .I(\tok.n6_adj_650 ));
    LocalMux I__4853 (
            .O(N__22161),
            .I(\tok.n6_adj_650 ));
    Odrv4 I__4852 (
            .O(N__22158),
            .I(\tok.n6_adj_650 ));
    InMux I__4851 (
            .O(N__22151),
            .I(N__22147));
    InMux I__4850 (
            .O(N__22150),
            .I(N__22136));
    LocalMux I__4849 (
            .O(N__22147),
            .I(N__22131));
    InMux I__4848 (
            .O(N__22146),
            .I(N__22126));
    InMux I__4847 (
            .O(N__22145),
            .I(N__22126));
    InMux I__4846 (
            .O(N__22144),
            .I(N__22123));
    InMux I__4845 (
            .O(N__22143),
            .I(N__22116));
    InMux I__4844 (
            .O(N__22142),
            .I(N__22116));
    InMux I__4843 (
            .O(N__22141),
            .I(N__22116));
    InMux I__4842 (
            .O(N__22140),
            .I(N__22111));
    InMux I__4841 (
            .O(N__22139),
            .I(N__22111));
    LocalMux I__4840 (
            .O(N__22136),
            .I(N__22104));
    InMux I__4839 (
            .O(N__22135),
            .I(N__22099));
    InMux I__4838 (
            .O(N__22134),
            .I(N__22099));
    Span4Mux_v I__4837 (
            .O(N__22131),
            .I(N__22094));
    LocalMux I__4836 (
            .O(N__22126),
            .I(N__22094));
    LocalMux I__4835 (
            .O(N__22123),
            .I(N__22089));
    LocalMux I__4834 (
            .O(N__22116),
            .I(N__22089));
    LocalMux I__4833 (
            .O(N__22111),
            .I(N__22086));
    InMux I__4832 (
            .O(N__22110),
            .I(N__22083));
    InMux I__4831 (
            .O(N__22109),
            .I(N__22078));
    InMux I__4830 (
            .O(N__22108),
            .I(N__22078));
    CascadeMux I__4829 (
            .O(N__22107),
            .I(N__22074));
    Span4Mux_s3_v I__4828 (
            .O(N__22104),
            .I(N__22069));
    LocalMux I__4827 (
            .O(N__22099),
            .I(N__22069));
    Span4Mux_h I__4826 (
            .O(N__22094),
            .I(N__22064));
    Span4Mux_v I__4825 (
            .O(N__22089),
            .I(N__22064));
    Span4Mux_h I__4824 (
            .O(N__22086),
            .I(N__22060));
    LocalMux I__4823 (
            .O(N__22083),
            .I(N__22057));
    LocalMux I__4822 (
            .O(N__22078),
            .I(N__22054));
    InMux I__4821 (
            .O(N__22077),
            .I(N__22049));
    InMux I__4820 (
            .O(N__22074),
            .I(N__22049));
    Span4Mux_v I__4819 (
            .O(N__22069),
            .I(N__22044));
    Span4Mux_h I__4818 (
            .O(N__22064),
            .I(N__22044));
    InMux I__4817 (
            .O(N__22063),
            .I(N__22041));
    Span4Mux_v I__4816 (
            .O(N__22060),
            .I(N__22038));
    Span4Mux_s3_v I__4815 (
            .O(N__22057),
            .I(N__22033));
    Span4Mux_v I__4814 (
            .O(N__22054),
            .I(N__22033));
    LocalMux I__4813 (
            .O(N__22049),
            .I(N__22030));
    Odrv4 I__4812 (
            .O(N__22044),
            .I(\tok.T_7 ));
    LocalMux I__4811 (
            .O(N__22041),
            .I(\tok.T_7 ));
    Odrv4 I__4810 (
            .O(N__22038),
            .I(\tok.T_7 ));
    Odrv4 I__4809 (
            .O(N__22033),
            .I(\tok.T_7 ));
    Odrv12 I__4808 (
            .O(N__22030),
            .I(\tok.T_7 ));
    InMux I__4807 (
            .O(N__22019),
            .I(N__22013));
    InMux I__4806 (
            .O(N__22018),
            .I(N__22013));
    LocalMux I__4805 (
            .O(N__22013),
            .I(\tok.A_stk.tail_8 ));
    CascadeMux I__4804 (
            .O(N__22010),
            .I(N__22006));
    CascadeMux I__4803 (
            .O(N__22009),
            .I(N__22003));
    InMux I__4802 (
            .O(N__22006),
            .I(N__21998));
    InMux I__4801 (
            .O(N__22003),
            .I(N__21998));
    LocalMux I__4800 (
            .O(N__21998),
            .I(\tok.A_stk.tail_24 ));
    InMux I__4799 (
            .O(N__21995),
            .I(N__21992));
    LocalMux I__4798 (
            .O(N__21992),
            .I(N__21989));
    Span4Mux_v I__4797 (
            .O(N__21989),
            .I(N__21985));
    InMux I__4796 (
            .O(N__21988),
            .I(N__21982));
    Odrv4 I__4795 (
            .O(N__21985),
            .I(\tok.A_stk.tail_56 ));
    LocalMux I__4794 (
            .O(N__21982),
            .I(\tok.A_stk.tail_56 ));
    InMux I__4793 (
            .O(N__21977),
            .I(N__21974));
    LocalMux I__4792 (
            .O(N__21974),
            .I(N__21970));
    InMux I__4791 (
            .O(N__21973),
            .I(N__21967));
    Span4Mux_h I__4790 (
            .O(N__21970),
            .I(N__21964));
    LocalMux I__4789 (
            .O(N__21967),
            .I(\tok.A_stk.tail_40 ));
    Odrv4 I__4788 (
            .O(N__21964),
            .I(\tok.A_stk.tail_40 ));
    InMux I__4787 (
            .O(N__21959),
            .I(N__21956));
    LocalMux I__4786 (
            .O(N__21956),
            .I(N__21953));
    Odrv4 I__4785 (
            .O(N__21953),
            .I(\tok.n22 ));
    CascadeMux I__4784 (
            .O(N__21950),
            .I(N__21947));
    InMux I__4783 (
            .O(N__21947),
            .I(N__21944));
    LocalMux I__4782 (
            .O(N__21944),
            .I(N__21941));
    Span4Mux_s3_h I__4781 (
            .O(N__21941),
            .I(N__21938));
    Span4Mux_v I__4780 (
            .O(N__21938),
            .I(N__21935));
    Odrv4 I__4779 (
            .O(N__21935),
            .I(\tok.n24 ));
    InMux I__4778 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__4777 (
            .O(N__21929),
            .I(N__21926));
    Span4Mux_s3_h I__4776 (
            .O(N__21926),
            .I(N__21923));
    Span4Mux_h I__4775 (
            .O(N__21923),
            .I(N__21920));
    Odrv4 I__4774 (
            .O(N__21920),
            .I(\tok.n21 ));
    CascadeMux I__4773 (
            .O(N__21917),
            .I(\tok.n30_cascade_ ));
    InMux I__4772 (
            .O(N__21914),
            .I(N__21911));
    LocalMux I__4771 (
            .O(N__21911),
            .I(N__21907));
    InMux I__4770 (
            .O(N__21910),
            .I(N__21904));
    Span12Mux_s8_v I__4769 (
            .O(N__21907),
            .I(N__21899));
    LocalMux I__4768 (
            .O(N__21904),
            .I(N__21899));
    Odrv12 I__4767 (
            .O(N__21899),
            .I(\tok.n15_adj_671 ));
    InMux I__4766 (
            .O(N__21896),
            .I(N__21890));
    InMux I__4765 (
            .O(N__21895),
            .I(N__21887));
    CascadeMux I__4764 (
            .O(N__21894),
            .I(N__21883));
    InMux I__4763 (
            .O(N__21893),
            .I(N__21880));
    LocalMux I__4762 (
            .O(N__21890),
            .I(N__21877));
    LocalMux I__4761 (
            .O(N__21887),
            .I(N__21872));
    InMux I__4760 (
            .O(N__21886),
            .I(N__21869));
    InMux I__4759 (
            .O(N__21883),
            .I(N__21861));
    LocalMux I__4758 (
            .O(N__21880),
            .I(N__21856));
    Span4Mux_h I__4757 (
            .O(N__21877),
            .I(N__21856));
    InMux I__4756 (
            .O(N__21876),
            .I(N__21851));
    InMux I__4755 (
            .O(N__21875),
            .I(N__21851));
    Span4Mux_v I__4754 (
            .O(N__21872),
            .I(N__21846));
    LocalMux I__4753 (
            .O(N__21869),
            .I(N__21846));
    InMux I__4752 (
            .O(N__21868),
            .I(N__21841));
    InMux I__4751 (
            .O(N__21867),
            .I(N__21841));
    InMux I__4750 (
            .O(N__21866),
            .I(N__21836));
    InMux I__4749 (
            .O(N__21865),
            .I(N__21836));
    InMux I__4748 (
            .O(N__21864),
            .I(N__21831));
    LocalMux I__4747 (
            .O(N__21861),
            .I(N__21827));
    Span4Mux_h I__4746 (
            .O(N__21856),
            .I(N__21818));
    LocalMux I__4745 (
            .O(N__21851),
            .I(N__21818));
    Span4Mux_h I__4744 (
            .O(N__21846),
            .I(N__21818));
    LocalMux I__4743 (
            .O(N__21841),
            .I(N__21818));
    LocalMux I__4742 (
            .O(N__21836),
            .I(N__21815));
    InMux I__4741 (
            .O(N__21835),
            .I(N__21812));
    InMux I__4740 (
            .O(N__21834),
            .I(N__21809));
    LocalMux I__4739 (
            .O(N__21831),
            .I(N__21806));
    InMux I__4738 (
            .O(N__21830),
            .I(N__21803));
    Span4Mux_h I__4737 (
            .O(N__21827),
            .I(N__21798));
    Span4Mux_v I__4736 (
            .O(N__21818),
            .I(N__21798));
    Span4Mux_v I__4735 (
            .O(N__21815),
            .I(N__21795));
    LocalMux I__4734 (
            .O(N__21812),
            .I(\tok.A_low_6 ));
    LocalMux I__4733 (
            .O(N__21809),
            .I(\tok.A_low_6 ));
    Odrv12 I__4732 (
            .O(N__21806),
            .I(\tok.A_low_6 ));
    LocalMux I__4731 (
            .O(N__21803),
            .I(\tok.A_low_6 ));
    Odrv4 I__4730 (
            .O(N__21798),
            .I(\tok.A_low_6 ));
    Odrv4 I__4729 (
            .O(N__21795),
            .I(\tok.A_low_6 ));
    InMux I__4728 (
            .O(N__21782),
            .I(N__21779));
    LocalMux I__4727 (
            .O(N__21779),
            .I(N__21776));
    Span4Mux_s3_h I__4726 (
            .O(N__21776),
            .I(N__21773));
    Span4Mux_v I__4725 (
            .O(N__21773),
            .I(N__21770));
    Odrv4 I__4724 (
            .O(N__21770),
            .I(\tok.n18 ));
    CascadeMux I__4723 (
            .O(N__21767),
            .I(\tok.n17_adj_661_cascade_ ));
    InMux I__4722 (
            .O(N__21764),
            .I(N__21761));
    LocalMux I__4721 (
            .O(N__21761),
            .I(\tok.n19 ));
    InMux I__4720 (
            .O(N__21758),
            .I(N__21755));
    LocalMux I__4719 (
            .O(N__21755),
            .I(\tok.n29 ));
    InMux I__4718 (
            .O(N__21752),
            .I(N__21749));
    LocalMux I__4717 (
            .O(N__21749),
            .I(N__21746));
    Span4Mux_h I__4716 (
            .O(N__21746),
            .I(N__21742));
    InMux I__4715 (
            .O(N__21745),
            .I(N__21739));
    Odrv4 I__4714 (
            .O(N__21742),
            .I(\tok.A_stk.tail_7 ));
    LocalMux I__4713 (
            .O(N__21739),
            .I(\tok.A_stk.tail_7 ));
    InMux I__4712 (
            .O(N__21734),
            .I(N__21728));
    InMux I__4711 (
            .O(N__21733),
            .I(N__21728));
    LocalMux I__4710 (
            .O(N__21728),
            .I(\tok.A_stk.tail_2 ));
    InMux I__4709 (
            .O(N__21725),
            .I(N__21719));
    InMux I__4708 (
            .O(N__21724),
            .I(N__21719));
    LocalMux I__4707 (
            .O(N__21719),
            .I(\tok.A_stk.tail_18 ));
    InMux I__4706 (
            .O(N__21716),
            .I(N__21710));
    InMux I__4705 (
            .O(N__21715),
            .I(N__21710));
    LocalMux I__4704 (
            .O(N__21710),
            .I(\tok.A_stk.tail_34 ));
    InMux I__4703 (
            .O(N__21707),
            .I(N__21704));
    LocalMux I__4702 (
            .O(N__21704),
            .I(N__21700));
    InMux I__4701 (
            .O(N__21703),
            .I(N__21697));
    Odrv4 I__4700 (
            .O(N__21700),
            .I(\tok.A_stk.tail_66 ));
    LocalMux I__4699 (
            .O(N__21697),
            .I(\tok.A_stk.tail_66 ));
    InMux I__4698 (
            .O(N__21692),
            .I(N__21688));
    InMux I__4697 (
            .O(N__21691),
            .I(N__21685));
    LocalMux I__4696 (
            .O(N__21688),
            .I(N__21682));
    LocalMux I__4695 (
            .O(N__21685),
            .I(\tok.A_stk.tail_50 ));
    Odrv4 I__4694 (
            .O(N__21682),
            .I(\tok.A_stk.tail_50 ));
    InMux I__4693 (
            .O(N__21677),
            .I(N__21674));
    LocalMux I__4692 (
            .O(N__21674),
            .I(N__21670));
    InMux I__4691 (
            .O(N__21673),
            .I(N__21667));
    Odrv4 I__4690 (
            .O(N__21670),
            .I(\tok.A_stk.tail_44 ));
    LocalMux I__4689 (
            .O(N__21667),
            .I(\tok.A_stk.tail_44 ));
    InMux I__4688 (
            .O(N__21662),
            .I(N__21658));
    InMux I__4687 (
            .O(N__21661),
            .I(N__21655));
    LocalMux I__4686 (
            .O(N__21658),
            .I(N__21652));
    LocalMux I__4685 (
            .O(N__21655),
            .I(\tok.A_stk.tail_28 ));
    Odrv4 I__4684 (
            .O(N__21652),
            .I(\tok.A_stk.tail_28 ));
    CascadeMux I__4683 (
            .O(N__21647),
            .I(N__21644));
    InMux I__4682 (
            .O(N__21644),
            .I(N__21638));
    InMux I__4681 (
            .O(N__21643),
            .I(N__21638));
    LocalMux I__4680 (
            .O(N__21638),
            .I(\tok.A_stk.tail_12 ));
    InMux I__4679 (
            .O(N__21635),
            .I(N__21626));
    InMux I__4678 (
            .O(N__21634),
            .I(N__21626));
    InMux I__4677 (
            .O(N__21633),
            .I(N__21623));
    InMux I__4676 (
            .O(N__21632),
            .I(N__21620));
    CascadeMux I__4675 (
            .O(N__21631),
            .I(N__21616));
    LocalMux I__4674 (
            .O(N__21626),
            .I(N__21613));
    LocalMux I__4673 (
            .O(N__21623),
            .I(N__21608));
    LocalMux I__4672 (
            .O(N__21620),
            .I(N__21605));
    InMux I__4671 (
            .O(N__21619),
            .I(N__21600));
    InMux I__4670 (
            .O(N__21616),
            .I(N__21600));
    Span4Mux_s3_h I__4669 (
            .O(N__21613),
            .I(N__21596));
    InMux I__4668 (
            .O(N__21612),
            .I(N__21592));
    InMux I__4667 (
            .O(N__21611),
            .I(N__21589));
    Span4Mux_h I__4666 (
            .O(N__21608),
            .I(N__21582));
    Span4Mux_v I__4665 (
            .O(N__21605),
            .I(N__21582));
    LocalMux I__4664 (
            .O(N__21600),
            .I(N__21582));
    InMux I__4663 (
            .O(N__21599),
            .I(N__21579));
    Span4Mux_v I__4662 (
            .O(N__21596),
            .I(N__21576));
    InMux I__4661 (
            .O(N__21595),
            .I(N__21573));
    LocalMux I__4660 (
            .O(N__21592),
            .I(N__21566));
    LocalMux I__4659 (
            .O(N__21589),
            .I(N__21566));
    Span4Mux_h I__4658 (
            .O(N__21582),
            .I(N__21566));
    LocalMux I__4657 (
            .O(N__21579),
            .I(\tok.A_12 ));
    Odrv4 I__4656 (
            .O(N__21576),
            .I(\tok.A_12 ));
    LocalMux I__4655 (
            .O(N__21573),
            .I(\tok.A_12 ));
    Odrv4 I__4654 (
            .O(N__21566),
            .I(\tok.A_12 ));
    InMux I__4653 (
            .O(N__21557),
            .I(N__21554));
    LocalMux I__4652 (
            .O(N__21554),
            .I(N__21550));
    InMux I__4651 (
            .O(N__21553),
            .I(N__21547));
    Odrv4 I__4650 (
            .O(N__21550),
            .I(tail_107));
    LocalMux I__4649 (
            .O(N__21547),
            .I(tail_107));
    InMux I__4648 (
            .O(N__21542),
            .I(N__21538));
    InMux I__4647 (
            .O(N__21541),
            .I(N__21535));
    LocalMux I__4646 (
            .O(N__21538),
            .I(\tok.A_stk.tail_91 ));
    LocalMux I__4645 (
            .O(N__21535),
            .I(\tok.A_stk.tail_91 ));
    CascadeMux I__4644 (
            .O(N__21530),
            .I(N__21526));
    InMux I__4643 (
            .O(N__21529),
            .I(N__21523));
    InMux I__4642 (
            .O(N__21526),
            .I(N__21520));
    LocalMux I__4641 (
            .O(N__21523),
            .I(N__21517));
    LocalMux I__4640 (
            .O(N__21520),
            .I(N__21514));
    Odrv4 I__4639 (
            .O(N__21517),
            .I(tail_124));
    Odrv4 I__4638 (
            .O(N__21514),
            .I(tail_124));
    InMux I__4637 (
            .O(N__21509),
            .I(N__21506));
    LocalMux I__4636 (
            .O(N__21506),
            .I(N__21502));
    InMux I__4635 (
            .O(N__21505),
            .I(N__21499));
    Odrv4 I__4634 (
            .O(N__21502),
            .I(tail_108));
    LocalMux I__4633 (
            .O(N__21499),
            .I(tail_108));
    InMux I__4632 (
            .O(N__21494),
            .I(N__21488));
    InMux I__4631 (
            .O(N__21493),
            .I(N__21488));
    LocalMux I__4630 (
            .O(N__21488),
            .I(\tok.A_stk.tail_92 ));
    InMux I__4629 (
            .O(N__21485),
            .I(N__21479));
    InMux I__4628 (
            .O(N__21484),
            .I(N__21479));
    LocalMux I__4627 (
            .O(N__21479),
            .I(\tok.A_stk.tail_76 ));
    InMux I__4626 (
            .O(N__21476),
            .I(N__21470));
    InMux I__4625 (
            .O(N__21475),
            .I(N__21470));
    LocalMux I__4624 (
            .O(N__21470),
            .I(\tok.A_stk.tail_60 ));
    InMux I__4623 (
            .O(N__21467),
            .I(N__21464));
    LocalMux I__4622 (
            .O(N__21464),
            .I(N__21461));
    Span4Mux_s2_v I__4621 (
            .O(N__21461),
            .I(N__21457));
    CascadeMux I__4620 (
            .O(N__21460),
            .I(N__21454));
    Span4Mux_s1_h I__4619 (
            .O(N__21457),
            .I(N__21451));
    InMux I__4618 (
            .O(N__21454),
            .I(N__21448));
    Odrv4 I__4617 (
            .O(N__21451),
            .I(tail_125));
    LocalMux I__4616 (
            .O(N__21448),
            .I(tail_125));
    InMux I__4615 (
            .O(N__21443),
            .I(N__21440));
    LocalMux I__4614 (
            .O(N__21440),
            .I(N__21437));
    Span4Mux_h I__4613 (
            .O(N__21437),
            .I(N__21433));
    InMux I__4612 (
            .O(N__21436),
            .I(N__21430));
    Odrv4 I__4611 (
            .O(N__21433),
            .I(tail_109));
    LocalMux I__4610 (
            .O(N__21430),
            .I(tail_109));
    InMux I__4609 (
            .O(N__21425),
            .I(N__21421));
    InMux I__4608 (
            .O(N__21424),
            .I(N__21418));
    LocalMux I__4607 (
            .O(N__21421),
            .I(\tok.A_stk.tail_93 ));
    LocalMux I__4606 (
            .O(N__21418),
            .I(\tok.A_stk.tail_93 ));
    InMux I__4605 (
            .O(N__21413),
            .I(N__21407));
    InMux I__4604 (
            .O(N__21412),
            .I(N__21407));
    LocalMux I__4603 (
            .O(N__21407),
            .I(\tok.A_stk.tail_77 ));
    InMux I__4602 (
            .O(N__21404),
            .I(N__21398));
    InMux I__4601 (
            .O(N__21403),
            .I(N__21398));
    LocalMux I__4600 (
            .O(N__21398),
            .I(\tok.A_stk.tail_61 ));
    InMux I__4599 (
            .O(N__21395),
            .I(N__21389));
    InMux I__4598 (
            .O(N__21394),
            .I(N__21389));
    LocalMux I__4597 (
            .O(N__21389),
            .I(\tok.A_stk.tail_45 ));
    InMux I__4596 (
            .O(N__21386),
            .I(N__21380));
    InMux I__4595 (
            .O(N__21385),
            .I(N__21380));
    LocalMux I__4594 (
            .O(N__21380),
            .I(\tok.A_stk.tail_29 ));
    CascadeMux I__4593 (
            .O(N__21377),
            .I(N__21374));
    InMux I__4592 (
            .O(N__21374),
            .I(N__21368));
    InMux I__4591 (
            .O(N__21373),
            .I(N__21368));
    LocalMux I__4590 (
            .O(N__21368),
            .I(\tok.A_stk.tail_13 ));
    InMux I__4589 (
            .O(N__21365),
            .I(N__21362));
    LocalMux I__4588 (
            .O(N__21362),
            .I(N__21358));
    InMux I__4587 (
            .O(N__21361),
            .I(N__21355));
    Odrv12 I__4586 (
            .O(N__21358),
            .I(tail_123));
    LocalMux I__4585 (
            .O(N__21355),
            .I(tail_123));
    CascadeMux I__4584 (
            .O(N__21350),
            .I(\tok.n13_adj_746_cascade_ ));
    InMux I__4583 (
            .O(N__21347),
            .I(N__21344));
    LocalMux I__4582 (
            .O(N__21344),
            .I(\tok.n12_adj_745 ));
    InMux I__4581 (
            .O(N__21341),
            .I(N__21338));
    LocalMux I__4580 (
            .O(N__21338),
            .I(N__21335));
    Span4Mux_v I__4579 (
            .O(N__21335),
            .I(N__21332));
    Odrv4 I__4578 (
            .O(N__21332),
            .I(\tok.n5525 ));
    InMux I__4577 (
            .O(N__21329),
            .I(N__21326));
    LocalMux I__4576 (
            .O(N__21326),
            .I(\tok.n16_adj_749 ));
    CascadeMux I__4575 (
            .O(N__21323),
            .I(\tok.n20_adj_753_cascade_ ));
    InMux I__4574 (
            .O(N__21320),
            .I(N__21317));
    LocalMux I__4573 (
            .O(N__21317),
            .I(\tok.n5522 ));
    CascadeMux I__4572 (
            .O(N__21314),
            .I(N__21308));
    CascadeMux I__4571 (
            .O(N__21313),
            .I(N__21305));
    CascadeMux I__4570 (
            .O(N__21312),
            .I(N__21301));
    InMux I__4569 (
            .O(N__21311),
            .I(N__21298));
    InMux I__4568 (
            .O(N__21308),
            .I(N__21295));
    InMux I__4567 (
            .O(N__21305),
            .I(N__21292));
    InMux I__4566 (
            .O(N__21304),
            .I(N__21289));
    InMux I__4565 (
            .O(N__21301),
            .I(N__21286));
    LocalMux I__4564 (
            .O(N__21298),
            .I(N__21275));
    LocalMux I__4563 (
            .O(N__21295),
            .I(N__21275));
    LocalMux I__4562 (
            .O(N__21292),
            .I(N__21275));
    LocalMux I__4561 (
            .O(N__21289),
            .I(N__21275));
    LocalMux I__4560 (
            .O(N__21286),
            .I(N__21275));
    Span4Mux_v I__4559 (
            .O(N__21275),
            .I(N__21272));
    Odrv4 I__4558 (
            .O(N__21272),
            .I(\tok.n8 ));
    InMux I__4557 (
            .O(N__21269),
            .I(N__21266));
    LocalMux I__4556 (
            .O(N__21266),
            .I(\tok.n14_adj_744 ));
    InMux I__4555 (
            .O(N__21263),
            .I(N__21260));
    LocalMux I__4554 (
            .O(N__21260),
            .I(\tok.n9_adj_748 ));
    InMux I__4553 (
            .O(N__21257),
            .I(N__21254));
    LocalMux I__4552 (
            .O(N__21254),
            .I(\tok.n2_adj_743 ));
    CascadeMux I__4551 (
            .O(N__21251),
            .I(\tok.n204_cascade_ ));
    InMux I__4550 (
            .O(N__21248),
            .I(N__21245));
    LocalMux I__4549 (
            .O(N__21245),
            .I(N__21242));
    Odrv12 I__4548 (
            .O(N__21242),
            .I(\tok.n16_adj_741 ));
    InMux I__4547 (
            .O(N__21239),
            .I(N__21236));
    LocalMux I__4546 (
            .O(N__21236),
            .I(N__21233));
    Odrv4 I__4545 (
            .O(N__21233),
            .I(\tok.n2 ));
    InMux I__4544 (
            .O(N__21230),
            .I(N__21227));
    LocalMux I__4543 (
            .O(N__21227),
            .I(\tok.n14_adj_722 ));
    InMux I__4542 (
            .O(N__21224),
            .I(N__21221));
    LocalMux I__4541 (
            .O(N__21221),
            .I(N__21218));
    Odrv12 I__4540 (
            .O(N__21218),
            .I(\tok.n20_adj_740 ));
    CascadeMux I__4539 (
            .O(N__21215),
            .I(\tok.n5527_cascade_ ));
    InMux I__4538 (
            .O(N__21212),
            .I(N__21209));
    LocalMux I__4537 (
            .O(N__21209),
            .I(\tok.n5513 ));
    InMux I__4536 (
            .O(N__21206),
            .I(N__21203));
    LocalMux I__4535 (
            .O(N__21203),
            .I(N__21200));
    Odrv4 I__4534 (
            .O(N__21200),
            .I(\tok.n5539 ));
    CascadeMux I__4533 (
            .O(N__21197),
            .I(N__21194));
    InMux I__4532 (
            .O(N__21194),
            .I(N__21191));
    LocalMux I__4531 (
            .O(N__21191),
            .I(\tok.n5348 ));
    InMux I__4530 (
            .O(N__21188),
            .I(N__21185));
    LocalMux I__4529 (
            .O(N__21185),
            .I(N__21180));
    InMux I__4528 (
            .O(N__21184),
            .I(N__21177));
    InMux I__4527 (
            .O(N__21183),
            .I(N__21174));
    Span4Mux_v I__4526 (
            .O(N__21180),
            .I(N__21171));
    LocalMux I__4525 (
            .O(N__21177),
            .I(N__21168));
    LocalMux I__4524 (
            .O(N__21174),
            .I(N__21165));
    Odrv4 I__4523 (
            .O(N__21171),
            .I(capture_2));
    Odrv4 I__4522 (
            .O(N__21168),
            .I(capture_2));
    Odrv4 I__4521 (
            .O(N__21165),
            .I(capture_2));
    InMux I__4520 (
            .O(N__21158),
            .I(N__21155));
    LocalMux I__4519 (
            .O(N__21155),
            .I(\tok.n9 ));
    CascadeMux I__4518 (
            .O(N__21152),
            .I(\tok.n5342_cascade_ ));
    InMux I__4517 (
            .O(N__21149),
            .I(N__21146));
    LocalMux I__4516 (
            .O(N__21146),
            .I(\tok.n10_adj_686 ));
    InMux I__4515 (
            .O(N__21143),
            .I(N__21137));
    InMux I__4514 (
            .O(N__21142),
            .I(N__21132));
    InMux I__4513 (
            .O(N__21141),
            .I(N__21128));
    InMux I__4512 (
            .O(N__21140),
            .I(N__21125));
    LocalMux I__4511 (
            .O(N__21137),
            .I(N__21122));
    InMux I__4510 (
            .O(N__21136),
            .I(N__21119));
    InMux I__4509 (
            .O(N__21135),
            .I(N__21116));
    LocalMux I__4508 (
            .O(N__21132),
            .I(N__21112));
    InMux I__4507 (
            .O(N__21131),
            .I(N__21104));
    LocalMux I__4506 (
            .O(N__21128),
            .I(N__21100));
    LocalMux I__4505 (
            .O(N__21125),
            .I(N__21097));
    Span4Mux_v I__4504 (
            .O(N__21122),
            .I(N__21094));
    LocalMux I__4503 (
            .O(N__21119),
            .I(N__21091));
    LocalMux I__4502 (
            .O(N__21116),
            .I(N__21088));
    InMux I__4501 (
            .O(N__21115),
            .I(N__21085));
    Span4Mux_h I__4500 (
            .O(N__21112),
            .I(N__21081));
    InMux I__4499 (
            .O(N__21111),
            .I(N__21076));
    InMux I__4498 (
            .O(N__21110),
            .I(N__21076));
    InMux I__4497 (
            .O(N__21109),
            .I(N__21073));
    CascadeMux I__4496 (
            .O(N__21108),
            .I(N__21070));
    InMux I__4495 (
            .O(N__21107),
            .I(N__21067));
    LocalMux I__4494 (
            .O(N__21104),
            .I(N__21064));
    InMux I__4493 (
            .O(N__21103),
            .I(N__21061));
    Span4Mux_v I__4492 (
            .O(N__21100),
            .I(N__21056));
    Span4Mux_v I__4491 (
            .O(N__21097),
            .I(N__21056));
    Span4Mux_v I__4490 (
            .O(N__21094),
            .I(N__21047));
    Span4Mux_h I__4489 (
            .O(N__21091),
            .I(N__21047));
    Span4Mux_h I__4488 (
            .O(N__21088),
            .I(N__21047));
    LocalMux I__4487 (
            .O(N__21085),
            .I(N__21047));
    InMux I__4486 (
            .O(N__21084),
            .I(N__21044));
    Span4Mux_v I__4485 (
            .O(N__21081),
            .I(N__21037));
    LocalMux I__4484 (
            .O(N__21076),
            .I(N__21037));
    LocalMux I__4483 (
            .O(N__21073),
            .I(N__21037));
    InMux I__4482 (
            .O(N__21070),
            .I(N__21034));
    LocalMux I__4481 (
            .O(N__21067),
            .I(N__21031));
    Span4Mux_h I__4480 (
            .O(N__21064),
            .I(N__21026));
    LocalMux I__4479 (
            .O(N__21061),
            .I(N__21026));
    Odrv4 I__4478 (
            .O(N__21056),
            .I(\tok.A_low_1 ));
    Odrv4 I__4477 (
            .O(N__21047),
            .I(\tok.A_low_1 ));
    LocalMux I__4476 (
            .O(N__21044),
            .I(\tok.A_low_1 ));
    Odrv4 I__4475 (
            .O(N__21037),
            .I(\tok.A_low_1 ));
    LocalMux I__4474 (
            .O(N__21034),
            .I(\tok.A_low_1 ));
    Odrv4 I__4473 (
            .O(N__21031),
            .I(\tok.A_low_1 ));
    Odrv4 I__4472 (
            .O(N__21026),
            .I(\tok.A_low_1 ));
    InMux I__4471 (
            .O(N__21011),
            .I(N__21008));
    LocalMux I__4470 (
            .O(N__21008),
            .I(\tok.n5336 ));
    InMux I__4469 (
            .O(N__21005),
            .I(N__21002));
    LocalMux I__4468 (
            .O(N__21002),
            .I(N__20999));
    Span4Mux_v I__4467 (
            .O(N__20999),
            .I(N__20996));
    Span4Mux_h I__4466 (
            .O(N__20996),
            .I(N__20993));
    Sp12to4 I__4465 (
            .O(N__20993),
            .I(N__20990));
    Odrv12 I__4464 (
            .O(N__20990),
            .I(\tok.table_rd_11 ));
    InMux I__4463 (
            .O(N__20987),
            .I(N__20984));
    LocalMux I__4462 (
            .O(N__20984),
            .I(N__20981));
    Span4Mux_v I__4461 (
            .O(N__20981),
            .I(N__20978));
    Odrv4 I__4460 (
            .O(N__20978),
            .I(\tok.n5_adj_726 ));
    CascadeMux I__4459 (
            .O(N__20975),
            .I(\tok.n13_adj_724_cascade_ ));
    InMux I__4458 (
            .O(N__20972),
            .I(N__20969));
    LocalMux I__4457 (
            .O(N__20969),
            .I(\tok.n12_adj_723 ));
    InMux I__4456 (
            .O(N__20966),
            .I(N__20963));
    LocalMux I__4455 (
            .O(N__20963),
            .I(N__20960));
    Odrv12 I__4454 (
            .O(N__20960),
            .I(\tok.n5534 ));
    InMux I__4453 (
            .O(N__20957),
            .I(N__20954));
    LocalMux I__4452 (
            .O(N__20954),
            .I(\tok.n16 ));
    CascadeMux I__4451 (
            .O(N__20951),
            .I(\tok.n20_adj_729_cascade_ ));
    InMux I__4450 (
            .O(N__20948),
            .I(N__20945));
    LocalMux I__4449 (
            .O(N__20945),
            .I(\tok.n9_adj_725 ));
    CascadeMux I__4448 (
            .O(N__20942),
            .I(N__20939));
    InMux I__4447 (
            .O(N__20939),
            .I(N__20936));
    LocalMux I__4446 (
            .O(N__20936),
            .I(N__20933));
    Odrv4 I__4445 (
            .O(N__20933),
            .I(\tok.n5531 ));
    CascadeMux I__4444 (
            .O(N__20930),
            .I(\tok.n1_cascade_ ));
    InMux I__4443 (
            .O(N__20927),
            .I(N__20924));
    LocalMux I__4442 (
            .O(N__20924),
            .I(N__20921));
    Span4Mux_h I__4441 (
            .O(N__20921),
            .I(N__20918));
    Odrv4 I__4440 (
            .O(N__20918),
            .I(\tok.n17_adj_656 ));
    InMux I__4439 (
            .O(N__20915),
            .I(N__20912));
    LocalMux I__4438 (
            .O(N__20912),
            .I(\tok.n12 ));
    InMux I__4437 (
            .O(N__20909),
            .I(N__20903));
    InMux I__4436 (
            .O(N__20908),
            .I(N__20903));
    LocalMux I__4435 (
            .O(N__20903),
            .I(uart_rx_data_7));
    CascadeMux I__4434 (
            .O(N__20900),
            .I(N__20897));
    InMux I__4433 (
            .O(N__20897),
            .I(N__20894));
    LocalMux I__4432 (
            .O(N__20894),
            .I(\tok.n177 ));
    InMux I__4431 (
            .O(N__20891),
            .I(N__20888));
    LocalMux I__4430 (
            .O(N__20888),
            .I(N__20885));
    Odrv4 I__4429 (
            .O(N__20885),
            .I(\tok.n17_adj_812 ));
    CascadeMux I__4428 (
            .O(N__20882),
            .I(N__20879));
    InMux I__4427 (
            .O(N__20879),
            .I(N__20876));
    LocalMux I__4426 (
            .O(N__20876),
            .I(\tok.n9_adj_838 ));
    InMux I__4425 (
            .O(N__20873),
            .I(N__20870));
    LocalMux I__4424 (
            .O(N__20870),
            .I(N__20867));
    Span4Mux_v I__4423 (
            .O(N__20867),
            .I(N__20864));
    Odrv4 I__4422 (
            .O(N__20864),
            .I(\tok.n23_adj_682 ));
    InMux I__4421 (
            .O(N__20861),
            .I(N__20858));
    LocalMux I__4420 (
            .O(N__20858),
            .I(\tok.n25 ));
    CascadeMux I__4419 (
            .O(N__20855),
            .I(\tok.n4_cascade_ ));
    InMux I__4418 (
            .O(N__20852),
            .I(N__20849));
    LocalMux I__4417 (
            .O(N__20849),
            .I(\tok.n5350 ));
    InMux I__4416 (
            .O(N__20846),
            .I(\tok.n4807 ));
    InMux I__4415 (
            .O(N__20843),
            .I(N__20833));
    InMux I__4414 (
            .O(N__20842),
            .I(N__20833));
    InMux I__4413 (
            .O(N__20841),
            .I(N__20830));
    InMux I__4412 (
            .O(N__20840),
            .I(N__20827));
    InMux I__4411 (
            .O(N__20839),
            .I(N__20822));
    InMux I__4410 (
            .O(N__20838),
            .I(N__20822));
    LocalMux I__4409 (
            .O(N__20833),
            .I(N__20813));
    LocalMux I__4408 (
            .O(N__20830),
            .I(N__20813));
    LocalMux I__4407 (
            .O(N__20827),
            .I(N__20813));
    LocalMux I__4406 (
            .O(N__20822),
            .I(N__20813));
    Span4Mux_v I__4405 (
            .O(N__20813),
            .I(N__20810));
    Span4Mux_h I__4404 (
            .O(N__20810),
            .I(N__20807));
    Odrv4 I__4403 (
            .O(N__20807),
            .I(\tok.n20_adj_663 ));
    InMux I__4402 (
            .O(N__20804),
            .I(\tok.n4808 ));
    InMux I__4401 (
            .O(N__20801),
            .I(\tok.n4809 ));
    InMux I__4400 (
            .O(N__20798),
            .I(N__20795));
    LocalMux I__4399 (
            .O(N__20795),
            .I(N__20792));
    Odrv4 I__4398 (
            .O(N__20792),
            .I(\tok.n10_adj_738 ));
    InMux I__4397 (
            .O(N__20789),
            .I(\tok.n4810 ));
    InMux I__4396 (
            .O(N__20786),
            .I(\tok.n4811 ));
    InMux I__4395 (
            .O(N__20783),
            .I(N__20780));
    LocalMux I__4394 (
            .O(N__20780),
            .I(N__20777));
    Span4Mux_v I__4393 (
            .O(N__20777),
            .I(N__20774));
    Odrv4 I__4392 (
            .O(N__20774),
            .I(\tok.n10_adj_768 ));
    InMux I__4391 (
            .O(N__20771),
            .I(\tok.n4812 ));
    InMux I__4390 (
            .O(N__20768),
            .I(N__20757));
    InMux I__4389 (
            .O(N__20767),
            .I(N__20757));
    InMux I__4388 (
            .O(N__20766),
            .I(N__20752));
    InMux I__4387 (
            .O(N__20765),
            .I(N__20752));
    SRMux I__4386 (
            .O(N__20764),
            .I(N__20745));
    InMux I__4385 (
            .O(N__20763),
            .I(N__20740));
    InMux I__4384 (
            .O(N__20762),
            .I(N__20740));
    LocalMux I__4383 (
            .O(N__20757),
            .I(N__20737));
    LocalMux I__4382 (
            .O(N__20752),
            .I(N__20734));
    InMux I__4381 (
            .O(N__20751),
            .I(N__20725));
    InMux I__4380 (
            .O(N__20750),
            .I(N__20725));
    InMux I__4379 (
            .O(N__20749),
            .I(N__20725));
    InMux I__4378 (
            .O(N__20748),
            .I(N__20725));
    LocalMux I__4377 (
            .O(N__20745),
            .I(N__20722));
    LocalMux I__4376 (
            .O(N__20740),
            .I(N__20713));
    Span4Mux_v I__4375 (
            .O(N__20737),
            .I(N__20713));
    Span4Mux_v I__4374 (
            .O(N__20734),
            .I(N__20713));
    LocalMux I__4373 (
            .O(N__20725),
            .I(N__20713));
    Span4Mux_v I__4372 (
            .O(N__20722),
            .I(N__20710));
    Span4Mux_h I__4371 (
            .O(N__20713),
            .I(N__20707));
    Odrv4 I__4370 (
            .O(N__20710),
            .I(\tok.write_flag ));
    Odrv4 I__4369 (
            .O(N__20707),
            .I(\tok.write_flag ));
    InMux I__4368 (
            .O(N__20702),
            .I(\tok.n4813 ));
    InMux I__4367 (
            .O(N__20699),
            .I(N__20696));
    LocalMux I__4366 (
            .O(N__20696),
            .I(N__20693));
    Span4Mux_h I__4365 (
            .O(N__20693),
            .I(N__20690));
    Span4Mux_v I__4364 (
            .O(N__20690),
            .I(N__20687));
    Odrv4 I__4363 (
            .O(N__20687),
            .I(\tok.n5516 ));
    InMux I__4362 (
            .O(N__20684),
            .I(N__20681));
    LocalMux I__4361 (
            .O(N__20681),
            .I(N__20678));
    Span4Mux_v I__4360 (
            .O(N__20678),
            .I(N__20675));
    Sp12to4 I__4359 (
            .O(N__20675),
            .I(N__20672));
    Odrv12 I__4358 (
            .O(N__20672),
            .I(\tok.n18_adj_739 ));
    CascadeMux I__4357 (
            .O(N__20669),
            .I(\tok.n12_adj_737_cascade_ ));
    InMux I__4356 (
            .O(N__20666),
            .I(bfn_9_6_0_));
    InMux I__4355 (
            .O(N__20663),
            .I(\tok.n4799 ));
    InMux I__4354 (
            .O(N__20660),
            .I(\tok.n4800 ));
    InMux I__4353 (
            .O(N__20657),
            .I(N__20654));
    LocalMux I__4352 (
            .O(N__20654),
            .I(N__20651));
    Span4Mux_h I__4351 (
            .O(N__20651),
            .I(N__20648));
    Odrv4 I__4350 (
            .O(N__20648),
            .I(\tok.n22_adj_829 ));
    InMux I__4349 (
            .O(N__20645),
            .I(\tok.n4801 ));
    InMux I__4348 (
            .O(N__20642),
            .I(N__20639));
    LocalMux I__4347 (
            .O(N__20639),
            .I(N__20636));
    Span4Mux_h I__4346 (
            .O(N__20636),
            .I(N__20633));
    Odrv4 I__4345 (
            .O(N__20633),
            .I(\tok.n10_adj_827 ));
    InMux I__4344 (
            .O(N__20630),
            .I(\tok.n4802 ));
    InMux I__4343 (
            .O(N__20627),
            .I(\tok.n4803 ));
    InMux I__4342 (
            .O(N__20624),
            .I(N__20621));
    LocalMux I__4341 (
            .O(N__20621),
            .I(\tok.n10_adj_820 ));
    InMux I__4340 (
            .O(N__20618),
            .I(\tok.n4804 ));
    InMux I__4339 (
            .O(N__20615),
            .I(N__20612));
    LocalMux I__4338 (
            .O(N__20612),
            .I(\tok.n10_adj_653 ));
    InMux I__4337 (
            .O(N__20609),
            .I(\tok.n4805 ));
    InMux I__4336 (
            .O(N__20606),
            .I(bfn_9_7_0_));
    InMux I__4335 (
            .O(N__20603),
            .I(N__20599));
    InMux I__4334 (
            .O(N__20602),
            .I(N__20596));
    LocalMux I__4333 (
            .O(N__20599),
            .I(N__20593));
    LocalMux I__4332 (
            .O(N__20596),
            .I(\tok.A_stk.tail_86 ));
    Odrv4 I__4331 (
            .O(N__20593),
            .I(\tok.A_stk.tail_86 ));
    InMux I__4330 (
            .O(N__20588),
            .I(N__20584));
    InMux I__4329 (
            .O(N__20587),
            .I(N__20581));
    LocalMux I__4328 (
            .O(N__20584),
            .I(\tok.A_stk.tail_55 ));
    LocalMux I__4327 (
            .O(N__20581),
            .I(\tok.A_stk.tail_55 ));
    InMux I__4326 (
            .O(N__20576),
            .I(N__20572));
    InMux I__4325 (
            .O(N__20575),
            .I(N__20569));
    LocalMux I__4324 (
            .O(N__20572),
            .I(\tok.A_stk.tail_39 ));
    LocalMux I__4323 (
            .O(N__20569),
            .I(\tok.A_stk.tail_39 ));
    InMux I__4322 (
            .O(N__20564),
            .I(N__20561));
    LocalMux I__4321 (
            .O(N__20561),
            .I(N__20557));
    InMux I__4320 (
            .O(N__20560),
            .I(N__20554));
    Odrv4 I__4319 (
            .O(N__20557),
            .I(\tok.A_stk.tail_83 ));
    LocalMux I__4318 (
            .O(N__20554),
            .I(\tok.A_stk.tail_83 ));
    InMux I__4317 (
            .O(N__20549),
            .I(N__20545));
    InMux I__4316 (
            .O(N__20548),
            .I(N__20542));
    LocalMux I__4315 (
            .O(N__20545),
            .I(\tok.A_stk.tail_4 ));
    LocalMux I__4314 (
            .O(N__20542),
            .I(\tok.A_stk.tail_4 ));
    InMux I__4313 (
            .O(N__20537),
            .I(N__20531));
    InMux I__4312 (
            .O(N__20536),
            .I(N__20531));
    LocalMux I__4311 (
            .O(N__20531),
            .I(\tok.A_stk.tail_6 ));
    CascadeMux I__4310 (
            .O(N__20528),
            .I(N__20525));
    InMux I__4309 (
            .O(N__20525),
            .I(N__20521));
    InMux I__4308 (
            .O(N__20524),
            .I(N__20518));
    LocalMux I__4307 (
            .O(N__20521),
            .I(\tok.A_stk.tail_54 ));
    LocalMux I__4306 (
            .O(N__20518),
            .I(\tok.A_stk.tail_54 ));
    InMux I__4305 (
            .O(N__20513),
            .I(N__20507));
    InMux I__4304 (
            .O(N__20512),
            .I(N__20507));
    LocalMux I__4303 (
            .O(N__20507),
            .I(\tok.A_stk.tail_22 ));
    InMux I__4302 (
            .O(N__20504),
            .I(N__20501));
    LocalMux I__4301 (
            .O(N__20501),
            .I(N__20497));
    InMux I__4300 (
            .O(N__20500),
            .I(N__20494));
    Odrv4 I__4299 (
            .O(N__20497),
            .I(\tok.A_stk.tail_38 ));
    LocalMux I__4298 (
            .O(N__20494),
            .I(\tok.A_stk.tail_38 ));
    InMux I__4297 (
            .O(N__20489),
            .I(N__20485));
    InMux I__4296 (
            .O(N__20488),
            .I(N__20482));
    LocalMux I__4295 (
            .O(N__20485),
            .I(\tok.A_stk.tail_23 ));
    LocalMux I__4294 (
            .O(N__20482),
            .I(\tok.A_stk.tail_23 ));
    InMux I__4293 (
            .O(N__20477),
            .I(N__20474));
    LocalMux I__4292 (
            .O(N__20474),
            .I(N__20471));
    Odrv4 I__4291 (
            .O(N__20471),
            .I(\tok.n3_adj_692 ));
    InMux I__4290 (
            .O(N__20468),
            .I(N__20465));
    LocalMux I__4289 (
            .O(N__20465),
            .I(N__20461));
    InMux I__4288 (
            .O(N__20464),
            .I(N__20458));
    Odrv4 I__4287 (
            .O(N__20461),
            .I(tail_100));
    LocalMux I__4286 (
            .O(N__20458),
            .I(tail_100));
    InMux I__4285 (
            .O(N__20453),
            .I(N__20450));
    LocalMux I__4284 (
            .O(N__20450),
            .I(N__20446));
    InMux I__4283 (
            .O(N__20449),
            .I(N__20443));
    Odrv4 I__4282 (
            .O(N__20446),
            .I(tail_116));
    LocalMux I__4281 (
            .O(N__20443),
            .I(tail_116));
    InMux I__4280 (
            .O(N__20438),
            .I(N__20434));
    CascadeMux I__4279 (
            .O(N__20437),
            .I(N__20431));
    LocalMux I__4278 (
            .O(N__20434),
            .I(N__20428));
    InMux I__4277 (
            .O(N__20431),
            .I(N__20425));
    Odrv4 I__4276 (
            .O(N__20428),
            .I(tail_114));
    LocalMux I__4275 (
            .O(N__20425),
            .I(tail_114));
    InMux I__4274 (
            .O(N__20420),
            .I(N__20416));
    InMux I__4273 (
            .O(N__20419),
            .I(N__20413));
    LocalMux I__4272 (
            .O(N__20416),
            .I(N__20410));
    LocalMux I__4271 (
            .O(N__20413),
            .I(tail_98));
    Odrv4 I__4270 (
            .O(N__20410),
            .I(tail_98));
    CascadeMux I__4269 (
            .O(N__20405),
            .I(N__20402));
    InMux I__4268 (
            .O(N__20402),
            .I(N__20396));
    InMux I__4267 (
            .O(N__20401),
            .I(N__20396));
    LocalMux I__4266 (
            .O(N__20396),
            .I(\tok.A_stk.tail_82 ));
    InMux I__4265 (
            .O(N__20393),
            .I(N__20389));
    InMux I__4264 (
            .O(N__20392),
            .I(N__20386));
    LocalMux I__4263 (
            .O(N__20389),
            .I(\tok.A_stk.tail_72 ));
    LocalMux I__4262 (
            .O(N__20386),
            .I(\tok.A_stk.tail_72 ));
    InMux I__4261 (
            .O(N__20381),
            .I(N__20377));
    InMux I__4260 (
            .O(N__20380),
            .I(N__20374));
    LocalMux I__4259 (
            .O(N__20377),
            .I(N__20371));
    LocalMux I__4258 (
            .O(N__20374),
            .I(tail_102));
    Odrv12 I__4257 (
            .O(N__20371),
            .I(tail_102));
    InMux I__4256 (
            .O(N__20366),
            .I(N__20360));
    InMux I__4255 (
            .O(N__20365),
            .I(N__20360));
    LocalMux I__4254 (
            .O(N__20360),
            .I(\tok.A_stk.tail_70 ));
    InMux I__4253 (
            .O(N__20357),
            .I(N__20354));
    LocalMux I__4252 (
            .O(N__20354),
            .I(\tok.n209 ));
    InMux I__4251 (
            .O(N__20351),
            .I(N__20348));
    LocalMux I__4250 (
            .O(N__20348),
            .I(N__20345));
    Odrv12 I__4249 (
            .O(N__20345),
            .I(\tok.n14_adj_658 ));
    InMux I__4248 (
            .O(N__20342),
            .I(N__20339));
    LocalMux I__4247 (
            .O(N__20339),
            .I(N__20336));
    Odrv4 I__4246 (
            .O(N__20336),
            .I(\tok.n2_adj_775 ));
    InMux I__4245 (
            .O(N__20333),
            .I(N__20329));
    InMux I__4244 (
            .O(N__20332),
            .I(N__20326));
    LocalMux I__4243 (
            .O(N__20329),
            .I(tail_118));
    LocalMux I__4242 (
            .O(N__20326),
            .I(tail_118));
    InMux I__4241 (
            .O(N__20321),
            .I(N__20318));
    LocalMux I__4240 (
            .O(N__20318),
            .I(\tok.n14_adj_764 ));
    InMux I__4239 (
            .O(N__20315),
            .I(N__20304));
    InMux I__4238 (
            .O(N__20314),
            .I(N__20304));
    InMux I__4237 (
            .O(N__20313),
            .I(N__20304));
    InMux I__4236 (
            .O(N__20312),
            .I(N__20299));
    InMux I__4235 (
            .O(N__20311),
            .I(N__20299));
    LocalMux I__4234 (
            .O(N__20304),
            .I(N__20286));
    LocalMux I__4233 (
            .O(N__20299),
            .I(N__20286));
    InMux I__4232 (
            .O(N__20298),
            .I(N__20281));
    InMux I__4231 (
            .O(N__20297),
            .I(N__20281));
    InMux I__4230 (
            .O(N__20296),
            .I(N__20273));
    InMux I__4229 (
            .O(N__20295),
            .I(N__20254));
    InMux I__4228 (
            .O(N__20294),
            .I(N__20254));
    InMux I__4227 (
            .O(N__20293),
            .I(N__20254));
    InMux I__4226 (
            .O(N__20292),
            .I(N__20254));
    InMux I__4225 (
            .O(N__20291),
            .I(N__20254));
    Span4Mux_v I__4224 (
            .O(N__20286),
            .I(N__20249));
    LocalMux I__4223 (
            .O(N__20281),
            .I(N__20249));
    CascadeMux I__4222 (
            .O(N__20280),
            .I(N__20246));
    CascadeMux I__4221 (
            .O(N__20279),
            .I(N__20241));
    InMux I__4220 (
            .O(N__20278),
            .I(N__20233));
    InMux I__4219 (
            .O(N__20277),
            .I(N__20233));
    InMux I__4218 (
            .O(N__20276),
            .I(N__20224));
    LocalMux I__4217 (
            .O(N__20273),
            .I(N__20221));
    InMux I__4216 (
            .O(N__20272),
            .I(N__20218));
    InMux I__4215 (
            .O(N__20271),
            .I(N__20213));
    InMux I__4214 (
            .O(N__20270),
            .I(N__20213));
    InMux I__4213 (
            .O(N__20269),
            .I(N__20208));
    InMux I__4212 (
            .O(N__20268),
            .I(N__20208));
    InMux I__4211 (
            .O(N__20267),
            .I(N__20201));
    InMux I__4210 (
            .O(N__20266),
            .I(N__20201));
    InMux I__4209 (
            .O(N__20265),
            .I(N__20201));
    LocalMux I__4208 (
            .O(N__20254),
            .I(N__20196));
    Span4Mux_h I__4207 (
            .O(N__20249),
            .I(N__20196));
    InMux I__4206 (
            .O(N__20246),
            .I(N__20183));
    InMux I__4205 (
            .O(N__20245),
            .I(N__20183));
    InMux I__4204 (
            .O(N__20244),
            .I(N__20183));
    InMux I__4203 (
            .O(N__20241),
            .I(N__20183));
    InMux I__4202 (
            .O(N__20240),
            .I(N__20183));
    InMux I__4201 (
            .O(N__20239),
            .I(N__20178));
    InMux I__4200 (
            .O(N__20238),
            .I(N__20178));
    LocalMux I__4199 (
            .O(N__20233),
            .I(N__20175));
    InMux I__4198 (
            .O(N__20232),
            .I(N__20172));
    InMux I__4197 (
            .O(N__20231),
            .I(N__20169));
    InMux I__4196 (
            .O(N__20230),
            .I(N__20159));
    InMux I__4195 (
            .O(N__20229),
            .I(N__20156));
    InMux I__4194 (
            .O(N__20228),
            .I(N__20151));
    InMux I__4193 (
            .O(N__20227),
            .I(N__20151));
    LocalMux I__4192 (
            .O(N__20224),
            .I(N__20146));
    Span4Mux_v I__4191 (
            .O(N__20221),
            .I(N__20146));
    LocalMux I__4190 (
            .O(N__20218),
            .I(N__20140));
    LocalMux I__4189 (
            .O(N__20213),
            .I(N__20140));
    LocalMux I__4188 (
            .O(N__20208),
            .I(N__20133));
    LocalMux I__4187 (
            .O(N__20201),
            .I(N__20133));
    Span4Mux_v I__4186 (
            .O(N__20196),
            .I(N__20133));
    CascadeMux I__4185 (
            .O(N__20195),
            .I(N__20129));
    CascadeMux I__4184 (
            .O(N__20194),
            .I(N__20126));
    LocalMux I__4183 (
            .O(N__20183),
            .I(N__20115));
    LocalMux I__4182 (
            .O(N__20178),
            .I(N__20108));
    Span4Mux_h I__4181 (
            .O(N__20175),
            .I(N__20108));
    LocalMux I__4180 (
            .O(N__20172),
            .I(N__20108));
    LocalMux I__4179 (
            .O(N__20169),
            .I(N__20105));
    InMux I__4178 (
            .O(N__20168),
            .I(N__20090));
    InMux I__4177 (
            .O(N__20167),
            .I(N__20090));
    InMux I__4176 (
            .O(N__20166),
            .I(N__20090));
    InMux I__4175 (
            .O(N__20165),
            .I(N__20090));
    InMux I__4174 (
            .O(N__20164),
            .I(N__20090));
    InMux I__4173 (
            .O(N__20163),
            .I(N__20090));
    InMux I__4172 (
            .O(N__20162),
            .I(N__20090));
    LocalMux I__4171 (
            .O(N__20159),
            .I(N__20085));
    LocalMux I__4170 (
            .O(N__20156),
            .I(N__20085));
    LocalMux I__4169 (
            .O(N__20151),
            .I(N__20082));
    Span4Mux_h I__4168 (
            .O(N__20146),
            .I(N__20079));
    InMux I__4167 (
            .O(N__20145),
            .I(N__20076));
    Span4Mux_h I__4166 (
            .O(N__20140),
            .I(N__20071));
    Span4Mux_v I__4165 (
            .O(N__20133),
            .I(N__20071));
    InMux I__4164 (
            .O(N__20132),
            .I(N__20060));
    InMux I__4163 (
            .O(N__20129),
            .I(N__20060));
    InMux I__4162 (
            .O(N__20126),
            .I(N__20060));
    InMux I__4161 (
            .O(N__20125),
            .I(N__20060));
    InMux I__4160 (
            .O(N__20124),
            .I(N__20060));
    InMux I__4159 (
            .O(N__20123),
            .I(N__20051));
    InMux I__4158 (
            .O(N__20122),
            .I(N__20051));
    InMux I__4157 (
            .O(N__20121),
            .I(N__20051));
    InMux I__4156 (
            .O(N__20120),
            .I(N__20051));
    InMux I__4155 (
            .O(N__20119),
            .I(N__20046));
    InMux I__4154 (
            .O(N__20118),
            .I(N__20046));
    Span4Mux_h I__4153 (
            .O(N__20115),
            .I(N__20043));
    Span4Mux_v I__4152 (
            .O(N__20108),
            .I(N__20034));
    Span4Mux_h I__4151 (
            .O(N__20105),
            .I(N__20034));
    LocalMux I__4150 (
            .O(N__20090),
            .I(N__20034));
    Span4Mux_h I__4149 (
            .O(N__20085),
            .I(N__20034));
    Span12Mux_s11_v I__4148 (
            .O(N__20082),
            .I(N__20031));
    Odrv4 I__4147 (
            .O(N__20079),
            .I(\tok.T_0 ));
    LocalMux I__4146 (
            .O(N__20076),
            .I(\tok.T_0 ));
    Odrv4 I__4145 (
            .O(N__20071),
            .I(\tok.T_0 ));
    LocalMux I__4144 (
            .O(N__20060),
            .I(\tok.T_0 ));
    LocalMux I__4143 (
            .O(N__20051),
            .I(\tok.T_0 ));
    LocalMux I__4142 (
            .O(N__20046),
            .I(\tok.T_0 ));
    Odrv4 I__4141 (
            .O(N__20043),
            .I(\tok.T_0 ));
    Odrv4 I__4140 (
            .O(N__20034),
            .I(\tok.T_0 ));
    Odrv12 I__4139 (
            .O(N__20031),
            .I(\tok.T_0 ));
    InMux I__4138 (
            .O(N__20012),
            .I(N__20009));
    LocalMux I__4137 (
            .O(N__20009),
            .I(N__20006));
    Odrv4 I__4136 (
            .O(N__20006),
            .I(\tok.n10_adj_858 ));
    InMux I__4135 (
            .O(N__20003),
            .I(N__20000));
    LocalMux I__4134 (
            .O(N__20000),
            .I(N__19997));
    Span4Mux_h I__4133 (
            .O(N__19997),
            .I(N__19994));
    Span4Mux_h I__4132 (
            .O(N__19994),
            .I(N__19991));
    Odrv4 I__4131 (
            .O(N__19991),
            .I(\tok.table_rd_13 ));
    InMux I__4130 (
            .O(N__19988),
            .I(N__19985));
    LocalMux I__4129 (
            .O(N__19985),
            .I(N__19982));
    Odrv12 I__4128 (
            .O(N__19982),
            .I(\tok.n5_adj_732 ));
    InMux I__4127 (
            .O(N__19979),
            .I(N__19976));
    LocalMux I__4126 (
            .O(N__19976),
            .I(\tok.n12_adj_779 ));
    CascadeMux I__4125 (
            .O(N__19973),
            .I(\tok.n14_adj_776_cascade_ ));
    InMux I__4124 (
            .O(N__19970),
            .I(N__19967));
    LocalMux I__4123 (
            .O(N__19967),
            .I(\tok.n13_adj_780 ));
    CascadeMux I__4122 (
            .O(N__19964),
            .I(\tok.n20_adj_784_cascade_ ));
    InMux I__4121 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__4120 (
            .O(N__19958),
            .I(\tok.n9_adj_781 ));
    InMux I__4119 (
            .O(N__19955),
            .I(N__19952));
    LocalMux I__4118 (
            .O(N__19952),
            .I(N__19949));
    Odrv12 I__4117 (
            .O(N__19949),
            .I(\tok.n5_adj_713 ));
    InMux I__4116 (
            .O(N__19946),
            .I(N__19943));
    LocalMux I__4115 (
            .O(N__19943),
            .I(N__19940));
    Span4Mux_v I__4114 (
            .O(N__19940),
            .I(N__19937));
    Span4Mux_h I__4113 (
            .O(N__19937),
            .I(N__19934));
    Span4Mux_h I__4112 (
            .O(N__19934),
            .I(N__19931));
    Odrv4 I__4111 (
            .O(N__19931),
            .I(\tok.table_rd_15 ));
    InMux I__4110 (
            .O(N__19928),
            .I(N__19925));
    LocalMux I__4109 (
            .O(N__19925),
            .I(\tok.n16_adj_782 ));
    CascadeMux I__4108 (
            .O(N__19922),
            .I(\tok.n10_adj_700_cascade_ ));
    InMux I__4107 (
            .O(N__19919),
            .I(N__19916));
    LocalMux I__4106 (
            .O(N__19916),
            .I(\tok.n5536 ));
    InMux I__4105 (
            .O(N__19913),
            .I(N__19910));
    LocalMux I__4104 (
            .O(N__19910),
            .I(\tok.n11_adj_730 ));
    CascadeMux I__4103 (
            .O(N__19907),
            .I(\tok.n26_cascade_ ));
    CascadeMux I__4102 (
            .O(N__19904),
            .I(N__19898));
    InMux I__4101 (
            .O(N__19903),
            .I(N__19892));
    InMux I__4100 (
            .O(N__19902),
            .I(N__19889));
    InMux I__4099 (
            .O(N__19901),
            .I(N__19885));
    InMux I__4098 (
            .O(N__19898),
            .I(N__19882));
    InMux I__4097 (
            .O(N__19897),
            .I(N__19879));
    InMux I__4096 (
            .O(N__19896),
            .I(N__19876));
    InMux I__4095 (
            .O(N__19895),
            .I(N__19873));
    LocalMux I__4094 (
            .O(N__19892),
            .I(N__19870));
    LocalMux I__4093 (
            .O(N__19889),
            .I(N__19867));
    InMux I__4092 (
            .O(N__19888),
            .I(N__19864));
    LocalMux I__4091 (
            .O(N__19885),
            .I(N__19861));
    LocalMux I__4090 (
            .O(N__19882),
            .I(N__19856));
    LocalMux I__4089 (
            .O(N__19879),
            .I(N__19856));
    LocalMux I__4088 (
            .O(N__19876),
            .I(N__19853));
    LocalMux I__4087 (
            .O(N__19873),
            .I(N__19848));
    Span4Mux_h I__4086 (
            .O(N__19870),
            .I(N__19848));
    Span4Mux_v I__4085 (
            .O(N__19867),
            .I(N__19845));
    LocalMux I__4084 (
            .O(N__19864),
            .I(N__19842));
    Span4Mux_v I__4083 (
            .O(N__19861),
            .I(N__19839));
    Span4Mux_h I__4082 (
            .O(N__19856),
            .I(N__19836));
    Span4Mux_h I__4081 (
            .O(N__19853),
            .I(N__19831));
    Span4Mux_v I__4080 (
            .O(N__19848),
            .I(N__19831));
    Span4Mux_h I__4079 (
            .O(N__19845),
            .I(N__19828));
    Span4Mux_h I__4078 (
            .O(N__19842),
            .I(N__19823));
    Span4Mux_h I__4077 (
            .O(N__19839),
            .I(N__19823));
    Span4Mux_v I__4076 (
            .O(N__19836),
            .I(N__19818));
    Span4Mux_h I__4075 (
            .O(N__19831),
            .I(N__19818));
    Odrv4 I__4074 (
            .O(N__19828),
            .I(\tok.tc__7__N_134 ));
    Odrv4 I__4073 (
            .O(N__19823),
            .I(\tok.tc__7__N_134 ));
    Odrv4 I__4072 (
            .O(N__19818),
            .I(\tok.tc__7__N_134 ));
    InMux I__4071 (
            .O(N__19811),
            .I(N__19808));
    LocalMux I__4070 (
            .O(N__19808),
            .I(\tok.n25_adj_710 ));
    InMux I__4069 (
            .O(N__19805),
            .I(N__19802));
    LocalMux I__4068 (
            .O(N__19802),
            .I(N__19799));
    Odrv4 I__4067 (
            .O(N__19799),
            .I(\tok.n28_adj_708 ));
    InMux I__4066 (
            .O(N__19796),
            .I(N__19793));
    LocalMux I__4065 (
            .O(N__19793),
            .I(\tok.n27_adj_709 ));
    InMux I__4064 (
            .O(N__19790),
            .I(N__19787));
    LocalMux I__4063 (
            .O(N__19787),
            .I(N__19784));
    Span4Mux_v I__4062 (
            .O(N__19784),
            .I(N__19781));
    Span4Mux_h I__4061 (
            .O(N__19781),
            .I(N__19778));
    Odrv4 I__4060 (
            .O(N__19778),
            .I(\tok.n16_adj_810 ));
    CascadeMux I__4059 (
            .O(N__19775),
            .I(\tok.n14_adj_841_cascade_ ));
    InMux I__4058 (
            .O(N__19772),
            .I(N__19769));
    LocalMux I__4057 (
            .O(N__19769),
            .I(N__19766));
    Span4Mux_h I__4056 (
            .O(N__19766),
            .I(N__19763));
    Odrv4 I__4055 (
            .O(N__19763),
            .I(\tok.n5571 ));
    InMux I__4054 (
            .O(N__19760),
            .I(N__19757));
    LocalMux I__4053 (
            .O(N__19757),
            .I(\tok.n5569 ));
    InMux I__4052 (
            .O(N__19754),
            .I(N__19751));
    LocalMux I__4051 (
            .O(N__19751),
            .I(N__19748));
    Odrv4 I__4050 (
            .O(N__19748),
            .I(\tok.n45_adj_849 ));
    InMux I__4049 (
            .O(N__19745),
            .I(N__19739));
    InMux I__4048 (
            .O(N__19744),
            .I(N__19739));
    LocalMux I__4047 (
            .O(N__19739),
            .I(N__19735));
    InMux I__4046 (
            .O(N__19738),
            .I(N__19732));
    Span4Mux_v I__4045 (
            .O(N__19735),
            .I(N__19727));
    LocalMux I__4044 (
            .O(N__19732),
            .I(N__19727));
    Odrv4 I__4043 (
            .O(N__19727),
            .I(\tok.n4848 ));
    InMux I__4042 (
            .O(N__19724),
            .I(N__19721));
    LocalMux I__4041 (
            .O(N__19721),
            .I(N__19718));
    Span4Mux_h I__4040 (
            .O(N__19718),
            .I(N__19715));
    Span4Mux_h I__4039 (
            .O(N__19715),
            .I(N__19712));
    Odrv4 I__4038 (
            .O(N__19712),
            .I(\tok.table_rd_9 ));
    CascadeMux I__4037 (
            .O(N__19709),
            .I(\tok.n45_cascade_ ));
    InMux I__4036 (
            .O(N__19706),
            .I(N__19703));
    LocalMux I__4035 (
            .O(N__19703),
            .I(\tok.n39 ));
    InMux I__4034 (
            .O(N__19700),
            .I(N__19694));
    InMux I__4033 (
            .O(N__19699),
            .I(N__19694));
    LocalMux I__4032 (
            .O(N__19694),
            .I(N__19690));
    InMux I__4031 (
            .O(N__19693),
            .I(N__19687));
    Span4Mux_v I__4030 (
            .O(N__19690),
            .I(N__19682));
    LocalMux I__4029 (
            .O(N__19687),
            .I(N__19682));
    Span4Mux_h I__4028 (
            .O(N__19682),
            .I(N__19677));
    InMux I__4027 (
            .O(N__19681),
            .I(N__19672));
    InMux I__4026 (
            .O(N__19680),
            .I(N__19672));
    Odrv4 I__4025 (
            .O(N__19677),
            .I(\tok.n11_adj_680 ));
    LocalMux I__4024 (
            .O(N__19672),
            .I(\tok.n11_adj_680 ));
    InMux I__4023 (
            .O(N__19667),
            .I(N__19664));
    LocalMux I__4022 (
            .O(N__19664),
            .I(N__19661));
    Span4Mux_v I__4021 (
            .O(N__19661),
            .I(N__19658));
    Span4Mux_h I__4020 (
            .O(N__19658),
            .I(N__19655));
    Span4Mux_h I__4019 (
            .O(N__19655),
            .I(N__19652));
    Span4Mux_s0_h I__4018 (
            .O(N__19652),
            .I(N__19649));
    Odrv4 I__4017 (
            .O(N__19649),
            .I(\tok.table_rd_10 ));
    CascadeMux I__4016 (
            .O(N__19646),
            .I(N__19643));
    InMux I__4015 (
            .O(N__19643),
            .I(N__19637));
    InMux I__4014 (
            .O(N__19642),
            .I(N__19637));
    LocalMux I__4013 (
            .O(N__19637),
            .I(\tok.n14_adj_679 ));
    InMux I__4012 (
            .O(N__19634),
            .I(N__19631));
    LocalMux I__4011 (
            .O(N__19631),
            .I(\tok.n45_adj_696 ));
    CascadeMux I__4010 (
            .O(N__19628),
            .I(\tok.n39_adj_697_cascade_ ));
    InMux I__4009 (
            .O(N__19625),
            .I(N__19622));
    LocalMux I__4008 (
            .O(N__19622),
            .I(\tok.n5_adj_734 ));
    InMux I__4007 (
            .O(N__19619),
            .I(\tok.n4795 ));
    InMux I__4006 (
            .O(N__19616),
            .I(\tok.n4796 ));
    InMux I__4005 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__4004 (
            .O(N__19610),
            .I(N__19607));
    Odrv4 I__4003 (
            .O(N__19607),
            .I(\tok.n5_adj_716 ));
    InMux I__4002 (
            .O(N__19604),
            .I(\tok.n4797 ));
    InMux I__4001 (
            .O(N__19601),
            .I(N__19579));
    InMux I__4000 (
            .O(N__19600),
            .I(N__19579));
    InMux I__3999 (
            .O(N__19599),
            .I(N__19579));
    InMux I__3998 (
            .O(N__19598),
            .I(N__19568));
    InMux I__3997 (
            .O(N__19597),
            .I(N__19568));
    InMux I__3996 (
            .O(N__19596),
            .I(N__19568));
    InMux I__3995 (
            .O(N__19595),
            .I(N__19568));
    InMux I__3994 (
            .O(N__19594),
            .I(N__19568));
    InMux I__3993 (
            .O(N__19593),
            .I(N__19561));
    InMux I__3992 (
            .O(N__19592),
            .I(N__19561));
    InMux I__3991 (
            .O(N__19591),
            .I(N__19561));
    InMux I__3990 (
            .O(N__19590),
            .I(N__19550));
    InMux I__3989 (
            .O(N__19589),
            .I(N__19550));
    InMux I__3988 (
            .O(N__19588),
            .I(N__19550));
    InMux I__3987 (
            .O(N__19587),
            .I(N__19550));
    InMux I__3986 (
            .O(N__19586),
            .I(N__19550));
    LocalMux I__3985 (
            .O(N__19579),
            .I(N__19545));
    LocalMux I__3984 (
            .O(N__19568),
            .I(N__19545));
    LocalMux I__3983 (
            .O(N__19561),
            .I(N__19540));
    LocalMux I__3982 (
            .O(N__19550),
            .I(N__19540));
    Span4Mux_v I__3981 (
            .O(N__19545),
            .I(N__19537));
    Span4Mux_v I__3980 (
            .O(N__19540),
            .I(N__19534));
    Span4Mux_h I__3979 (
            .O(N__19537),
            .I(N__19529));
    Span4Mux_h I__3978 (
            .O(N__19534),
            .I(N__19529));
    Odrv4 I__3977 (
            .O(N__19529),
            .I(\tok.n399 ));
    InMux I__3976 (
            .O(N__19526),
            .I(\tok.n4798 ));
    InMux I__3975 (
            .O(N__19523),
            .I(N__19520));
    LocalMux I__3974 (
            .O(N__19520),
            .I(\tok.n8_adj_837 ));
    InMux I__3973 (
            .O(N__19517),
            .I(N__19514));
    LocalMux I__3972 (
            .O(N__19514),
            .I(\tok.n5574 ));
    InMux I__3971 (
            .O(N__19511),
            .I(N__19507));
    InMux I__3970 (
            .O(N__19510),
            .I(N__19504));
    LocalMux I__3969 (
            .O(N__19507),
            .I(\tok.n5334 ));
    LocalMux I__3968 (
            .O(N__19504),
            .I(\tok.n5334 ));
    InMux I__3967 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__3966 (
            .O(N__19496),
            .I(N__19493));
    Span4Mux_v I__3965 (
            .O(N__19493),
            .I(N__19490));
    Odrv4 I__3964 (
            .O(N__19490),
            .I(\tok.n5254 ));
    CascadeMux I__3963 (
            .O(N__19487),
            .I(\tok.n5414_cascade_ ));
    InMux I__3962 (
            .O(N__19484),
            .I(N__19481));
    LocalMux I__3961 (
            .O(N__19481),
            .I(\tok.n8_adj_767 ));
    CascadeMux I__3960 (
            .O(N__19478),
            .I(\tok.n904_cascade_ ));
    InMux I__3959 (
            .O(N__19475),
            .I(N__19472));
    LocalMux I__3958 (
            .O(N__19472),
            .I(N__19469));
    Span4Mux_v I__3957 (
            .O(N__19469),
            .I(N__19466));
    Span4Mux_s2_v I__3956 (
            .O(N__19466),
            .I(N__19463));
    Odrv4 I__3955 (
            .O(N__19463),
            .I(\tok.n11_adj_840 ));
    CascadeMux I__3954 (
            .O(N__19460),
            .I(\tok.n5346_cascade_ ));
    InMux I__3953 (
            .O(N__19457),
            .I(N__19454));
    LocalMux I__3952 (
            .O(N__19454),
            .I(N__19451));
    Sp12to4 I__3951 (
            .O(N__19451),
            .I(N__19448));
    Odrv12 I__3950 (
            .O(N__19448),
            .I(\tok.n4_adj_806 ));
    InMux I__3949 (
            .O(N__19445),
            .I(\tok.n4786 ));
    InMux I__3948 (
            .O(N__19442),
            .I(N__19439));
    LocalMux I__3947 (
            .O(N__19439),
            .I(\tok.n5564 ));
    InMux I__3946 (
            .O(N__19436),
            .I(\tok.n4787 ));
    InMux I__3945 (
            .O(N__19433),
            .I(\tok.n4788 ));
    CascadeMux I__3944 (
            .O(N__19430),
            .I(N__19427));
    InMux I__3943 (
            .O(N__19427),
            .I(N__19424));
    LocalMux I__3942 (
            .O(N__19424),
            .I(\tok.n5554 ));
    InMux I__3941 (
            .O(N__19421),
            .I(\tok.n4789 ));
    CascadeMux I__3940 (
            .O(N__19418),
            .I(N__19415));
    InMux I__3939 (
            .O(N__19415),
            .I(N__19412));
    LocalMux I__3938 (
            .O(N__19412),
            .I(N__19409));
    Odrv12 I__3937 (
            .O(N__19409),
            .I(\tok.n5549 ));
    InMux I__3936 (
            .O(N__19406),
            .I(\tok.n4790 ));
    InMux I__3935 (
            .O(N__19403),
            .I(bfn_8_8_0_));
    InMux I__3934 (
            .O(N__19400),
            .I(\tok.n4792 ));
    InMux I__3933 (
            .O(N__19397),
            .I(\tok.n4793 ));
    InMux I__3932 (
            .O(N__19394),
            .I(\tok.n4794 ));
    CascadeMux I__3931 (
            .O(N__19391),
            .I(\tok.n13_adj_654_cascade_ ));
    InMux I__3930 (
            .O(N__19388),
            .I(N__19385));
    LocalMux I__3929 (
            .O(N__19385),
            .I(\tok.n5547 ));
    CascadeMux I__3928 (
            .O(N__19382),
            .I(\tok.n5546_cascade_ ));
    InMux I__3927 (
            .O(N__19379),
            .I(N__19376));
    LocalMux I__3926 (
            .O(N__19376),
            .I(N__19373));
    Span4Mux_h I__3925 (
            .O(N__19373),
            .I(N__19370));
    Odrv4 I__3924 (
            .O(N__19370),
            .I(\tok.n14 ));
    InMux I__3923 (
            .O(N__19367),
            .I(N__19364));
    LocalMux I__3922 (
            .O(N__19364),
            .I(\tok.n17 ));
    CascadeMux I__3921 (
            .O(N__19361),
            .I(\tok.n13_adj_641_cascade_ ));
    InMux I__3920 (
            .O(N__19358),
            .I(N__19355));
    LocalMux I__3919 (
            .O(N__19355),
            .I(\tok.n5552 ));
    CascadeMux I__3918 (
            .O(N__19352),
            .I(\tok.n5551_cascade_ ));
    InMux I__3917 (
            .O(N__19349),
            .I(N__19346));
    LocalMux I__3916 (
            .O(N__19346),
            .I(N__19343));
    Odrv4 I__3915 (
            .O(N__19343),
            .I(\tok.n5465 ));
    InMux I__3914 (
            .O(N__19340),
            .I(\tok.n4784 ));
    InMux I__3913 (
            .O(N__19337),
            .I(\tok.n4785 ));
    CascadeMux I__3912 (
            .O(N__19334),
            .I(N__19330));
    InMux I__3911 (
            .O(N__19333),
            .I(N__19325));
    InMux I__3910 (
            .O(N__19330),
            .I(N__19325));
    LocalMux I__3909 (
            .O(N__19325),
            .I(N__19320));
    InMux I__3908 (
            .O(N__19324),
            .I(N__19315));
    InMux I__3907 (
            .O(N__19323),
            .I(N__19315));
    Span12Mux_s4_v I__3906 (
            .O(N__19320),
            .I(N__19312));
    LocalMux I__3905 (
            .O(N__19315),
            .I(\tok.n9_adj_786 ));
    Odrv12 I__3904 (
            .O(N__19312),
            .I(\tok.n9_adj_786 ));
    InMux I__3903 (
            .O(N__19307),
            .I(N__19304));
    LocalMux I__3902 (
            .O(N__19304),
            .I(N__19301));
    Span4Mux_v I__3901 (
            .O(N__19301),
            .I(N__19297));
    CascadeMux I__3900 (
            .O(N__19300),
            .I(N__19294));
    Span4Mux_h I__3899 (
            .O(N__19297),
            .I(N__19291));
    InMux I__3898 (
            .O(N__19294),
            .I(N__19288));
    Odrv4 I__3897 (
            .O(N__19291),
            .I(\tok.table_rd_7 ));
    LocalMux I__3896 (
            .O(N__19288),
            .I(\tok.table_rd_7 ));
    CascadeMux I__3895 (
            .O(N__19283),
            .I(\tok.n5548_cascade_ ));
    CascadeMux I__3894 (
            .O(N__19280),
            .I(\tok.n285_cascade_ ));
    InMux I__3893 (
            .O(N__19277),
            .I(N__19274));
    LocalMux I__3892 (
            .O(N__19274),
            .I(N__19271));
    Span4Mux_v I__3891 (
            .O(N__19271),
            .I(N__19268));
    Span4Mux_h I__3890 (
            .O(N__19268),
            .I(N__19265));
    Odrv4 I__3889 (
            .O(N__19265),
            .I(\tok.n12_adj_824 ));
    CascadeMux I__3888 (
            .O(N__19262),
            .I(\tok.n1_adj_862_cascade_ ));
    InMux I__3887 (
            .O(N__19259),
            .I(N__19252));
    InMux I__3886 (
            .O(N__19258),
            .I(N__19247));
    InMux I__3885 (
            .O(N__19257),
            .I(N__19247));
    InMux I__3884 (
            .O(N__19256),
            .I(N__19241));
    CascadeMux I__3883 (
            .O(N__19255),
            .I(N__19233));
    LocalMux I__3882 (
            .O(N__19252),
            .I(N__19227));
    LocalMux I__3881 (
            .O(N__19247),
            .I(N__19227));
    InMux I__3880 (
            .O(N__19246),
            .I(N__19224));
    InMux I__3879 (
            .O(N__19245),
            .I(N__19221));
    InMux I__3878 (
            .O(N__19244),
            .I(N__19218));
    LocalMux I__3877 (
            .O(N__19241),
            .I(N__19211));
    InMux I__3876 (
            .O(N__19240),
            .I(N__19208));
    InMux I__3875 (
            .O(N__19239),
            .I(N__19205));
    InMux I__3874 (
            .O(N__19238),
            .I(N__19200));
    InMux I__3873 (
            .O(N__19237),
            .I(N__19200));
    InMux I__3872 (
            .O(N__19236),
            .I(N__19191));
    InMux I__3871 (
            .O(N__19233),
            .I(N__19191));
    InMux I__3870 (
            .O(N__19232),
            .I(N__19191));
    Span4Mux_v I__3869 (
            .O(N__19227),
            .I(N__19186));
    LocalMux I__3868 (
            .O(N__19224),
            .I(N__19186));
    LocalMux I__3867 (
            .O(N__19221),
            .I(N__19183));
    LocalMux I__3866 (
            .O(N__19218),
            .I(N__19180));
    InMux I__3865 (
            .O(N__19217),
            .I(N__19175));
    InMux I__3864 (
            .O(N__19216),
            .I(N__19175));
    InMux I__3863 (
            .O(N__19215),
            .I(N__19172));
    InMux I__3862 (
            .O(N__19214),
            .I(N__19169));
    Span4Mux_v I__3861 (
            .O(N__19211),
            .I(N__19163));
    LocalMux I__3860 (
            .O(N__19208),
            .I(N__19158));
    LocalMux I__3859 (
            .O(N__19205),
            .I(N__19158));
    LocalMux I__3858 (
            .O(N__19200),
            .I(N__19155));
    InMux I__3857 (
            .O(N__19199),
            .I(N__19148));
    InMux I__3856 (
            .O(N__19198),
            .I(N__19148));
    LocalMux I__3855 (
            .O(N__19191),
            .I(N__19143));
    Span4Mux_h I__3854 (
            .O(N__19186),
            .I(N__19143));
    Span4Mux_h I__3853 (
            .O(N__19183),
            .I(N__19140));
    Span4Mux_v I__3852 (
            .O(N__19180),
            .I(N__19135));
    LocalMux I__3851 (
            .O(N__19175),
            .I(N__19135));
    LocalMux I__3850 (
            .O(N__19172),
            .I(N__19130));
    LocalMux I__3849 (
            .O(N__19169),
            .I(N__19130));
    InMux I__3848 (
            .O(N__19168),
            .I(N__19125));
    InMux I__3847 (
            .O(N__19167),
            .I(N__19125));
    InMux I__3846 (
            .O(N__19166),
            .I(N__19122));
    Span4Mux_v I__3845 (
            .O(N__19163),
            .I(N__19119));
    Span4Mux_v I__3844 (
            .O(N__19158),
            .I(N__19116));
    Span12Mux_s10_v I__3843 (
            .O(N__19155),
            .I(N__19113));
    InMux I__3842 (
            .O(N__19154),
            .I(N__19110));
    InMux I__3841 (
            .O(N__19153),
            .I(N__19107));
    LocalMux I__3840 (
            .O(N__19148),
            .I(N__19102));
    Span4Mux_v I__3839 (
            .O(N__19143),
            .I(N__19102));
    Span4Mux_v I__3838 (
            .O(N__19140),
            .I(N__19097));
    Span4Mux_h I__3837 (
            .O(N__19135),
            .I(N__19097));
    Span4Mux_s3_v I__3836 (
            .O(N__19130),
            .I(N__19092));
    LocalMux I__3835 (
            .O(N__19125),
            .I(N__19092));
    LocalMux I__3834 (
            .O(N__19122),
            .I(\tok.T_6 ));
    Odrv4 I__3833 (
            .O(N__19119),
            .I(\tok.T_6 ));
    Odrv4 I__3832 (
            .O(N__19116),
            .I(\tok.T_6 ));
    Odrv12 I__3831 (
            .O(N__19113),
            .I(\tok.T_6 ));
    LocalMux I__3830 (
            .O(N__19110),
            .I(\tok.T_6 ));
    LocalMux I__3829 (
            .O(N__19107),
            .I(\tok.T_6 ));
    Odrv4 I__3828 (
            .O(N__19102),
            .I(\tok.T_6 ));
    Odrv4 I__3827 (
            .O(N__19097),
            .I(\tok.T_6 ));
    Odrv4 I__3826 (
            .O(N__19092),
            .I(\tok.T_6 ));
    CascadeMux I__3825 (
            .O(N__19073),
            .I(N__19067));
    InMux I__3824 (
            .O(N__19072),
            .I(N__19061));
    InMux I__3823 (
            .O(N__19071),
            .I(N__19061));
    InMux I__3822 (
            .O(N__19070),
            .I(N__19039));
    InMux I__3821 (
            .O(N__19067),
            .I(N__19032));
    InMux I__3820 (
            .O(N__19066),
            .I(N__19032));
    LocalMux I__3819 (
            .O(N__19061),
            .I(N__19029));
    InMux I__3818 (
            .O(N__19060),
            .I(N__19024));
    InMux I__3817 (
            .O(N__19059),
            .I(N__19024));
    InMux I__3816 (
            .O(N__19058),
            .I(N__19019));
    InMux I__3815 (
            .O(N__19057),
            .I(N__19019));
    InMux I__3814 (
            .O(N__19056),
            .I(N__19010));
    InMux I__3813 (
            .O(N__19055),
            .I(N__19010));
    InMux I__3812 (
            .O(N__19054),
            .I(N__19010));
    InMux I__3811 (
            .O(N__19053),
            .I(N__19007));
    InMux I__3810 (
            .O(N__19052),
            .I(N__19004));
    InMux I__3809 (
            .O(N__19051),
            .I(N__18999));
    InMux I__3808 (
            .O(N__19050),
            .I(N__18999));
    InMux I__3807 (
            .O(N__19049),
            .I(N__18994));
    InMux I__3806 (
            .O(N__19048),
            .I(N__18994));
    InMux I__3805 (
            .O(N__19047),
            .I(N__18987));
    InMux I__3804 (
            .O(N__19046),
            .I(N__18987));
    InMux I__3803 (
            .O(N__19045),
            .I(N__18987));
    InMux I__3802 (
            .O(N__19044),
            .I(N__18984));
    CascadeMux I__3801 (
            .O(N__19043),
            .I(N__18980));
    InMux I__3800 (
            .O(N__19042),
            .I(N__18976));
    LocalMux I__3799 (
            .O(N__19039),
            .I(N__18973));
    InMux I__3798 (
            .O(N__19038),
            .I(N__18970));
    InMux I__3797 (
            .O(N__19037),
            .I(N__18967));
    LocalMux I__3796 (
            .O(N__19032),
            .I(N__18964));
    Span4Mux_v I__3795 (
            .O(N__19029),
            .I(N__18955));
    LocalMux I__3794 (
            .O(N__19024),
            .I(N__18955));
    LocalMux I__3793 (
            .O(N__19019),
            .I(N__18955));
    InMux I__3792 (
            .O(N__19018),
            .I(N__18950));
    InMux I__3791 (
            .O(N__19017),
            .I(N__18950));
    LocalMux I__3790 (
            .O(N__19010),
            .I(N__18947));
    LocalMux I__3789 (
            .O(N__19007),
            .I(N__18942));
    LocalMux I__3788 (
            .O(N__19004),
            .I(N__18942));
    LocalMux I__3787 (
            .O(N__18999),
            .I(N__18937));
    LocalMux I__3786 (
            .O(N__18994),
            .I(N__18937));
    LocalMux I__3785 (
            .O(N__18987),
            .I(N__18932));
    LocalMux I__3784 (
            .O(N__18984),
            .I(N__18932));
    InMux I__3783 (
            .O(N__18983),
            .I(N__18925));
    InMux I__3782 (
            .O(N__18980),
            .I(N__18925));
    InMux I__3781 (
            .O(N__18979),
            .I(N__18925));
    LocalMux I__3780 (
            .O(N__18976),
            .I(N__18921));
    Span4Mux_h I__3779 (
            .O(N__18973),
            .I(N__18918));
    LocalMux I__3778 (
            .O(N__18970),
            .I(N__18915));
    LocalMux I__3777 (
            .O(N__18967),
            .I(N__18910));
    Span4Mux_v I__3776 (
            .O(N__18964),
            .I(N__18910));
    CascadeMux I__3775 (
            .O(N__18963),
            .I(N__18905));
    CascadeMux I__3774 (
            .O(N__18962),
            .I(N__18902));
    Span4Mux_h I__3773 (
            .O(N__18955),
            .I(N__18897));
    LocalMux I__3772 (
            .O(N__18950),
            .I(N__18897));
    Span4Mux_s3_h I__3771 (
            .O(N__18947),
            .I(N__18894));
    Span4Mux_v I__3770 (
            .O(N__18942),
            .I(N__18891));
    Span4Mux_v I__3769 (
            .O(N__18937),
            .I(N__18884));
    Span4Mux_v I__3768 (
            .O(N__18932),
            .I(N__18884));
    LocalMux I__3767 (
            .O(N__18925),
            .I(N__18884));
    InMux I__3766 (
            .O(N__18924),
            .I(N__18881));
    Span4Mux_h I__3765 (
            .O(N__18921),
            .I(N__18876));
    Span4Mux_v I__3764 (
            .O(N__18918),
            .I(N__18876));
    Span4Mux_v I__3763 (
            .O(N__18915),
            .I(N__18871));
    Span4Mux_h I__3762 (
            .O(N__18910),
            .I(N__18871));
    InMux I__3761 (
            .O(N__18909),
            .I(N__18866));
    InMux I__3760 (
            .O(N__18908),
            .I(N__18866));
    InMux I__3759 (
            .O(N__18905),
            .I(N__18863));
    InMux I__3758 (
            .O(N__18902),
            .I(N__18860));
    Span4Mux_v I__3757 (
            .O(N__18897),
            .I(N__18851));
    Span4Mux_v I__3756 (
            .O(N__18894),
            .I(N__18851));
    Span4Mux_h I__3755 (
            .O(N__18891),
            .I(N__18851));
    Span4Mux_h I__3754 (
            .O(N__18884),
            .I(N__18851));
    LocalMux I__3753 (
            .O(N__18881),
            .I(\tok.T_4 ));
    Odrv4 I__3752 (
            .O(N__18876),
            .I(\tok.T_4 ));
    Odrv4 I__3751 (
            .O(N__18871),
            .I(\tok.T_4 ));
    LocalMux I__3750 (
            .O(N__18866),
            .I(\tok.T_4 ));
    LocalMux I__3749 (
            .O(N__18863),
            .I(\tok.T_4 ));
    LocalMux I__3748 (
            .O(N__18860),
            .I(\tok.T_4 ));
    Odrv4 I__3747 (
            .O(N__18851),
            .I(\tok.T_4 ));
    CascadeMux I__3746 (
            .O(N__18836),
            .I(N__18827));
    InMux I__3745 (
            .O(N__18835),
            .I(N__18822));
    InMux I__3744 (
            .O(N__18834),
            .I(N__18822));
    InMux I__3743 (
            .O(N__18833),
            .I(N__18819));
    InMux I__3742 (
            .O(N__18832),
            .I(N__18808));
    InMux I__3741 (
            .O(N__18831),
            .I(N__18808));
    InMux I__3740 (
            .O(N__18830),
            .I(N__18808));
    InMux I__3739 (
            .O(N__18827),
            .I(N__18805));
    LocalMux I__3738 (
            .O(N__18822),
            .I(N__18799));
    LocalMux I__3737 (
            .O(N__18819),
            .I(N__18799));
    InMux I__3736 (
            .O(N__18818),
            .I(N__18792));
    InMux I__3735 (
            .O(N__18817),
            .I(N__18792));
    InMux I__3734 (
            .O(N__18816),
            .I(N__18792));
    CascadeMux I__3733 (
            .O(N__18815),
            .I(N__18788));
    LocalMux I__3732 (
            .O(N__18808),
            .I(N__18785));
    LocalMux I__3731 (
            .O(N__18805),
            .I(N__18782));
    InMux I__3730 (
            .O(N__18804),
            .I(N__18779));
    Span4Mux_v I__3729 (
            .O(N__18799),
            .I(N__18774));
    LocalMux I__3728 (
            .O(N__18792),
            .I(N__18771));
    InMux I__3727 (
            .O(N__18791),
            .I(N__18766));
    InMux I__3726 (
            .O(N__18788),
            .I(N__18766));
    Span4Mux_v I__3725 (
            .O(N__18785),
            .I(N__18762));
    Span4Mux_v I__3724 (
            .O(N__18782),
            .I(N__18758));
    LocalMux I__3723 (
            .O(N__18779),
            .I(N__18755));
    InMux I__3722 (
            .O(N__18778),
            .I(N__18750));
    InMux I__3721 (
            .O(N__18777),
            .I(N__18750));
    Span4Mux_v I__3720 (
            .O(N__18774),
            .I(N__18743));
    Span4Mux_v I__3719 (
            .O(N__18771),
            .I(N__18743));
    LocalMux I__3718 (
            .O(N__18766),
            .I(N__18743));
    InMux I__3717 (
            .O(N__18765),
            .I(N__18740));
    Span4Mux_h I__3716 (
            .O(N__18762),
            .I(N__18737));
    InMux I__3715 (
            .O(N__18761),
            .I(N__18734));
    Span4Mux_v I__3714 (
            .O(N__18758),
            .I(N__18727));
    Span4Mux_s3_v I__3713 (
            .O(N__18755),
            .I(N__18727));
    LocalMux I__3712 (
            .O(N__18750),
            .I(N__18727));
    Span4Mux_h I__3711 (
            .O(N__18743),
            .I(N__18724));
    LocalMux I__3710 (
            .O(N__18740),
            .I(\tok.T_5 ));
    Odrv4 I__3709 (
            .O(N__18737),
            .I(\tok.T_5 ));
    LocalMux I__3708 (
            .O(N__18734),
            .I(\tok.T_5 ));
    Odrv4 I__3707 (
            .O(N__18727),
            .I(\tok.T_5 ));
    Odrv4 I__3706 (
            .O(N__18724),
            .I(\tok.T_5 ));
    CascadeMux I__3705 (
            .O(N__18713),
            .I(\tok.n6_adj_650_cascade_ ));
    InMux I__3704 (
            .O(N__18710),
            .I(N__18704));
    InMux I__3703 (
            .O(N__18709),
            .I(N__18704));
    LocalMux I__3702 (
            .O(N__18704),
            .I(\tok.A_stk.tail_68 ));
    InMux I__3701 (
            .O(N__18701),
            .I(N__18695));
    InMux I__3700 (
            .O(N__18700),
            .I(N__18695));
    LocalMux I__3699 (
            .O(N__18695),
            .I(\tok.A_stk.tail_52 ));
    InMux I__3698 (
            .O(N__18692),
            .I(N__18686));
    InMux I__3697 (
            .O(N__18691),
            .I(N__18686));
    LocalMux I__3696 (
            .O(N__18686),
            .I(\tok.A_stk.tail_36 ));
    InMux I__3695 (
            .O(N__18683),
            .I(N__18679));
    CascadeMux I__3694 (
            .O(N__18682),
            .I(N__18676));
    LocalMux I__3693 (
            .O(N__18679),
            .I(N__18673));
    InMux I__3692 (
            .O(N__18676),
            .I(N__18670));
    Odrv4 I__3691 (
            .O(N__18673),
            .I(tail_119));
    LocalMux I__3690 (
            .O(N__18670),
            .I(tail_119));
    InMux I__3689 (
            .O(N__18665),
            .I(N__18661));
    InMux I__3688 (
            .O(N__18664),
            .I(N__18658));
    LocalMux I__3687 (
            .O(N__18661),
            .I(\tok.A_stk.tail_20 ));
    LocalMux I__3686 (
            .O(N__18658),
            .I(\tok.A_stk.tail_20 ));
    InMux I__3685 (
            .O(N__18653),
            .I(N__18649));
    InMux I__3684 (
            .O(N__18652),
            .I(N__18646));
    LocalMux I__3683 (
            .O(N__18649),
            .I(tail_103));
    LocalMux I__3682 (
            .O(N__18646),
            .I(tail_103));
    CascadeMux I__3681 (
            .O(N__18641),
            .I(N__18638));
    InMux I__3680 (
            .O(N__18638),
            .I(N__18632));
    InMux I__3679 (
            .O(N__18637),
            .I(N__18632));
    LocalMux I__3678 (
            .O(N__18632),
            .I(\tok.A_stk.tail_71 ));
    InMux I__3677 (
            .O(N__18629),
            .I(N__18625));
    InMux I__3676 (
            .O(N__18628),
            .I(N__18622));
    LocalMux I__3675 (
            .O(N__18625),
            .I(\tok.A_stk.tail_87 ));
    LocalMux I__3674 (
            .O(N__18622),
            .I(\tok.A_stk.tail_87 ));
    InMux I__3673 (
            .O(N__18617),
            .I(N__18613));
    InMux I__3672 (
            .O(N__18616),
            .I(N__18610));
    LocalMux I__3671 (
            .O(N__18613),
            .I(tail_120));
    LocalMux I__3670 (
            .O(N__18610),
            .I(tail_120));
    InMux I__3669 (
            .O(N__18605),
            .I(N__18599));
    InMux I__3668 (
            .O(N__18604),
            .I(N__18599));
    LocalMux I__3667 (
            .O(N__18599),
            .I(\tok.A_stk.tail_88 ));
    InMux I__3666 (
            .O(N__18596),
            .I(N__18593));
    LocalMux I__3665 (
            .O(N__18593),
            .I(N__18589));
    InMux I__3664 (
            .O(N__18592),
            .I(N__18586));
    Odrv4 I__3663 (
            .O(N__18589),
            .I(tail_104));
    LocalMux I__3662 (
            .O(N__18586),
            .I(tail_104));
    InMux I__3661 (
            .O(N__18581),
            .I(N__18575));
    InMux I__3660 (
            .O(N__18580),
            .I(N__18575));
    LocalMux I__3659 (
            .O(N__18575),
            .I(\tok.A_stk.tail_41 ));
    InMux I__3658 (
            .O(N__18572),
            .I(N__18566));
    InMux I__3657 (
            .O(N__18571),
            .I(N__18566));
    LocalMux I__3656 (
            .O(N__18566),
            .I(\tok.A_stk.tail_25 ));
    CascadeMux I__3655 (
            .O(N__18563),
            .I(N__18560));
    InMux I__3654 (
            .O(N__18560),
            .I(N__18554));
    InMux I__3653 (
            .O(N__18559),
            .I(N__18554));
    LocalMux I__3652 (
            .O(N__18554),
            .I(\tok.A_stk.tail_9 ));
    CascadeMux I__3651 (
            .O(N__18551),
            .I(N__18547));
    InMux I__3650 (
            .O(N__18550),
            .I(N__18544));
    InMux I__3649 (
            .O(N__18547),
            .I(N__18541));
    LocalMux I__3648 (
            .O(N__18544),
            .I(tail_115));
    LocalMux I__3647 (
            .O(N__18541),
            .I(tail_115));
    InMux I__3646 (
            .O(N__18536),
            .I(N__18532));
    InMux I__3645 (
            .O(N__18535),
            .I(N__18529));
    LocalMux I__3644 (
            .O(N__18532),
            .I(tail_99));
    LocalMux I__3643 (
            .O(N__18529),
            .I(tail_99));
    InMux I__3642 (
            .O(N__18524),
            .I(N__18520));
    InMux I__3641 (
            .O(N__18523),
            .I(N__18517));
    LocalMux I__3640 (
            .O(N__18520),
            .I(\tok.A_stk.tail_84 ));
    LocalMux I__3639 (
            .O(N__18517),
            .I(\tok.A_stk.tail_84 ));
    InMux I__3638 (
            .O(N__18512),
            .I(\tok.n4765 ));
    CascadeMux I__3637 (
            .O(N__18509),
            .I(N__18506));
    InMux I__3636 (
            .O(N__18506),
            .I(N__18503));
    LocalMux I__3635 (
            .O(N__18503),
            .I(N__18500));
    Sp12to4 I__3634 (
            .O(N__18500),
            .I(N__18497));
    Odrv12 I__3633 (
            .O(N__18497),
            .I(\tok.n210 ));
    InMux I__3632 (
            .O(N__18494),
            .I(\tok.n4766 ));
    InMux I__3631 (
            .O(N__18491),
            .I(\tok.n4767 ));
    InMux I__3630 (
            .O(N__18488),
            .I(bfn_7_14_0_));
    InMux I__3629 (
            .O(N__18485),
            .I(N__18482));
    LocalMux I__3628 (
            .O(N__18482),
            .I(N__18478));
    InMux I__3627 (
            .O(N__18481),
            .I(N__18475));
    Odrv4 I__3626 (
            .O(N__18478),
            .I(tail_121));
    LocalMux I__3625 (
            .O(N__18475),
            .I(tail_121));
    InMux I__3624 (
            .O(N__18470),
            .I(N__18467));
    LocalMux I__3623 (
            .O(N__18467),
            .I(N__18464));
    Span4Mux_h I__3622 (
            .O(N__18464),
            .I(N__18460));
    InMux I__3621 (
            .O(N__18463),
            .I(N__18457));
    Odrv4 I__3620 (
            .O(N__18460),
            .I(tail_105));
    LocalMux I__3619 (
            .O(N__18457),
            .I(tail_105));
    InMux I__3618 (
            .O(N__18452),
            .I(N__18446));
    InMux I__3617 (
            .O(N__18451),
            .I(N__18446));
    LocalMux I__3616 (
            .O(N__18446),
            .I(\tok.A_stk.tail_89 ));
    InMux I__3615 (
            .O(N__18443),
            .I(N__18437));
    InMux I__3614 (
            .O(N__18442),
            .I(N__18437));
    LocalMux I__3613 (
            .O(N__18437),
            .I(\tok.A_stk.tail_73 ));
    InMux I__3612 (
            .O(N__18434),
            .I(N__18428));
    InMux I__3611 (
            .O(N__18433),
            .I(N__18428));
    LocalMux I__3610 (
            .O(N__18428),
            .I(\tok.A_stk.tail_57 ));
    CascadeMux I__3609 (
            .O(N__18425),
            .I(\tok.n82_cascade_ ));
    InMux I__3608 (
            .O(N__18422),
            .I(N__18415));
    InMux I__3607 (
            .O(N__18421),
            .I(N__18415));
    InMux I__3606 (
            .O(N__18420),
            .I(N__18411));
    LocalMux I__3605 (
            .O(N__18415),
            .I(N__18408));
    InMux I__3604 (
            .O(N__18414),
            .I(N__18405));
    LocalMux I__3603 (
            .O(N__18411),
            .I(\tok.n878 ));
    Odrv4 I__3602 (
            .O(N__18408),
            .I(\tok.n878 ));
    LocalMux I__3601 (
            .O(N__18405),
            .I(\tok.n878 ));
    InMux I__3600 (
            .O(N__18398),
            .I(N__18395));
    LocalMux I__3599 (
            .O(N__18395),
            .I(N__18392));
    Span4Mux_h I__3598 (
            .O(N__18392),
            .I(N__18389));
    Odrv4 I__3597 (
            .O(N__18389),
            .I(\tok.n8_adj_846 ));
    InMux I__3596 (
            .O(N__18386),
            .I(N__18380));
    InMux I__3595 (
            .O(N__18385),
            .I(N__18380));
    LocalMux I__3594 (
            .O(N__18380),
            .I(N__18377));
    Span4Mux_h I__3593 (
            .O(N__18377),
            .I(N__18374));
    Span4Mux_v I__3592 (
            .O(N__18374),
            .I(N__18371));
    Odrv4 I__3591 (
            .O(N__18371),
            .I(\tok.n41 ));
    InMux I__3590 (
            .O(N__18368),
            .I(N__18362));
    InMux I__3589 (
            .O(N__18367),
            .I(N__18362));
    LocalMux I__3588 (
            .O(N__18362),
            .I(N__18347));
    InMux I__3587 (
            .O(N__18361),
            .I(N__18342));
    InMux I__3586 (
            .O(N__18360),
            .I(N__18342));
    CascadeMux I__3585 (
            .O(N__18359),
            .I(N__18336));
    InMux I__3584 (
            .O(N__18358),
            .I(N__18331));
    InMux I__3583 (
            .O(N__18357),
            .I(N__18322));
    InMux I__3582 (
            .O(N__18356),
            .I(N__18322));
    InMux I__3581 (
            .O(N__18355),
            .I(N__18322));
    InMux I__3580 (
            .O(N__18354),
            .I(N__18322));
    CascadeMux I__3579 (
            .O(N__18353),
            .I(N__18319));
    InMux I__3578 (
            .O(N__18352),
            .I(N__18308));
    InMux I__3577 (
            .O(N__18351),
            .I(N__18308));
    InMux I__3576 (
            .O(N__18350),
            .I(N__18301));
    Span4Mux_v I__3575 (
            .O(N__18347),
            .I(N__18296));
    LocalMux I__3574 (
            .O(N__18342),
            .I(N__18296));
    InMux I__3573 (
            .O(N__18341),
            .I(N__18284));
    InMux I__3572 (
            .O(N__18340),
            .I(N__18284));
    InMux I__3571 (
            .O(N__18339),
            .I(N__18284));
    InMux I__3570 (
            .O(N__18336),
            .I(N__18284));
    InMux I__3569 (
            .O(N__18335),
            .I(N__18276));
    InMux I__3568 (
            .O(N__18334),
            .I(N__18273));
    LocalMux I__3567 (
            .O(N__18331),
            .I(N__18268));
    LocalMux I__3566 (
            .O(N__18322),
            .I(N__18268));
    InMux I__3565 (
            .O(N__18319),
            .I(N__18263));
    InMux I__3564 (
            .O(N__18318),
            .I(N__18263));
    CascadeMux I__3563 (
            .O(N__18317),
            .I(N__18259));
    CascadeMux I__3562 (
            .O(N__18316),
            .I(N__18255));
    CascadeMux I__3561 (
            .O(N__18315),
            .I(N__18252));
    CascadeMux I__3560 (
            .O(N__18314),
            .I(N__18247));
    InMux I__3559 (
            .O(N__18313),
            .I(N__18244));
    LocalMux I__3558 (
            .O(N__18308),
            .I(N__18241));
    InMux I__3557 (
            .O(N__18307),
            .I(N__18232));
    InMux I__3556 (
            .O(N__18306),
            .I(N__18232));
    InMux I__3555 (
            .O(N__18305),
            .I(N__18232));
    InMux I__3554 (
            .O(N__18304),
            .I(N__18232));
    LocalMux I__3553 (
            .O(N__18301),
            .I(N__18229));
    Span4Mux_h I__3552 (
            .O(N__18296),
            .I(N__18226));
    InMux I__3551 (
            .O(N__18295),
            .I(N__18223));
    InMux I__3550 (
            .O(N__18294),
            .I(N__18218));
    InMux I__3549 (
            .O(N__18293),
            .I(N__18218));
    LocalMux I__3548 (
            .O(N__18284),
            .I(N__18215));
    CascadeMux I__3547 (
            .O(N__18283),
            .I(N__18210));
    CascadeMux I__3546 (
            .O(N__18282),
            .I(N__18205));
    CascadeMux I__3545 (
            .O(N__18281),
            .I(N__18202));
    CascadeMux I__3544 (
            .O(N__18280),
            .I(N__18198));
    CascadeMux I__3543 (
            .O(N__18279),
            .I(N__18195));
    LocalMux I__3542 (
            .O(N__18276),
            .I(N__18189));
    LocalMux I__3541 (
            .O(N__18273),
            .I(N__18182));
    Span4Mux_v I__3540 (
            .O(N__18268),
            .I(N__18182));
    LocalMux I__3539 (
            .O(N__18263),
            .I(N__18182));
    InMux I__3538 (
            .O(N__18262),
            .I(N__18179));
    InMux I__3537 (
            .O(N__18259),
            .I(N__18164));
    InMux I__3536 (
            .O(N__18258),
            .I(N__18164));
    InMux I__3535 (
            .O(N__18255),
            .I(N__18164));
    InMux I__3534 (
            .O(N__18252),
            .I(N__18164));
    InMux I__3533 (
            .O(N__18251),
            .I(N__18164));
    InMux I__3532 (
            .O(N__18250),
            .I(N__18164));
    InMux I__3531 (
            .O(N__18247),
            .I(N__18164));
    LocalMux I__3530 (
            .O(N__18244),
            .I(N__18157));
    Span4Mux_h I__3529 (
            .O(N__18241),
            .I(N__18157));
    LocalMux I__3528 (
            .O(N__18232),
            .I(N__18157));
    Span12Mux_s10_h I__3527 (
            .O(N__18229),
            .I(N__18154));
    Span4Mux_v I__3526 (
            .O(N__18226),
            .I(N__18151));
    LocalMux I__3525 (
            .O(N__18223),
            .I(N__18144));
    LocalMux I__3524 (
            .O(N__18218),
            .I(N__18144));
    Span4Mux_v I__3523 (
            .O(N__18215),
            .I(N__18144));
    InMux I__3522 (
            .O(N__18214),
            .I(N__18141));
    InMux I__3521 (
            .O(N__18213),
            .I(N__18128));
    InMux I__3520 (
            .O(N__18210),
            .I(N__18128));
    InMux I__3519 (
            .O(N__18209),
            .I(N__18128));
    InMux I__3518 (
            .O(N__18208),
            .I(N__18128));
    InMux I__3517 (
            .O(N__18205),
            .I(N__18128));
    InMux I__3516 (
            .O(N__18202),
            .I(N__18128));
    InMux I__3515 (
            .O(N__18201),
            .I(N__18115));
    InMux I__3514 (
            .O(N__18198),
            .I(N__18115));
    InMux I__3513 (
            .O(N__18195),
            .I(N__18115));
    InMux I__3512 (
            .O(N__18194),
            .I(N__18115));
    InMux I__3511 (
            .O(N__18193),
            .I(N__18115));
    InMux I__3510 (
            .O(N__18192),
            .I(N__18115));
    Span4Mux_v I__3509 (
            .O(N__18189),
            .I(N__18110));
    Span4Mux_s2_v I__3508 (
            .O(N__18182),
            .I(N__18110));
    LocalMux I__3507 (
            .O(N__18179),
            .I(N__18103));
    LocalMux I__3506 (
            .O(N__18164),
            .I(N__18103));
    Span4Mux_v I__3505 (
            .O(N__18157),
            .I(N__18103));
    Odrv12 I__3504 (
            .O(N__18154),
            .I(\tok.T_1 ));
    Odrv4 I__3503 (
            .O(N__18151),
            .I(\tok.T_1 ));
    Odrv4 I__3502 (
            .O(N__18144),
            .I(\tok.T_1 ));
    LocalMux I__3501 (
            .O(N__18141),
            .I(\tok.T_1 ));
    LocalMux I__3500 (
            .O(N__18128),
            .I(\tok.T_1 ));
    LocalMux I__3499 (
            .O(N__18115),
            .I(\tok.T_1 ));
    Odrv4 I__3498 (
            .O(N__18110),
            .I(\tok.T_1 ));
    Odrv4 I__3497 (
            .O(N__18103),
            .I(\tok.T_1 ));
    InMux I__3496 (
            .O(N__18086),
            .I(\tok.n4761 ));
    InMux I__3495 (
            .O(N__18083),
            .I(N__18080));
    LocalMux I__3494 (
            .O(N__18080),
            .I(\tok.n15_adj_664 ));
    InMux I__3493 (
            .O(N__18077),
            .I(\tok.n4762 ));
    InMux I__3492 (
            .O(N__18074),
            .I(N__18069));
    InMux I__3491 (
            .O(N__18073),
            .I(N__18064));
    InMux I__3490 (
            .O(N__18072),
            .I(N__18064));
    LocalMux I__3489 (
            .O(N__18069),
            .I(\tok.n82 ));
    LocalMux I__3488 (
            .O(N__18064),
            .I(\tok.n82 ));
    InMux I__3487 (
            .O(N__18059),
            .I(N__18055));
    CascadeMux I__3486 (
            .O(N__18058),
            .I(N__18048));
    LocalMux I__3485 (
            .O(N__18055),
            .I(N__18043));
    InMux I__3484 (
            .O(N__18054),
            .I(N__18038));
    InMux I__3483 (
            .O(N__18053),
            .I(N__18038));
    InMux I__3482 (
            .O(N__18052),
            .I(N__18035));
    InMux I__3481 (
            .O(N__18051),
            .I(N__18031));
    InMux I__3480 (
            .O(N__18048),
            .I(N__18028));
    InMux I__3479 (
            .O(N__18047),
            .I(N__18013));
    InMux I__3478 (
            .O(N__18046),
            .I(N__18010));
    Span4Mux_s3_v I__3477 (
            .O(N__18043),
            .I(N__18003));
    LocalMux I__3476 (
            .O(N__18038),
            .I(N__18003));
    LocalMux I__3475 (
            .O(N__18035),
            .I(N__18003));
    InMux I__3474 (
            .O(N__18034),
            .I(N__17999));
    LocalMux I__3473 (
            .O(N__18031),
            .I(N__17991));
    LocalMux I__3472 (
            .O(N__18028),
            .I(N__17991));
    InMux I__3471 (
            .O(N__18027),
            .I(N__17986));
    InMux I__3470 (
            .O(N__18026),
            .I(N__17986));
    InMux I__3469 (
            .O(N__18025),
            .I(N__17983));
    CascadeMux I__3468 (
            .O(N__18024),
            .I(N__17979));
    CascadeMux I__3467 (
            .O(N__18023),
            .I(N__17976));
    CascadeMux I__3466 (
            .O(N__18022),
            .I(N__17971));
    InMux I__3465 (
            .O(N__18021),
            .I(N__17968));
    InMux I__3464 (
            .O(N__18020),
            .I(N__17951));
    InMux I__3463 (
            .O(N__18019),
            .I(N__17951));
    InMux I__3462 (
            .O(N__18018),
            .I(N__17951));
    InMux I__3461 (
            .O(N__18017),
            .I(N__17951));
    InMux I__3460 (
            .O(N__18016),
            .I(N__17951));
    LocalMux I__3459 (
            .O(N__18013),
            .I(N__17944));
    LocalMux I__3458 (
            .O(N__18010),
            .I(N__17944));
    Span4Mux_h I__3457 (
            .O(N__18003),
            .I(N__17944));
    InMux I__3456 (
            .O(N__18002),
            .I(N__17941));
    LocalMux I__3455 (
            .O(N__17999),
            .I(N__17938));
    CascadeMux I__3454 (
            .O(N__17998),
            .I(N__17935));
    CascadeMux I__3453 (
            .O(N__17997),
            .I(N__17930));
    CascadeMux I__3452 (
            .O(N__17996),
            .I(N__17927));
    Span4Mux_v I__3451 (
            .O(N__17991),
            .I(N__17921));
    LocalMux I__3450 (
            .O(N__17986),
            .I(N__17921));
    LocalMux I__3449 (
            .O(N__17983),
            .I(N__17918));
    InMux I__3448 (
            .O(N__17982),
            .I(N__17905));
    InMux I__3447 (
            .O(N__17979),
            .I(N__17905));
    InMux I__3446 (
            .O(N__17976),
            .I(N__17905));
    InMux I__3445 (
            .O(N__17975),
            .I(N__17905));
    InMux I__3444 (
            .O(N__17974),
            .I(N__17905));
    InMux I__3443 (
            .O(N__17971),
            .I(N__17905));
    LocalMux I__3442 (
            .O(N__17968),
            .I(N__17902));
    InMux I__3441 (
            .O(N__17967),
            .I(N__17889));
    InMux I__3440 (
            .O(N__17966),
            .I(N__17889));
    InMux I__3439 (
            .O(N__17965),
            .I(N__17889));
    InMux I__3438 (
            .O(N__17964),
            .I(N__17889));
    InMux I__3437 (
            .O(N__17963),
            .I(N__17889));
    InMux I__3436 (
            .O(N__17962),
            .I(N__17889));
    LocalMux I__3435 (
            .O(N__17951),
            .I(N__17886));
    Span4Mux_v I__3434 (
            .O(N__17944),
            .I(N__17881));
    LocalMux I__3433 (
            .O(N__17941),
            .I(N__17881));
    Span12Mux_s10_h I__3432 (
            .O(N__17938),
            .I(N__17878));
    InMux I__3431 (
            .O(N__17935),
            .I(N__17869));
    InMux I__3430 (
            .O(N__17934),
            .I(N__17869));
    InMux I__3429 (
            .O(N__17933),
            .I(N__17869));
    InMux I__3428 (
            .O(N__17930),
            .I(N__17869));
    InMux I__3427 (
            .O(N__17927),
            .I(N__17864));
    InMux I__3426 (
            .O(N__17926),
            .I(N__17864));
    Span4Mux_v I__3425 (
            .O(N__17921),
            .I(N__17857));
    Span4Mux_h I__3424 (
            .O(N__17918),
            .I(N__17857));
    LocalMux I__3423 (
            .O(N__17905),
            .I(N__17857));
    Span4Mux_h I__3422 (
            .O(N__17902),
            .I(N__17848));
    LocalMux I__3421 (
            .O(N__17889),
            .I(N__17848));
    Span4Mux_v I__3420 (
            .O(N__17886),
            .I(N__17848));
    Span4Mux_v I__3419 (
            .O(N__17881),
            .I(N__17848));
    Odrv12 I__3418 (
            .O(N__17878),
            .I(\tok.T_3 ));
    LocalMux I__3417 (
            .O(N__17869),
            .I(\tok.T_3 ));
    LocalMux I__3416 (
            .O(N__17864),
            .I(\tok.T_3 ));
    Odrv4 I__3415 (
            .O(N__17857),
            .I(\tok.T_3 ));
    Odrv4 I__3414 (
            .O(N__17848),
            .I(\tok.T_3 ));
    InMux I__3413 (
            .O(N__17837),
            .I(N__17834));
    LocalMux I__3412 (
            .O(N__17834),
            .I(N__17831));
    Odrv4 I__3411 (
            .O(N__17831),
            .I(\tok.n11_adj_830 ));
    InMux I__3410 (
            .O(N__17828),
            .I(\tok.n4763 ));
    InMux I__3409 (
            .O(N__17825),
            .I(N__17822));
    LocalMux I__3408 (
            .O(N__17822),
            .I(N__17819));
    Odrv12 I__3407 (
            .O(N__17819),
            .I(\tok.n212 ));
    InMux I__3406 (
            .O(N__17816),
            .I(\tok.n4764 ));
    InMux I__3405 (
            .O(N__17813),
            .I(N__17809));
    CascadeMux I__3404 (
            .O(N__17812),
            .I(N__17804));
    LocalMux I__3403 (
            .O(N__17809),
            .I(N__17801));
    InMux I__3402 (
            .O(N__17808),
            .I(N__17794));
    InMux I__3401 (
            .O(N__17807),
            .I(N__17794));
    InMux I__3400 (
            .O(N__17804),
            .I(N__17794));
    Span4Mux_v I__3399 (
            .O(N__17801),
            .I(N__17791));
    LocalMux I__3398 (
            .O(N__17794),
            .I(N__17788));
    Span4Mux_h I__3397 (
            .O(N__17791),
            .I(N__17785));
    Span4Mux_h I__3396 (
            .O(N__17788),
            .I(N__17782));
    Span4Mux_v I__3395 (
            .O(N__17785),
            .I(N__17779));
    Odrv4 I__3394 (
            .O(N__17782),
            .I(\tok.uart_tx_busy ));
    Odrv4 I__3393 (
            .O(N__17779),
            .I(\tok.uart_tx_busy ));
    CascadeMux I__3392 (
            .O(N__17774),
            .I(\tok.n15_adj_655_cascade_ ));
    InMux I__3391 (
            .O(N__17771),
            .I(N__17759));
    InMux I__3390 (
            .O(N__17770),
            .I(N__17759));
    InMux I__3389 (
            .O(N__17769),
            .I(N__17759));
    InMux I__3388 (
            .O(N__17768),
            .I(N__17759));
    LocalMux I__3387 (
            .O(N__17759),
            .I(N__17756));
    Sp12to4 I__3386 (
            .O(N__17756),
            .I(N__17753));
    Odrv12 I__3385 (
            .O(N__17753),
            .I(\tok.uart_stall ));
    CascadeMux I__3384 (
            .O(N__17750),
            .I(N__17746));
    InMux I__3383 (
            .O(N__17749),
            .I(N__17742));
    InMux I__3382 (
            .O(N__17746),
            .I(N__17737));
    InMux I__3381 (
            .O(N__17745),
            .I(N__17737));
    LocalMux I__3380 (
            .O(N__17742),
            .I(\tok.uart_rx_valid ));
    LocalMux I__3379 (
            .O(N__17737),
            .I(\tok.uart_rx_valid ));
    CEMux I__3378 (
            .O(N__17732),
            .I(N__17729));
    LocalMux I__3377 (
            .O(N__17729),
            .I(N__17726));
    Odrv4 I__3376 (
            .O(N__17726),
            .I(\tok.uart.n953 ));
    CascadeMux I__3375 (
            .O(N__17723),
            .I(\tok.n15_adj_667_cascade_ ));
    CascadeMux I__3374 (
            .O(N__17720),
            .I(N__17716));
    CascadeMux I__3373 (
            .O(N__17719),
            .I(N__17713));
    InMux I__3372 (
            .O(N__17716),
            .I(N__17710));
    InMux I__3371 (
            .O(N__17713),
            .I(N__17707));
    LocalMux I__3370 (
            .O(N__17710),
            .I(N__17704));
    LocalMux I__3369 (
            .O(N__17707),
            .I(N__17701));
    Span4Mux_h I__3368 (
            .O(N__17704),
            .I(N__17698));
    Span4Mux_s3_h I__3367 (
            .O(N__17701),
            .I(N__17695));
    Odrv4 I__3366 (
            .O(N__17698),
            .I(\tok.table_rd_2 ));
    Odrv4 I__3365 (
            .O(N__17695),
            .I(\tok.table_rd_2 ));
    CascadeMux I__3364 (
            .O(N__17690),
            .I(\tok.n28_adj_771_cascade_ ));
    InMux I__3363 (
            .O(N__17687),
            .I(N__17684));
    LocalMux I__3362 (
            .O(N__17684),
            .I(\tok.n5470 ));
    CascadeMux I__3361 (
            .O(N__17681),
            .I(\tok.n5467_cascade_ ));
    CascadeMux I__3360 (
            .O(N__17678),
            .I(N__17674));
    InMux I__3359 (
            .O(N__17677),
            .I(N__17669));
    InMux I__3358 (
            .O(N__17674),
            .I(N__17669));
    LocalMux I__3357 (
            .O(N__17669),
            .I(N__17666));
    Odrv12 I__3356 (
            .O(N__17666),
            .I(\tok.n34 ));
    CascadeMux I__3355 (
            .O(N__17663),
            .I(N__17660));
    InMux I__3354 (
            .O(N__17660),
            .I(N__17657));
    LocalMux I__3353 (
            .O(N__17657),
            .I(\tok.n5462 ));
    InMux I__3352 (
            .O(N__17654),
            .I(N__17651));
    LocalMux I__3351 (
            .O(N__17651),
            .I(\tok.n5566 ));
    InMux I__3350 (
            .O(N__17648),
            .I(N__17645));
    LocalMux I__3349 (
            .O(N__17645),
            .I(N__17642));
    Odrv4 I__3348 (
            .O(N__17642),
            .I(\tok.n5561 ));
    InMux I__3347 (
            .O(N__17639),
            .I(N__17635));
    CascadeMux I__3346 (
            .O(N__17638),
            .I(N__17632));
    LocalMux I__3345 (
            .O(N__17635),
            .I(N__17629));
    InMux I__3344 (
            .O(N__17632),
            .I(N__17626));
    Span4Mux_v I__3343 (
            .O(N__17629),
            .I(N__17621));
    LocalMux I__3342 (
            .O(N__17626),
            .I(N__17621));
    Span4Mux_v I__3341 (
            .O(N__17621),
            .I(N__17618));
    Odrv4 I__3340 (
            .O(N__17618),
            .I(\tok.n9_adj_766 ));
    InMux I__3339 (
            .O(N__17615),
            .I(N__17607));
    InMux I__3338 (
            .O(N__17614),
            .I(N__17602));
    InMux I__3337 (
            .O(N__17613),
            .I(N__17602));
    CascadeMux I__3336 (
            .O(N__17612),
            .I(N__17599));
    InMux I__3335 (
            .O(N__17611),
            .I(N__17593));
    InMux I__3334 (
            .O(N__17610),
            .I(N__17593));
    LocalMux I__3333 (
            .O(N__17607),
            .I(N__17590));
    LocalMux I__3332 (
            .O(N__17602),
            .I(N__17587));
    InMux I__3331 (
            .O(N__17599),
            .I(N__17582));
    InMux I__3330 (
            .O(N__17598),
            .I(N__17582));
    LocalMux I__3329 (
            .O(N__17593),
            .I(N__17579));
    Odrv4 I__3328 (
            .O(N__17590),
            .I(\tok.n10_adj_643 ));
    Odrv4 I__3327 (
            .O(N__17587),
            .I(\tok.n10_adj_643 ));
    LocalMux I__3326 (
            .O(N__17582),
            .I(\tok.n10_adj_643 ));
    Odrv4 I__3325 (
            .O(N__17579),
            .I(\tok.n10_adj_643 ));
    CascadeMux I__3324 (
            .O(N__17570),
            .I(N__17567));
    InMux I__3323 (
            .O(N__17567),
            .I(N__17564));
    LocalMux I__3322 (
            .O(N__17564),
            .I(N__17561));
    Span4Mux_h I__3321 (
            .O(N__17561),
            .I(N__17557));
    CascadeMux I__3320 (
            .O(N__17560),
            .I(N__17554));
    Span4Mux_h I__3319 (
            .O(N__17557),
            .I(N__17551));
    InMux I__3318 (
            .O(N__17554),
            .I(N__17548));
    Odrv4 I__3317 (
            .O(N__17551),
            .I(\tok.table_rd_0 ));
    LocalMux I__3316 (
            .O(N__17548),
            .I(\tok.table_rd_0 ));
    InMux I__3315 (
            .O(N__17543),
            .I(N__17540));
    LocalMux I__3314 (
            .O(N__17540),
            .I(N__17537));
    Odrv12 I__3313 (
            .O(N__17537),
            .I(\tok.n31 ));
    CascadeMux I__3312 (
            .O(N__17534),
            .I(\tok.n5463_cascade_ ));
    CascadeMux I__3311 (
            .O(N__17531),
            .I(N__17525));
    InMux I__3310 (
            .O(N__17530),
            .I(N__17522));
    InMux I__3309 (
            .O(N__17529),
            .I(N__17517));
    InMux I__3308 (
            .O(N__17528),
            .I(N__17517));
    InMux I__3307 (
            .O(N__17525),
            .I(N__17514));
    LocalMux I__3306 (
            .O(N__17522),
            .I(N__17509));
    LocalMux I__3305 (
            .O(N__17517),
            .I(N__17509));
    LocalMux I__3304 (
            .O(N__17514),
            .I(N__17506));
    Span4Mux_h I__3303 (
            .O(N__17509),
            .I(N__17503));
    Odrv4 I__3302 (
            .O(N__17506),
            .I(\tok.n2607 ));
    Odrv4 I__3301 (
            .O(N__17503),
            .I(\tok.n2607 ));
    InMux I__3300 (
            .O(N__17498),
            .I(N__17495));
    LocalMux I__3299 (
            .O(N__17495),
            .I(N__17492));
    Span4Mux_s2_h I__3298 (
            .O(N__17492),
            .I(N__17488));
    InMux I__3297 (
            .O(N__17491),
            .I(N__17484));
    Span4Mux_h I__3296 (
            .O(N__17488),
            .I(N__17479));
    InMux I__3295 (
            .O(N__17487),
            .I(N__17476));
    LocalMux I__3294 (
            .O(N__17484),
            .I(N__17473));
    InMux I__3293 (
            .O(N__17483),
            .I(N__17468));
    InMux I__3292 (
            .O(N__17482),
            .I(N__17468));
    Odrv4 I__3291 (
            .O(N__17479),
            .I(\tok.n14_adj_765 ));
    LocalMux I__3290 (
            .O(N__17476),
            .I(\tok.n14_adj_765 ));
    Odrv4 I__3289 (
            .O(N__17473),
            .I(\tok.n14_adj_765 ));
    LocalMux I__3288 (
            .O(N__17468),
            .I(\tok.n14_adj_765 ));
    CascadeMux I__3287 (
            .O(N__17459),
            .I(N__17455));
    InMux I__3286 (
            .O(N__17458),
            .I(N__17452));
    InMux I__3285 (
            .O(N__17455),
            .I(N__17449));
    LocalMux I__3284 (
            .O(N__17452),
            .I(N__17446));
    LocalMux I__3283 (
            .O(N__17449),
            .I(N__17443));
    Span4Mux_v I__3282 (
            .O(N__17446),
            .I(N__17440));
    Span4Mux_h I__3281 (
            .O(N__17443),
            .I(N__17437));
    Span4Mux_h I__3280 (
            .O(N__17440),
            .I(N__17434));
    Span4Mux_v I__3279 (
            .O(N__17437),
            .I(N__17431));
    Odrv4 I__3278 (
            .O(N__17434),
            .I(\tok.table_rd_1 ));
    Odrv4 I__3277 (
            .O(N__17431),
            .I(\tok.table_rd_1 ));
    CascadeMux I__3276 (
            .O(N__17426),
            .I(\tok.n5334_cascade_ ));
    CascadeMux I__3275 (
            .O(N__17423),
            .I(\tok.n14_adj_735_cascade_ ));
    CascadeMux I__3274 (
            .O(N__17420),
            .I(N__17417));
    InMux I__3273 (
            .O(N__17417),
            .I(N__17411));
    InMux I__3272 (
            .O(N__17416),
            .I(N__17411));
    LocalMux I__3271 (
            .O(N__17411),
            .I(N__17408));
    Span4Mux_h I__3270 (
            .O(N__17408),
            .I(N__17405));
    Odrv4 I__3269 (
            .O(N__17405),
            .I(\tok.n6_adj_754 ));
    CascadeMux I__3268 (
            .O(N__17402),
            .I(N__17398));
    InMux I__3267 (
            .O(N__17401),
            .I(N__17395));
    InMux I__3266 (
            .O(N__17398),
            .I(N__17392));
    LocalMux I__3265 (
            .O(N__17395),
            .I(N__17389));
    LocalMux I__3264 (
            .O(N__17392),
            .I(N__17386));
    Span4Mux_v I__3263 (
            .O(N__17389),
            .I(N__17383));
    Span4Mux_h I__3262 (
            .O(N__17386),
            .I(N__17380));
    Odrv4 I__3261 (
            .O(N__17383),
            .I(\tok.table_rd_4 ));
    Odrv4 I__3260 (
            .O(N__17380),
            .I(\tok.table_rd_4 ));
    CascadeMux I__3259 (
            .O(N__17375),
            .I(\tok.n16_adj_851_cascade_ ));
    InMux I__3258 (
            .O(N__17372),
            .I(N__17369));
    LocalMux I__3257 (
            .O(N__17369),
            .I(N__17366));
    Span4Mux_h I__3256 (
            .O(N__17366),
            .I(N__17363));
    Odrv4 I__3255 (
            .O(N__17363),
            .I(\tok.n17_adj_853 ));
    CascadeMux I__3254 (
            .O(N__17360),
            .I(\tok.n5562_cascade_ ));
    InMux I__3253 (
            .O(N__17357),
            .I(N__17354));
    LocalMux I__3252 (
            .O(N__17354),
            .I(\tok.n13_adj_852 ));
    InMux I__3251 (
            .O(N__17351),
            .I(N__17348));
    LocalMux I__3250 (
            .O(N__17348),
            .I(\tok.n14_adj_854 ));
    InMux I__3249 (
            .O(N__17345),
            .I(N__17340));
    InMux I__3248 (
            .O(N__17344),
            .I(N__17335));
    InMux I__3247 (
            .O(N__17343),
            .I(N__17335));
    LocalMux I__3246 (
            .O(N__17340),
            .I(capture_3));
    LocalMux I__3245 (
            .O(N__17335),
            .I(capture_3));
    CascadeMux I__3244 (
            .O(N__17330),
            .I(N__17327));
    InMux I__3243 (
            .O(N__17327),
            .I(N__17324));
    LocalMux I__3242 (
            .O(N__17324),
            .I(N__17321));
    Span4Mux_h I__3241 (
            .O(N__17321),
            .I(N__17317));
    InMux I__3240 (
            .O(N__17320),
            .I(N__17314));
    Sp12to4 I__3239 (
            .O(N__17317),
            .I(N__17311));
    LocalMux I__3238 (
            .O(N__17314),
            .I(capture_0));
    Odrv12 I__3237 (
            .O(N__17311),
            .I(capture_0));
    InMux I__3236 (
            .O(N__17306),
            .I(N__17297));
    InMux I__3235 (
            .O(N__17305),
            .I(N__17297));
    InMux I__3234 (
            .O(N__17304),
            .I(N__17297));
    LocalMux I__3233 (
            .O(N__17297),
            .I(capture_1));
    CascadeMux I__3232 (
            .O(N__17294),
            .I(N__17290));
    InMux I__3231 (
            .O(N__17293),
            .I(N__17285));
    InMux I__3230 (
            .O(N__17290),
            .I(N__17285));
    LocalMux I__3229 (
            .O(N__17285),
            .I(uart_rx_data_0));
    CascadeMux I__3228 (
            .O(N__17282),
            .I(\tok.n6_adj_794_cascade_ ));
    CascadeMux I__3227 (
            .O(N__17279),
            .I(N__17276));
    InMux I__3226 (
            .O(N__17276),
            .I(N__17272));
    InMux I__3225 (
            .O(N__17275),
            .I(N__17269));
    LocalMux I__3224 (
            .O(N__17272),
            .I(N__17266));
    LocalMux I__3223 (
            .O(N__17269),
            .I(N__17263));
    Span4Mux_v I__3222 (
            .O(N__17266),
            .I(N__17260));
    Span4Mux_v I__3221 (
            .O(N__17263),
            .I(N__17257));
    Span4Mux_v I__3220 (
            .O(N__17260),
            .I(N__17254));
    Odrv4 I__3219 (
            .O(N__17257),
            .I(\tok.table_rd_6 ));
    Odrv4 I__3218 (
            .O(N__17254),
            .I(\tok.table_rd_6 ));
    CascadeMux I__3217 (
            .O(N__17249),
            .I(\tok.n5553_cascade_ ));
    InMux I__3216 (
            .O(N__17246),
            .I(N__17243));
    LocalMux I__3215 (
            .O(N__17243),
            .I(N__17240));
    Span4Mux_v I__3214 (
            .O(N__17240),
            .I(N__17237));
    Odrv4 I__3213 (
            .O(N__17237),
            .I(\tok.table_rd_14 ));
    InMux I__3212 (
            .O(N__17234),
            .I(N__17231));
    LocalMux I__3211 (
            .O(N__17231),
            .I(N__17228));
    Span4Mux_v I__3210 (
            .O(N__17228),
            .I(N__17225));
    Span4Mux_h I__3209 (
            .O(N__17225),
            .I(N__17222));
    Odrv4 I__3208 (
            .O(N__17222),
            .I(\tok.table_rd_12 ));
    InMux I__3207 (
            .O(N__17219),
            .I(N__17216));
    LocalMux I__3206 (
            .O(N__17216),
            .I(N__17212));
    InMux I__3205 (
            .O(N__17215),
            .I(N__17209));
    Span4Mux_v I__3204 (
            .O(N__17212),
            .I(N__17206));
    LocalMux I__3203 (
            .O(N__17209),
            .I(tail_110));
    Odrv4 I__3202 (
            .O(N__17206),
            .I(tail_110));
    InMux I__3201 (
            .O(N__17201),
            .I(N__17198));
    LocalMux I__3200 (
            .O(N__17198),
            .I(N__17194));
    InMux I__3199 (
            .O(N__17197),
            .I(N__17191));
    Odrv12 I__3198 (
            .O(N__17194),
            .I(tail_126));
    LocalMux I__3197 (
            .O(N__17191),
            .I(tail_126));
    CascadeMux I__3196 (
            .O(N__17186),
            .I(N__17183));
    InMux I__3195 (
            .O(N__17183),
            .I(N__17180));
    LocalMux I__3194 (
            .O(N__17180),
            .I(N__17177));
    Span4Mux_v I__3193 (
            .O(N__17177),
            .I(N__17173));
    InMux I__3192 (
            .O(N__17176),
            .I(N__17170));
    Sp12to4 I__3191 (
            .O(N__17173),
            .I(N__17167));
    LocalMux I__3190 (
            .O(N__17170),
            .I(N__17164));
    Odrv12 I__3189 (
            .O(N__17167),
            .I(tail_111));
    Odrv12 I__3188 (
            .O(N__17164),
            .I(tail_111));
    InMux I__3187 (
            .O(N__17159),
            .I(N__17155));
    InMux I__3186 (
            .O(N__17158),
            .I(N__17152));
    LocalMux I__3185 (
            .O(N__17155),
            .I(N__17148));
    LocalMux I__3184 (
            .O(N__17152),
            .I(N__17145));
    InMux I__3183 (
            .O(N__17151),
            .I(N__17142));
    Span4Mux_h I__3182 (
            .O(N__17148),
            .I(N__17137));
    Span4Mux_h I__3181 (
            .O(N__17145),
            .I(N__17137));
    LocalMux I__3180 (
            .O(N__17142),
            .I(N__17134));
    Sp12to4 I__3179 (
            .O(N__17137),
            .I(N__17131));
    Span4Mux_h I__3178 (
            .O(N__17134),
            .I(N__17128));
    Odrv12 I__3177 (
            .O(N__17131),
            .I(rx_c));
    Odrv4 I__3176 (
            .O(N__17128),
            .I(rx_c));
    InMux I__3175 (
            .O(N__17123),
            .I(N__17120));
    LocalMux I__3174 (
            .O(N__17120),
            .I(N__17117));
    Span4Mux_h I__3173 (
            .O(N__17117),
            .I(N__17114));
    Odrv4 I__3172 (
            .O(N__17114),
            .I(\tok.uart.n5235 ));
    CascadeMux I__3171 (
            .O(N__17111),
            .I(N__17108));
    InMux I__3170 (
            .O(N__17108),
            .I(N__17102));
    InMux I__3169 (
            .O(N__17107),
            .I(N__17102));
    LocalMux I__3168 (
            .O(N__17102),
            .I(N__17098));
    InMux I__3167 (
            .O(N__17101),
            .I(N__17094));
    Span4Mux_h I__3166 (
            .O(N__17098),
            .I(N__17091));
    InMux I__3165 (
            .O(N__17097),
            .I(N__17088));
    LocalMux I__3164 (
            .O(N__17094),
            .I(N__17083));
    Span4Mux_h I__3163 (
            .O(N__17091),
            .I(N__17083));
    LocalMux I__3162 (
            .O(N__17088),
            .I(\tok.uart.bytephase_5 ));
    Odrv4 I__3161 (
            .O(N__17083),
            .I(\tok.uart.bytephase_5 ));
    CascadeMux I__3160 (
            .O(N__17078),
            .I(N__17073));
    InMux I__3159 (
            .O(N__17077),
            .I(N__17068));
    InMux I__3158 (
            .O(N__17076),
            .I(N__17068));
    InMux I__3157 (
            .O(N__17073),
            .I(N__17064));
    LocalMux I__3156 (
            .O(N__17068),
            .I(N__17061));
    InMux I__3155 (
            .O(N__17067),
            .I(N__17058));
    LocalMux I__3154 (
            .O(N__17064),
            .I(N__17053));
    Span12Mux_s11_h I__3153 (
            .O(N__17061),
            .I(N__17053));
    LocalMux I__3152 (
            .O(N__17058),
            .I(\tok.uart.bytephase_3 ));
    Odrv12 I__3151 (
            .O(N__17053),
            .I(\tok.uart.bytephase_3 ));
    InMux I__3150 (
            .O(N__17048),
            .I(N__17045));
    LocalMux I__3149 (
            .O(N__17045),
            .I(N__17042));
    Span4Mux_v I__3148 (
            .O(N__17042),
            .I(N__17039));
    Odrv4 I__3147 (
            .O(N__17039),
            .I(\tok.uart.n5374 ));
    InMux I__3146 (
            .O(N__17036),
            .I(N__17032));
    InMux I__3145 (
            .O(N__17035),
            .I(N__17029));
    LocalMux I__3144 (
            .O(N__17032),
            .I(N__17024));
    LocalMux I__3143 (
            .O(N__17029),
            .I(N__17024));
    Span4Mux_h I__3142 (
            .O(N__17024),
            .I(N__17021));
    Odrv4 I__3141 (
            .O(N__17021),
            .I(\tok.key_rd_13 ));
    InMux I__3140 (
            .O(N__17018),
            .I(N__17015));
    LocalMux I__3139 (
            .O(N__17015),
            .I(N__17012));
    Odrv4 I__3138 (
            .O(N__17012),
            .I(\tok.n14_adj_647 ));
    CascadeMux I__3137 (
            .O(N__17009),
            .I(\tok.n27_adj_818_cascade_ ));
    CascadeMux I__3136 (
            .O(N__17006),
            .I(N__17002));
    CascadeMux I__3135 (
            .O(N__17005),
            .I(N__16999));
    CascadeBuf I__3134 (
            .O(N__17002),
            .I(N__16996));
    CascadeBuf I__3133 (
            .O(N__16999),
            .I(N__16993));
    CascadeMux I__3132 (
            .O(N__16996),
            .I(N__16990));
    CascadeMux I__3131 (
            .O(N__16993),
            .I(N__16987));
    InMux I__3130 (
            .O(N__16990),
            .I(N__16984));
    InMux I__3129 (
            .O(N__16987),
            .I(N__16981));
    LocalMux I__3128 (
            .O(N__16984),
            .I(N__16976));
    LocalMux I__3127 (
            .O(N__16981),
            .I(N__16976));
    Span4Mux_v I__3126 (
            .O(N__16976),
            .I(N__16970));
    InMux I__3125 (
            .O(N__16975),
            .I(N__16967));
    InMux I__3124 (
            .O(N__16974),
            .I(N__16964));
    InMux I__3123 (
            .O(N__16973),
            .I(N__16961));
    Span4Mux_h I__3122 (
            .O(N__16970),
            .I(N__16958));
    LocalMux I__3121 (
            .O(N__16967),
            .I(\tok.idx_2 ));
    LocalMux I__3120 (
            .O(N__16964),
            .I(\tok.idx_2 ));
    LocalMux I__3119 (
            .O(N__16961),
            .I(\tok.idx_2 ));
    Odrv4 I__3118 (
            .O(N__16958),
            .I(\tok.idx_2 ));
    InMux I__3117 (
            .O(N__16949),
            .I(N__16945));
    CascadeMux I__3116 (
            .O(N__16948),
            .I(N__16936));
    LocalMux I__3115 (
            .O(N__16945),
            .I(N__16927));
    InMux I__3114 (
            .O(N__16944),
            .I(N__16924));
    InMux I__3113 (
            .O(N__16943),
            .I(N__16917));
    InMux I__3112 (
            .O(N__16942),
            .I(N__16917));
    InMux I__3111 (
            .O(N__16941),
            .I(N__16912));
    InMux I__3110 (
            .O(N__16940),
            .I(N__16912));
    InMux I__3109 (
            .O(N__16939),
            .I(N__16909));
    InMux I__3108 (
            .O(N__16936),
            .I(N__16902));
    InMux I__3107 (
            .O(N__16935),
            .I(N__16902));
    InMux I__3106 (
            .O(N__16934),
            .I(N__16902));
    InMux I__3105 (
            .O(N__16933),
            .I(N__16893));
    InMux I__3104 (
            .O(N__16932),
            .I(N__16893));
    InMux I__3103 (
            .O(N__16931),
            .I(N__16893));
    InMux I__3102 (
            .O(N__16930),
            .I(N__16893));
    Span4Mux_v I__3101 (
            .O(N__16927),
            .I(N__16890));
    LocalMux I__3100 (
            .O(N__16924),
            .I(N__16887));
    InMux I__3099 (
            .O(N__16923),
            .I(N__16882));
    InMux I__3098 (
            .O(N__16922),
            .I(N__16882));
    LocalMux I__3097 (
            .O(N__16917),
            .I(\tok.stall ));
    LocalMux I__3096 (
            .O(N__16912),
            .I(\tok.stall ));
    LocalMux I__3095 (
            .O(N__16909),
            .I(\tok.stall ));
    LocalMux I__3094 (
            .O(N__16902),
            .I(\tok.stall ));
    LocalMux I__3093 (
            .O(N__16893),
            .I(\tok.stall ));
    Odrv4 I__3092 (
            .O(N__16890),
            .I(\tok.stall ));
    Odrv12 I__3091 (
            .O(N__16887),
            .I(\tok.stall ));
    LocalMux I__3090 (
            .O(N__16882),
            .I(\tok.stall ));
    InMux I__3089 (
            .O(N__16865),
            .I(N__16862));
    LocalMux I__3088 (
            .O(N__16862),
            .I(\tok.n33_adj_821 ));
    CascadeMux I__3087 (
            .O(N__16859),
            .I(N__16850));
    CascadeMux I__3086 (
            .O(N__16858),
            .I(N__16845));
    CascadeMux I__3085 (
            .O(N__16857),
            .I(N__16841));
    CascadeMux I__3084 (
            .O(N__16856),
            .I(N__16838));
    InMux I__3083 (
            .O(N__16855),
            .I(N__16828));
    InMux I__3082 (
            .O(N__16854),
            .I(N__16828));
    InMux I__3081 (
            .O(N__16853),
            .I(N__16828));
    InMux I__3080 (
            .O(N__16850),
            .I(N__16828));
    InMux I__3079 (
            .O(N__16849),
            .I(N__16821));
    InMux I__3078 (
            .O(N__16848),
            .I(N__16821));
    InMux I__3077 (
            .O(N__16845),
            .I(N__16821));
    InMux I__3076 (
            .O(N__16844),
            .I(N__16812));
    InMux I__3075 (
            .O(N__16841),
            .I(N__16812));
    InMux I__3074 (
            .O(N__16838),
            .I(N__16812));
    InMux I__3073 (
            .O(N__16837),
            .I(N__16812));
    LocalMux I__3072 (
            .O(N__16828),
            .I(\tok.search_clk ));
    LocalMux I__3071 (
            .O(N__16821),
            .I(\tok.search_clk ));
    LocalMux I__3070 (
            .O(N__16812),
            .I(\tok.search_clk ));
    CascadeMux I__3069 (
            .O(N__16805),
            .I(\tok.n27_adj_822_cascade_ ));
    CascadeMux I__3068 (
            .O(N__16802),
            .I(N__16799));
    CascadeBuf I__3067 (
            .O(N__16799),
            .I(N__16795));
    CascadeMux I__3066 (
            .O(N__16798),
            .I(N__16792));
    CascadeMux I__3065 (
            .O(N__16795),
            .I(N__16789));
    CascadeBuf I__3064 (
            .O(N__16792),
            .I(N__16786));
    InMux I__3063 (
            .O(N__16789),
            .I(N__16783));
    CascadeMux I__3062 (
            .O(N__16786),
            .I(N__16780));
    LocalMux I__3061 (
            .O(N__16783),
            .I(N__16777));
    InMux I__3060 (
            .O(N__16780),
            .I(N__16774));
    Span4Mux_h I__3059 (
            .O(N__16777),
            .I(N__16771));
    LocalMux I__3058 (
            .O(N__16774),
            .I(N__16765));
    Span4Mux_h I__3057 (
            .O(N__16771),
            .I(N__16762));
    InMux I__3056 (
            .O(N__16770),
            .I(N__16759));
    InMux I__3055 (
            .O(N__16769),
            .I(N__16756));
    InMux I__3054 (
            .O(N__16768),
            .I(N__16753));
    Span12Mux_s7_h I__3053 (
            .O(N__16765),
            .I(N__16750));
    Span4Mux_v I__3052 (
            .O(N__16762),
            .I(N__16747));
    LocalMux I__3051 (
            .O(N__16759),
            .I(\tok.idx_3 ));
    LocalMux I__3050 (
            .O(N__16756),
            .I(\tok.idx_3 ));
    LocalMux I__3049 (
            .O(N__16753),
            .I(\tok.idx_3 ));
    Odrv12 I__3048 (
            .O(N__16750),
            .I(\tok.idx_3 ));
    Odrv4 I__3047 (
            .O(N__16747),
            .I(\tok.idx_3 ));
    InMux I__3046 (
            .O(N__16736),
            .I(N__16720));
    InMux I__3045 (
            .O(N__16735),
            .I(N__16720));
    InMux I__3044 (
            .O(N__16734),
            .I(N__16720));
    InMux I__3043 (
            .O(N__16733),
            .I(N__16720));
    InMux I__3042 (
            .O(N__16732),
            .I(N__16713));
    InMux I__3041 (
            .O(N__16731),
            .I(N__16713));
    InMux I__3040 (
            .O(N__16730),
            .I(N__16713));
    InMux I__3039 (
            .O(N__16729),
            .I(N__16710));
    LocalMux I__3038 (
            .O(N__16720),
            .I(\tok.n2699 ));
    LocalMux I__3037 (
            .O(N__16713),
            .I(\tok.n2699 ));
    LocalMux I__3036 (
            .O(N__16710),
            .I(\tok.n2699 ));
    CascadeMux I__3035 (
            .O(N__16703),
            .I(N__16694));
    InMux I__3034 (
            .O(N__16702),
            .I(N__16684));
    InMux I__3033 (
            .O(N__16701),
            .I(N__16684));
    InMux I__3032 (
            .O(N__16700),
            .I(N__16684));
    InMux I__3031 (
            .O(N__16699),
            .I(N__16684));
    InMux I__3030 (
            .O(N__16698),
            .I(N__16677));
    InMux I__3029 (
            .O(N__16697),
            .I(N__16677));
    InMux I__3028 (
            .O(N__16694),
            .I(N__16677));
    InMux I__3027 (
            .O(N__16693),
            .I(N__16674));
    LocalMux I__3026 (
            .O(N__16684),
            .I(\tok.n5282 ));
    LocalMux I__3025 (
            .O(N__16677),
            .I(\tok.n5282 ));
    LocalMux I__3024 (
            .O(N__16674),
            .I(\tok.n5282 ));
    InMux I__3023 (
            .O(N__16667),
            .I(N__16664));
    LocalMux I__3022 (
            .O(N__16664),
            .I(\tok.n27_adj_815 ));
    CascadeMux I__3021 (
            .O(N__16661),
            .I(N__16658));
    CascadeBuf I__3020 (
            .O(N__16658),
            .I(N__16654));
    CascadeMux I__3019 (
            .O(N__16657),
            .I(N__16651));
    CascadeMux I__3018 (
            .O(N__16654),
            .I(N__16648));
    CascadeBuf I__3017 (
            .O(N__16651),
            .I(N__16645));
    InMux I__3016 (
            .O(N__16648),
            .I(N__16642));
    CascadeMux I__3015 (
            .O(N__16645),
            .I(N__16639));
    LocalMux I__3014 (
            .O(N__16642),
            .I(N__16636));
    InMux I__3013 (
            .O(N__16639),
            .I(N__16633));
    Span4Mux_h I__3012 (
            .O(N__16636),
            .I(N__16627));
    LocalMux I__3011 (
            .O(N__16633),
            .I(N__16624));
    InMux I__3010 (
            .O(N__16632),
            .I(N__16621));
    InMux I__3009 (
            .O(N__16631),
            .I(N__16618));
    InMux I__3008 (
            .O(N__16630),
            .I(N__16615));
    Sp12to4 I__3007 (
            .O(N__16627),
            .I(N__16610));
    Span12Mux_s7_h I__3006 (
            .O(N__16624),
            .I(N__16610));
    LocalMux I__3005 (
            .O(N__16621),
            .I(\tok.idx_1 ));
    LocalMux I__3004 (
            .O(N__16618),
            .I(\tok.idx_1 ));
    LocalMux I__3003 (
            .O(N__16615),
            .I(\tok.idx_1 ));
    Odrv12 I__3002 (
            .O(N__16610),
            .I(\tok.idx_1 ));
    CascadeMux I__3001 (
            .O(N__16601),
            .I(rd_15__N_301_cascade_));
    CascadeMux I__3000 (
            .O(N__16598),
            .I(N__16595));
    InMux I__2999 (
            .O(N__16595),
            .I(N__16589));
    InMux I__2998 (
            .O(N__16594),
            .I(N__16589));
    LocalMux I__2997 (
            .O(N__16589),
            .I(\tok.n797 ));
    InMux I__2996 (
            .O(N__16586),
            .I(N__16579));
    InMux I__2995 (
            .O(N__16585),
            .I(N__16579));
    InMux I__2994 (
            .O(N__16584),
            .I(N__16576));
    LocalMux I__2993 (
            .O(N__16579),
            .I(N__16573));
    LocalMux I__2992 (
            .O(N__16576),
            .I(N__16570));
    Odrv4 I__2991 (
            .O(N__16573),
            .I(\tok.n2585 ));
    Odrv4 I__2990 (
            .O(N__16570),
            .I(\tok.n2585 ));
    CascadeMux I__2989 (
            .O(N__16565),
            .I(A_stk_delta_1_cascade_));
    InMux I__2988 (
            .O(N__16562),
            .I(N__16556));
    InMux I__2987 (
            .O(N__16561),
            .I(N__16556));
    LocalMux I__2986 (
            .O(N__16556),
            .I(\tok.A_stk.tail_78 ));
    InMux I__2985 (
            .O(N__16553),
            .I(N__16547));
    InMux I__2984 (
            .O(N__16552),
            .I(N__16547));
    LocalMux I__2983 (
            .O(N__16547),
            .I(\tok.A_stk.tail_62 ));
    InMux I__2982 (
            .O(N__16544),
            .I(N__16538));
    InMux I__2981 (
            .O(N__16543),
            .I(N__16538));
    LocalMux I__2980 (
            .O(N__16538),
            .I(\tok.A_stk.tail_46 ));
    InMux I__2979 (
            .O(N__16535),
            .I(N__16529));
    InMux I__2978 (
            .O(N__16534),
            .I(N__16529));
    LocalMux I__2977 (
            .O(N__16529),
            .I(\tok.A_stk.tail_30 ));
    InMux I__2976 (
            .O(N__16526),
            .I(N__16523));
    LocalMux I__2975 (
            .O(N__16523),
            .I(N__16520));
    Span4Mux_s2_v I__2974 (
            .O(N__16520),
            .I(N__16517));
    Span4Mux_h I__2973 (
            .O(N__16517),
            .I(N__16513));
    InMux I__2972 (
            .O(N__16516),
            .I(N__16510));
    Odrv4 I__2971 (
            .O(N__16513),
            .I(tail_127));
    LocalMux I__2970 (
            .O(N__16510),
            .I(tail_127));
    InMux I__2969 (
            .O(N__16505),
            .I(N__16502));
    LocalMux I__2968 (
            .O(N__16502),
            .I(\tok.n33_adj_814 ));
    CascadeMux I__2967 (
            .O(N__16499),
            .I(N__16494));
    InMux I__2966 (
            .O(N__16498),
            .I(N__16489));
    CascadeMux I__2965 (
            .O(N__16497),
            .I(N__16485));
    InMux I__2964 (
            .O(N__16494),
            .I(N__16481));
    CascadeMux I__2963 (
            .O(N__16493),
            .I(N__16477));
    CascadeMux I__2962 (
            .O(N__16492),
            .I(N__16473));
    LocalMux I__2961 (
            .O(N__16489),
            .I(N__16470));
    InMux I__2960 (
            .O(N__16488),
            .I(N__16463));
    InMux I__2959 (
            .O(N__16485),
            .I(N__16463));
    InMux I__2958 (
            .O(N__16484),
            .I(N__16463));
    LocalMux I__2957 (
            .O(N__16481),
            .I(N__16460));
    InMux I__2956 (
            .O(N__16480),
            .I(N__16451));
    InMux I__2955 (
            .O(N__16477),
            .I(N__16451));
    InMux I__2954 (
            .O(N__16476),
            .I(N__16451));
    InMux I__2953 (
            .O(N__16473),
            .I(N__16451));
    Odrv4 I__2952 (
            .O(N__16470),
            .I(\tok.n62 ));
    LocalMux I__2951 (
            .O(N__16463),
            .I(\tok.n62 ));
    Odrv4 I__2950 (
            .O(N__16460),
            .I(\tok.n62 ));
    LocalMux I__2949 (
            .O(N__16451),
            .I(\tok.n62 ));
    InMux I__2948 (
            .O(N__16442),
            .I(N__16439));
    LocalMux I__2947 (
            .O(N__16439),
            .I(N__16436));
    Span4Mux_h I__2946 (
            .O(N__16436),
            .I(N__16429));
    InMux I__2945 (
            .O(N__16435),
            .I(N__16422));
    InMux I__2944 (
            .O(N__16434),
            .I(N__16422));
    InMux I__2943 (
            .O(N__16433),
            .I(N__16422));
    InMux I__2942 (
            .O(N__16432),
            .I(N__16419));
    Odrv4 I__2941 (
            .O(N__16429),
            .I(\tok.n1_adj_715 ));
    LocalMux I__2940 (
            .O(N__16422),
            .I(\tok.n1_adj_715 ));
    LocalMux I__2939 (
            .O(N__16419),
            .I(\tok.n1_adj_715 ));
    CascadeMux I__2938 (
            .O(N__16412),
            .I(\tok.depth_0_cascade_ ));
    InMux I__2937 (
            .O(N__16409),
            .I(N__16406));
    LocalMux I__2936 (
            .O(N__16406),
            .I(N__16403));
    Odrv12 I__2935 (
            .O(N__16403),
            .I(\tok.n5408 ));
    InMux I__2934 (
            .O(N__16400),
            .I(N__16397));
    LocalMux I__2933 (
            .O(N__16397),
            .I(\tok.n33_adj_816 ));
    InMux I__2932 (
            .O(N__16394),
            .I(N__16391));
    LocalMux I__2931 (
            .O(N__16391),
            .I(N__16387));
    InMux I__2930 (
            .O(N__16390),
            .I(N__16384));
    Span4Mux_h I__2929 (
            .O(N__16387),
            .I(N__16377));
    LocalMux I__2928 (
            .O(N__16384),
            .I(N__16377));
    CascadeMux I__2927 (
            .O(N__16383),
            .I(N__16374));
    CascadeMux I__2926 (
            .O(N__16382),
            .I(N__16371));
    Span4Mux_v I__2925 (
            .O(N__16377),
            .I(N__16366));
    InMux I__2924 (
            .O(N__16374),
            .I(N__16361));
    InMux I__2923 (
            .O(N__16371),
            .I(N__16361));
    InMux I__2922 (
            .O(N__16370),
            .I(N__16358));
    InMux I__2921 (
            .O(N__16369),
            .I(N__16354));
    Span4Mux_s3_h I__2920 (
            .O(N__16366),
            .I(N__16348));
    LocalMux I__2919 (
            .O(N__16361),
            .I(N__16348));
    LocalMux I__2918 (
            .O(N__16358),
            .I(N__16345));
    InMux I__2917 (
            .O(N__16357),
            .I(N__16342));
    LocalMux I__2916 (
            .O(N__16354),
            .I(N__16339));
    InMux I__2915 (
            .O(N__16353),
            .I(N__16336));
    Span4Mux_v I__2914 (
            .O(N__16348),
            .I(N__16333));
    Span4Mux_h I__2913 (
            .O(N__16345),
            .I(N__16330));
    LocalMux I__2912 (
            .O(N__16342),
            .I(N__16327));
    Odrv12 I__2911 (
            .O(N__16339),
            .I(\tok.n820 ));
    LocalMux I__2910 (
            .O(N__16336),
            .I(\tok.n820 ));
    Odrv4 I__2909 (
            .O(N__16333),
            .I(\tok.n820 ));
    Odrv4 I__2908 (
            .O(N__16330),
            .I(\tok.n820 ));
    Odrv4 I__2907 (
            .O(N__16327),
            .I(\tok.n820 ));
    InMux I__2906 (
            .O(N__16316),
            .I(N__16313));
    LocalMux I__2905 (
            .O(N__16313),
            .I(N__16306));
    InMux I__2904 (
            .O(N__16312),
            .I(N__16303));
    InMux I__2903 (
            .O(N__16311),
            .I(N__16298));
    InMux I__2902 (
            .O(N__16310),
            .I(N__16298));
    InMux I__2901 (
            .O(N__16309),
            .I(N__16295));
    Span4Mux_v I__2900 (
            .O(N__16306),
            .I(N__16290));
    LocalMux I__2899 (
            .O(N__16303),
            .I(N__16285));
    LocalMux I__2898 (
            .O(N__16298),
            .I(N__16285));
    LocalMux I__2897 (
            .O(N__16295),
            .I(N__16282));
    InMux I__2896 (
            .O(N__16294),
            .I(N__16278));
    InMux I__2895 (
            .O(N__16293),
            .I(N__16275));
    Span4Mux_v I__2894 (
            .O(N__16290),
            .I(N__16268));
    Span4Mux_v I__2893 (
            .O(N__16285),
            .I(N__16268));
    Span4Mux_v I__2892 (
            .O(N__16282),
            .I(N__16268));
    InMux I__2891 (
            .O(N__16281),
            .I(N__16265));
    LocalMux I__2890 (
            .O(N__16278),
            .I(\tok.n5298 ));
    LocalMux I__2889 (
            .O(N__16275),
            .I(\tok.n5298 ));
    Odrv4 I__2888 (
            .O(N__16268),
            .I(\tok.n5298 ));
    LocalMux I__2887 (
            .O(N__16265),
            .I(\tok.n5298 ));
    CascadeMux I__2886 (
            .O(N__16256),
            .I(\tok.n13_adj_673_cascade_ ));
    InMux I__2885 (
            .O(N__16253),
            .I(N__16248));
    InMux I__2884 (
            .O(N__16252),
            .I(N__16243));
    InMux I__2883 (
            .O(N__16251),
            .I(N__16243));
    LocalMux I__2882 (
            .O(N__16248),
            .I(N__16239));
    LocalMux I__2881 (
            .O(N__16243),
            .I(N__16236));
    InMux I__2880 (
            .O(N__16242),
            .I(N__16233));
    Span4Mux_h I__2879 (
            .O(N__16239),
            .I(N__16228));
    Span4Mux_s3_v I__2878 (
            .O(N__16236),
            .I(N__16228));
    LocalMux I__2877 (
            .O(N__16233),
            .I(\tok.tc_plus_1_4 ));
    Odrv4 I__2876 (
            .O(N__16228),
            .I(\tok.tc_plus_1_4 ));
    CascadeMux I__2875 (
            .O(N__16223),
            .I(n10_adj_870_cascade_));
    CascadeMux I__2874 (
            .O(N__16220),
            .I(N__16217));
    InMux I__2873 (
            .O(N__16217),
            .I(N__16214));
    LocalMux I__2872 (
            .O(N__16214),
            .I(N__16211));
    Span4Mux_h I__2871 (
            .O(N__16211),
            .I(N__16208));
    Odrv4 I__2870 (
            .O(N__16208),
            .I(\tok.tc_4 ));
    CascadeMux I__2869 (
            .O(N__16205),
            .I(N__16198));
    InMux I__2868 (
            .O(N__16204),
            .I(N__16191));
    InMux I__2867 (
            .O(N__16203),
            .I(N__16186));
    InMux I__2866 (
            .O(N__16202),
            .I(N__16186));
    InMux I__2865 (
            .O(N__16201),
            .I(N__16173));
    InMux I__2864 (
            .O(N__16198),
            .I(N__16173));
    InMux I__2863 (
            .O(N__16197),
            .I(N__16173));
    InMux I__2862 (
            .O(N__16196),
            .I(N__16173));
    InMux I__2861 (
            .O(N__16195),
            .I(N__16173));
    InMux I__2860 (
            .O(N__16194),
            .I(N__16173));
    LocalMux I__2859 (
            .O(N__16191),
            .I(N__16168));
    LocalMux I__2858 (
            .O(N__16186),
            .I(N__16165));
    LocalMux I__2857 (
            .O(N__16173),
            .I(N__16159));
    InMux I__2856 (
            .O(N__16172),
            .I(N__16154));
    InMux I__2855 (
            .O(N__16171),
            .I(N__16154));
    Span4Mux_v I__2854 (
            .O(N__16168),
            .I(N__16149));
    Span4Mux_h I__2853 (
            .O(N__16165),
            .I(N__16149));
    InMux I__2852 (
            .O(N__16164),
            .I(N__16144));
    InMux I__2851 (
            .O(N__16163),
            .I(N__16144));
    InMux I__2850 (
            .O(N__16162),
            .I(N__16141));
    Span4Mux_h I__2849 (
            .O(N__16159),
            .I(N__16136));
    LocalMux I__2848 (
            .O(N__16154),
            .I(N__16136));
    Sp12to4 I__2847 (
            .O(N__16149),
            .I(N__16127));
    LocalMux I__2846 (
            .O(N__16144),
            .I(N__16127));
    LocalMux I__2845 (
            .O(N__16141),
            .I(N__16127));
    Span4Mux_v I__2844 (
            .O(N__16136),
            .I(N__16124));
    InMux I__2843 (
            .O(N__16135),
            .I(N__16119));
    InMux I__2842 (
            .O(N__16134),
            .I(N__16119));
    Odrv12 I__2841 (
            .O(N__16127),
            .I(stall_));
    Odrv4 I__2840 (
            .O(N__16124),
            .I(stall_));
    LocalMux I__2839 (
            .O(N__16119),
            .I(stall_));
    InMux I__2838 (
            .O(N__16112),
            .I(N__16109));
    LocalMux I__2837 (
            .O(N__16109),
            .I(n10_adj_870));
    InMux I__2836 (
            .O(N__16106),
            .I(N__16101));
    InMux I__2835 (
            .O(N__16105),
            .I(N__16098));
    CascadeMux I__2834 (
            .O(N__16104),
            .I(N__16095));
    LocalMux I__2833 (
            .O(N__16101),
            .I(N__16091));
    LocalMux I__2832 (
            .O(N__16098),
            .I(N__16088));
    InMux I__2831 (
            .O(N__16095),
            .I(N__16083));
    InMux I__2830 (
            .O(N__16094),
            .I(N__16083));
    Span4Mux_v I__2829 (
            .O(N__16091),
            .I(N__16080));
    Odrv12 I__2828 (
            .O(N__16088),
            .I(tc_4));
    LocalMux I__2827 (
            .O(N__16083),
            .I(tc_4));
    Odrv4 I__2826 (
            .O(N__16080),
            .I(tc_4));
    InMux I__2825 (
            .O(N__16073),
            .I(N__16068));
    CascadeMux I__2824 (
            .O(N__16072),
            .I(N__16064));
    CascadeMux I__2823 (
            .O(N__16071),
            .I(N__16061));
    LocalMux I__2822 (
            .O(N__16068),
            .I(N__16058));
    InMux I__2821 (
            .O(N__16067),
            .I(N__16053));
    InMux I__2820 (
            .O(N__16064),
            .I(N__16053));
    InMux I__2819 (
            .O(N__16061),
            .I(N__16050));
    Span4Mux_s2_v I__2818 (
            .O(N__16058),
            .I(N__16047));
    LocalMux I__2817 (
            .O(N__16053),
            .I(N__16044));
    LocalMux I__2816 (
            .O(N__16050),
            .I(\tok.c_stk_r_4 ));
    Odrv4 I__2815 (
            .O(N__16047),
            .I(\tok.c_stk_r_4 ));
    Odrv12 I__2814 (
            .O(N__16044),
            .I(\tok.c_stk_r_4 ));
    CascadeMux I__2813 (
            .O(N__16037),
            .I(\tok.n83_adj_665_cascade_ ));
    CascadeMux I__2812 (
            .O(N__16034),
            .I(N__16031));
    InMux I__2811 (
            .O(N__16031),
            .I(N__16028));
    LocalMux I__2810 (
            .O(N__16028),
            .I(\tok.n5487 ));
    InMux I__2809 (
            .O(N__16025),
            .I(N__16021));
    InMux I__2808 (
            .O(N__16024),
            .I(N__16018));
    LocalMux I__2807 (
            .O(N__16021),
            .I(\tok.A_stk.tail_94 ));
    LocalMux I__2806 (
            .O(N__16018),
            .I(\tok.A_stk.tail_94 ));
    CascadeMux I__2805 (
            .O(N__16013),
            .I(N__16010));
    InMux I__2804 (
            .O(N__16010),
            .I(N__16007));
    LocalMux I__2803 (
            .O(N__16007),
            .I(\tok.n5423 ));
    CascadeMux I__2802 (
            .O(N__16004),
            .I(N__16001));
    InMux I__2801 (
            .O(N__16001),
            .I(N__15998));
    LocalMux I__2800 (
            .O(N__15998),
            .I(\tok.n42_adj_751 ));
    InMux I__2799 (
            .O(N__15995),
            .I(N__15992));
    LocalMux I__2798 (
            .O(N__15992),
            .I(N__15987));
    InMux I__2797 (
            .O(N__15991),
            .I(N__15984));
    InMux I__2796 (
            .O(N__15990),
            .I(N__15981));
    Span4Mux_v I__2795 (
            .O(N__15987),
            .I(N__15978));
    LocalMux I__2794 (
            .O(N__15984),
            .I(capture_9));
    LocalMux I__2793 (
            .O(N__15981),
            .I(capture_9));
    Odrv4 I__2792 (
            .O(N__15978),
            .I(capture_9));
    InMux I__2791 (
            .O(N__15971),
            .I(N__15968));
    LocalMux I__2790 (
            .O(N__15968),
            .I(\tok.n2609 ));
    InMux I__2789 (
            .O(N__15965),
            .I(N__15957));
    InMux I__2788 (
            .O(N__15964),
            .I(N__15954));
    InMux I__2787 (
            .O(N__15963),
            .I(N__15950));
    InMux I__2786 (
            .O(N__15962),
            .I(N__15947));
    InMux I__2785 (
            .O(N__15961),
            .I(N__15943));
    InMux I__2784 (
            .O(N__15960),
            .I(N__15940));
    LocalMux I__2783 (
            .O(N__15957),
            .I(N__15935));
    LocalMux I__2782 (
            .O(N__15954),
            .I(N__15935));
    InMux I__2781 (
            .O(N__15953),
            .I(N__15932));
    LocalMux I__2780 (
            .O(N__15950),
            .I(N__15929));
    LocalMux I__2779 (
            .O(N__15947),
            .I(N__15926));
    InMux I__2778 (
            .O(N__15946),
            .I(N__15923));
    LocalMux I__2777 (
            .O(N__15943),
            .I(N__15920));
    LocalMux I__2776 (
            .O(N__15940),
            .I(N__15911));
    Span4Mux_h I__2775 (
            .O(N__15935),
            .I(N__15911));
    LocalMux I__2774 (
            .O(N__15932),
            .I(N__15911));
    Span4Mux_h I__2773 (
            .O(N__15929),
            .I(N__15911));
    Span4Mux_h I__2772 (
            .O(N__15926),
            .I(N__15908));
    LocalMux I__2771 (
            .O(N__15923),
            .I(N__15905));
    Span4Mux_h I__2770 (
            .O(N__15920),
            .I(N__15900));
    Span4Mux_v I__2769 (
            .O(N__15911),
            .I(N__15900));
    Odrv4 I__2768 (
            .O(N__15908),
            .I(\tok.n4_adj_712 ));
    Odrv12 I__2767 (
            .O(N__15905),
            .I(\tok.n4_adj_712 ));
    Odrv4 I__2766 (
            .O(N__15900),
            .I(\tok.n4_adj_712 ));
    CascadeMux I__2765 (
            .O(N__15893),
            .I(\tok.ram.n5577_cascade_ ));
    InMux I__2764 (
            .O(N__15890),
            .I(N__15886));
    CascadeMux I__2763 (
            .O(N__15889),
            .I(N__15883));
    LocalMux I__2762 (
            .O(N__15886),
            .I(N__15879));
    InMux I__2761 (
            .O(N__15883),
            .I(N__15876));
    InMux I__2760 (
            .O(N__15882),
            .I(N__15870));
    Span4Mux_v I__2759 (
            .O(N__15879),
            .I(N__15865));
    LocalMux I__2758 (
            .O(N__15876),
            .I(N__15865));
    InMux I__2757 (
            .O(N__15875),
            .I(N__15862));
    InMux I__2756 (
            .O(N__15874),
            .I(N__15857));
    InMux I__2755 (
            .O(N__15873),
            .I(N__15854));
    LocalMux I__2754 (
            .O(N__15870),
            .I(N__15851));
    Span4Mux_v I__2753 (
            .O(N__15865),
            .I(N__15846));
    LocalMux I__2752 (
            .O(N__15862),
            .I(N__15846));
    InMux I__2751 (
            .O(N__15861),
            .I(N__15843));
    InMux I__2750 (
            .O(N__15860),
            .I(N__15840));
    LocalMux I__2749 (
            .O(N__15857),
            .I(N__15835));
    LocalMux I__2748 (
            .O(N__15854),
            .I(N__15835));
    Span4Mux_v I__2747 (
            .O(N__15851),
            .I(N__15830));
    Span4Mux_h I__2746 (
            .O(N__15846),
            .I(N__15830));
    LocalMux I__2745 (
            .O(N__15843),
            .I(\tok.n101 ));
    LocalMux I__2744 (
            .O(N__15840),
            .I(\tok.n101 ));
    Odrv4 I__2743 (
            .O(N__15835),
            .I(\tok.n101 ));
    Odrv4 I__2742 (
            .O(N__15830),
            .I(\tok.n101 ));
    InMux I__2741 (
            .O(N__15821),
            .I(N__15818));
    LocalMux I__2740 (
            .O(N__15818),
            .I(\tok.n3_adj_672 ));
    InMux I__2739 (
            .O(N__15815),
            .I(N__15809));
    InMux I__2738 (
            .O(N__15814),
            .I(N__15809));
    LocalMux I__2737 (
            .O(N__15809),
            .I(\tok.n14_adj_701 ));
    InMux I__2736 (
            .O(N__15806),
            .I(N__15803));
    LocalMux I__2735 (
            .O(N__15803),
            .I(N__15800));
    Span4Mux_h I__2734 (
            .O(N__15800),
            .I(N__15797));
    Odrv4 I__2733 (
            .O(N__15797),
            .I(\tok.n5429 ));
    InMux I__2732 (
            .O(N__15794),
            .I(N__15791));
    LocalMux I__2731 (
            .O(N__15791),
            .I(\tok.n5406 ));
    CascadeMux I__2730 (
            .O(N__15788),
            .I(\tok.n5433_cascade_ ));
    InMux I__2729 (
            .O(N__15785),
            .I(N__15782));
    LocalMux I__2728 (
            .O(N__15782),
            .I(\tok.n5272 ));
    CascadeMux I__2727 (
            .O(N__15779),
            .I(N__15776));
    InMux I__2726 (
            .O(N__15776),
            .I(N__15773));
    LocalMux I__2725 (
            .O(N__15773),
            .I(N__15770));
    Odrv4 I__2724 (
            .O(N__15770),
            .I(\tok.n10_adj_796 ));
    InMux I__2723 (
            .O(N__15767),
            .I(N__15761));
    InMux I__2722 (
            .O(N__15766),
            .I(N__15761));
    LocalMux I__2721 (
            .O(N__15761),
            .I(\tok.n14_adj_807 ));
    InMux I__2720 (
            .O(N__15758),
            .I(N__15755));
    LocalMux I__2719 (
            .O(N__15755),
            .I(\tok.n5175 ));
    InMux I__2718 (
            .O(N__15752),
            .I(N__15749));
    LocalMux I__2717 (
            .O(N__15749),
            .I(N__15745));
    InMux I__2716 (
            .O(N__15748),
            .I(N__15742));
    Span4Mux_h I__2715 (
            .O(N__15745),
            .I(N__15737));
    LocalMux I__2714 (
            .O(N__15742),
            .I(N__15737));
    Span4Mux_v I__2713 (
            .O(N__15737),
            .I(N__15734));
    Odrv4 I__2712 (
            .O(N__15734),
            .I(n10_adj_866));
    InMux I__2711 (
            .O(N__15731),
            .I(N__15728));
    LocalMux I__2710 (
            .O(N__15728),
            .I(N__15723));
    InMux I__2709 (
            .O(N__15727),
            .I(N__15719));
    InMux I__2708 (
            .O(N__15726),
            .I(N__15716));
    Span12Mux_v I__2707 (
            .O(N__15723),
            .I(N__15713));
    InMux I__2706 (
            .O(N__15722),
            .I(N__15710));
    LocalMux I__2705 (
            .O(N__15719),
            .I(N__15707));
    LocalMux I__2704 (
            .O(N__15716),
            .I(N__15704));
    Odrv12 I__2703 (
            .O(N__15713),
            .I(tc_1));
    LocalMux I__2702 (
            .O(N__15710),
            .I(tc_1));
    Odrv4 I__2701 (
            .O(N__15707),
            .I(tc_1));
    Odrv12 I__2700 (
            .O(N__15704),
            .I(tc_1));
    CascadeMux I__2699 (
            .O(N__15695),
            .I(N__15692));
    InMux I__2698 (
            .O(N__15692),
            .I(N__15689));
    LocalMux I__2697 (
            .O(N__15689),
            .I(N__15686));
    Span4Mux_h I__2696 (
            .O(N__15686),
            .I(N__15683));
    Odrv4 I__2695 (
            .O(N__15683),
            .I(\tok.tc_1 ));
    InMux I__2694 (
            .O(N__15680),
            .I(N__15677));
    LocalMux I__2693 (
            .O(N__15677),
            .I(\tok.n2_adj_808 ));
    CascadeMux I__2692 (
            .O(N__15674),
            .I(N__15668));
    CascadeMux I__2691 (
            .O(N__15673),
            .I(N__15664));
    CascadeMux I__2690 (
            .O(N__15672),
            .I(N__15660));
    InMux I__2689 (
            .O(N__15671),
            .I(N__15647));
    InMux I__2688 (
            .O(N__15668),
            .I(N__15647));
    InMux I__2687 (
            .O(N__15667),
            .I(N__15647));
    InMux I__2686 (
            .O(N__15664),
            .I(N__15647));
    InMux I__2685 (
            .O(N__15663),
            .I(N__15647));
    InMux I__2684 (
            .O(N__15660),
            .I(N__15647));
    LocalMux I__2683 (
            .O(N__15647),
            .I(N__15644));
    Odrv12 I__2682 (
            .O(N__15644),
            .I(\tok.n10_adj_747 ));
    InMux I__2681 (
            .O(N__15641),
            .I(N__15635));
    InMux I__2680 (
            .O(N__15640),
            .I(N__15635));
    LocalMux I__2679 (
            .O(N__15635),
            .I(N__15632));
    Odrv4 I__2678 (
            .O(N__15632),
            .I(\tok.n2635 ));
    InMux I__2677 (
            .O(N__15629),
            .I(N__15612));
    InMux I__2676 (
            .O(N__15628),
            .I(N__15612));
    InMux I__2675 (
            .O(N__15627),
            .I(N__15612));
    InMux I__2674 (
            .O(N__15626),
            .I(N__15595));
    InMux I__2673 (
            .O(N__15625),
            .I(N__15595));
    InMux I__2672 (
            .O(N__15624),
            .I(N__15595));
    InMux I__2671 (
            .O(N__15623),
            .I(N__15595));
    InMux I__2670 (
            .O(N__15622),
            .I(N__15595));
    InMux I__2669 (
            .O(N__15621),
            .I(N__15595));
    InMux I__2668 (
            .O(N__15620),
            .I(N__15595));
    InMux I__2667 (
            .O(N__15619),
            .I(N__15595));
    LocalMux I__2666 (
            .O(N__15612),
            .I(N__15591));
    LocalMux I__2665 (
            .O(N__15595),
            .I(N__15586));
    InMux I__2664 (
            .O(N__15594),
            .I(N__15583));
    Span4Mux_v I__2663 (
            .O(N__15591),
            .I(N__15580));
    InMux I__2662 (
            .O(N__15590),
            .I(N__15575));
    InMux I__2661 (
            .O(N__15589),
            .I(N__15575));
    Odrv4 I__2660 (
            .O(N__15586),
            .I(\tok.n11 ));
    LocalMux I__2659 (
            .O(N__15583),
            .I(\tok.n11 ));
    Odrv4 I__2658 (
            .O(N__15580),
            .I(\tok.n11 ));
    LocalMux I__2657 (
            .O(N__15575),
            .I(\tok.n11 ));
    CascadeMux I__2656 (
            .O(N__15566),
            .I(N__15563));
    InMux I__2655 (
            .O(N__15563),
            .I(N__15551));
    InMux I__2654 (
            .O(N__15562),
            .I(N__15551));
    InMux I__2653 (
            .O(N__15561),
            .I(N__15551));
    InMux I__2652 (
            .O(N__15560),
            .I(N__15551));
    LocalMux I__2651 (
            .O(N__15551),
            .I(N__15548));
    Odrv12 I__2650 (
            .O(N__15548),
            .I(\tok.n2697 ));
    InMux I__2649 (
            .O(N__15545),
            .I(N__15539));
    InMux I__2648 (
            .O(N__15544),
            .I(N__15536));
    InMux I__2647 (
            .O(N__15543),
            .I(N__15532));
    InMux I__2646 (
            .O(N__15542),
            .I(N__15529));
    LocalMux I__2645 (
            .O(N__15539),
            .I(N__15524));
    LocalMux I__2644 (
            .O(N__15536),
            .I(N__15521));
    InMux I__2643 (
            .O(N__15535),
            .I(N__15518));
    LocalMux I__2642 (
            .O(N__15532),
            .I(N__15512));
    LocalMux I__2641 (
            .O(N__15529),
            .I(N__15512));
    InMux I__2640 (
            .O(N__15528),
            .I(N__15509));
    InMux I__2639 (
            .O(N__15527),
            .I(N__15505));
    Span4Mux_v I__2638 (
            .O(N__15524),
            .I(N__15500));
    Span4Mux_s1_h I__2637 (
            .O(N__15521),
            .I(N__15500));
    LocalMux I__2636 (
            .O(N__15518),
            .I(N__15497));
    InMux I__2635 (
            .O(N__15517),
            .I(N__15494));
    Span4Mux_s2_h I__2634 (
            .O(N__15512),
            .I(N__15489));
    LocalMux I__2633 (
            .O(N__15509),
            .I(N__15489));
    InMux I__2632 (
            .O(N__15508),
            .I(N__15486));
    LocalMux I__2631 (
            .O(N__15505),
            .I(N__15483));
    Span4Mux_h I__2630 (
            .O(N__15500),
            .I(N__15476));
    Span4Mux_h I__2629 (
            .O(N__15497),
            .I(N__15476));
    LocalMux I__2628 (
            .O(N__15494),
            .I(N__15476));
    Span4Mux_h I__2627 (
            .O(N__15489),
            .I(N__15471));
    LocalMux I__2626 (
            .O(N__15486),
            .I(N__15471));
    Odrv12 I__2625 (
            .O(N__15483),
            .I(\tok.n15_adj_789 ));
    Odrv4 I__2624 (
            .O(N__15476),
            .I(\tok.n15_adj_789 ));
    Odrv4 I__2623 (
            .O(N__15471),
            .I(\tok.n15_adj_789 ));
    InMux I__2622 (
            .O(N__15464),
            .I(N__15461));
    LocalMux I__2621 (
            .O(N__15461),
            .I(\tok.n2520 ));
    InMux I__2620 (
            .O(N__15458),
            .I(N__15455));
    LocalMux I__2619 (
            .O(N__15455),
            .I(N__15452));
    Span4Mux_v I__2618 (
            .O(N__15452),
            .I(N__15447));
    InMux I__2617 (
            .O(N__15451),
            .I(N__15442));
    InMux I__2616 (
            .O(N__15450),
            .I(N__15442));
    Odrv4 I__2615 (
            .O(N__15447),
            .I(\tok.n10_adj_803 ));
    LocalMux I__2614 (
            .O(N__15442),
            .I(\tok.n10_adj_803 ));
    CascadeMux I__2613 (
            .O(N__15437),
            .I(\tok.n2520_cascade_ ));
    InMux I__2612 (
            .O(N__15434),
            .I(N__15425));
    InMux I__2611 (
            .O(N__15433),
            .I(N__15425));
    InMux I__2610 (
            .O(N__15432),
            .I(N__15425));
    LocalMux I__2609 (
            .O(N__15425),
            .I(N__15420));
    InMux I__2608 (
            .O(N__15424),
            .I(N__15412));
    InMux I__2607 (
            .O(N__15423),
            .I(N__15412));
    Span4Mux_h I__2606 (
            .O(N__15420),
            .I(N__15409));
    InMux I__2605 (
            .O(N__15419),
            .I(N__15402));
    InMux I__2604 (
            .O(N__15418),
            .I(N__15402));
    InMux I__2603 (
            .O(N__15417),
            .I(N__15402));
    LocalMux I__2602 (
            .O(N__15412),
            .I(\tok.n9_adj_802 ));
    Odrv4 I__2601 (
            .O(N__15409),
            .I(\tok.n9_adj_802 ));
    LocalMux I__2600 (
            .O(N__15402),
            .I(\tok.n9_adj_802 ));
    CascadeMux I__2599 (
            .O(N__15395),
            .I(N__15392));
    InMux I__2598 (
            .O(N__15392),
            .I(N__15388));
    InMux I__2597 (
            .O(N__15391),
            .I(N__15385));
    LocalMux I__2596 (
            .O(N__15388),
            .I(N__15382));
    LocalMux I__2595 (
            .O(N__15385),
            .I(N__15379));
    Span4Mux_h I__2594 (
            .O(N__15382),
            .I(N__15376));
    Span4Mux_h I__2593 (
            .O(N__15379),
            .I(N__15371));
    Span4Mux_v I__2592 (
            .O(N__15376),
            .I(N__15371));
    Odrv4 I__2591 (
            .O(N__15371),
            .I(\tok.table_rd_3 ));
    CascadeMux I__2590 (
            .O(N__15368),
            .I(\tok.n2661_cascade_ ));
    InMux I__2589 (
            .O(N__15365),
            .I(N__15362));
    LocalMux I__2588 (
            .O(N__15362),
            .I(\tok.n10_adj_845 ));
    CascadeMux I__2587 (
            .O(N__15359),
            .I(\tok.n9_adj_847_cascade_ ));
    InMux I__2586 (
            .O(N__15356),
            .I(N__15350));
    InMux I__2585 (
            .O(N__15355),
            .I(N__15350));
    LocalMux I__2584 (
            .O(N__15350),
            .I(uart_rx_data_6));
    InMux I__2583 (
            .O(N__15347),
            .I(N__15344));
    LocalMux I__2582 (
            .O(N__15344),
            .I(\tok.n6_adj_843 ));
    CascadeMux I__2581 (
            .O(N__15341),
            .I(\tok.n31_adj_844_cascade_ ));
    InMux I__2580 (
            .O(N__15338),
            .I(N__15332));
    InMux I__2579 (
            .O(N__15337),
            .I(N__15332));
    LocalMux I__2578 (
            .O(N__15332),
            .I(uart_rx_data_3));
    CascadeMux I__2577 (
            .O(N__15329),
            .I(N__15326));
    InMux I__2576 (
            .O(N__15326),
            .I(N__15317));
    InMux I__2575 (
            .O(N__15325),
            .I(N__15317));
    InMux I__2574 (
            .O(N__15324),
            .I(N__15317));
    LocalMux I__2573 (
            .O(N__15317),
            .I(capture_4));
    InMux I__2572 (
            .O(N__15314),
            .I(N__15308));
    InMux I__2571 (
            .O(N__15313),
            .I(N__15303));
    InMux I__2570 (
            .O(N__15312),
            .I(N__15303));
    InMux I__2569 (
            .O(N__15311),
            .I(N__15300));
    LocalMux I__2568 (
            .O(N__15308),
            .I(N__15295));
    LocalMux I__2567 (
            .O(N__15303),
            .I(N__15295));
    LocalMux I__2566 (
            .O(N__15300),
            .I(\tok.tc_plus_1_6 ));
    Odrv12 I__2565 (
            .O(N__15295),
            .I(\tok.tc_plus_1_6 ));
    InMux I__2564 (
            .O(N__15290),
            .I(N__15287));
    LocalMux I__2563 (
            .O(N__15287),
            .I(N__15284));
    Span4Mux_v I__2562 (
            .O(N__15284),
            .I(N__15281));
    Span4Mux_h I__2561 (
            .O(N__15281),
            .I(N__15278));
    Odrv4 I__2560 (
            .O(N__15278),
            .I(\tok.table_wr_data_6 ));
    CascadeMux I__2559 (
            .O(N__15275),
            .I(N__15271));
    InMux I__2558 (
            .O(N__15274),
            .I(N__15266));
    InMux I__2557 (
            .O(N__15271),
            .I(N__15266));
    LocalMux I__2556 (
            .O(N__15266),
            .I(N__15263));
    Span4Mux_h I__2555 (
            .O(N__15263),
            .I(N__15260));
    Odrv4 I__2554 (
            .O(N__15260),
            .I(\tok.key_rd_8 ));
    InMux I__2553 (
            .O(N__15257),
            .I(N__15254));
    LocalMux I__2552 (
            .O(N__15254),
            .I(\tok.n28_adj_755 ));
    CascadeMux I__2551 (
            .O(N__15251),
            .I(\tok.n26_adj_756_cascade_ ));
    InMux I__2550 (
            .O(N__15248),
            .I(N__15245));
    LocalMux I__2549 (
            .O(N__15245),
            .I(\tok.n27_adj_757 ));
    InMux I__2548 (
            .O(N__15242),
            .I(N__15239));
    LocalMux I__2547 (
            .O(N__15239),
            .I(\tok.found_slot_N_145 ));
    CascadeMux I__2546 (
            .O(N__15236),
            .I(N__15226));
    CascadeMux I__2545 (
            .O(N__15235),
            .I(N__15223));
    CascadeMux I__2544 (
            .O(N__15234),
            .I(N__15220));
    CascadeMux I__2543 (
            .O(N__15233),
            .I(N__15217));
    CascadeMux I__2542 (
            .O(N__15232),
            .I(N__15214));
    CascadeMux I__2541 (
            .O(N__15231),
            .I(N__15211));
    CascadeMux I__2540 (
            .O(N__15230),
            .I(N__15208));
    CascadeMux I__2539 (
            .O(N__15229),
            .I(N__15205));
    InMux I__2538 (
            .O(N__15226),
            .I(N__15196));
    InMux I__2537 (
            .O(N__15223),
            .I(N__15196));
    InMux I__2536 (
            .O(N__15220),
            .I(N__15196));
    InMux I__2535 (
            .O(N__15217),
            .I(N__15196));
    InMux I__2534 (
            .O(N__15214),
            .I(N__15187));
    InMux I__2533 (
            .O(N__15211),
            .I(N__15187));
    InMux I__2532 (
            .O(N__15208),
            .I(N__15187));
    InMux I__2531 (
            .O(N__15205),
            .I(N__15187));
    LocalMux I__2530 (
            .O(N__15196),
            .I(N__15180));
    LocalMux I__2529 (
            .O(N__15187),
            .I(N__15180));
    InMux I__2528 (
            .O(N__15186),
            .I(N__15177));
    InMux I__2527 (
            .O(N__15185),
            .I(N__15174));
    Span4Mux_s2_v I__2526 (
            .O(N__15180),
            .I(N__15169));
    LocalMux I__2525 (
            .O(N__15177),
            .I(N__15169));
    LocalMux I__2524 (
            .O(N__15174),
            .I(\tok.found_slot ));
    Odrv4 I__2523 (
            .O(N__15169),
            .I(\tok.found_slot ));
    SRMux I__2522 (
            .O(N__15164),
            .I(N__15160));
    SRMux I__2521 (
            .O(N__15163),
            .I(N__15157));
    LocalMux I__2520 (
            .O(N__15160),
            .I(N__15152));
    LocalMux I__2519 (
            .O(N__15157),
            .I(N__15152));
    Span4Mux_v I__2518 (
            .O(N__15152),
            .I(N__15149));
    Span4Mux_h I__2517 (
            .O(N__15149),
            .I(N__15146));
    Odrv4 I__2516 (
            .O(N__15146),
            .I(\tok.write_slot ));
    InMux I__2515 (
            .O(N__15143),
            .I(N__15137));
    InMux I__2514 (
            .O(N__15142),
            .I(N__15137));
    LocalMux I__2513 (
            .O(N__15137),
            .I(N__15134));
    Span4Mux_h I__2512 (
            .O(N__15134),
            .I(N__15131));
    Odrv4 I__2511 (
            .O(N__15131),
            .I(\tok.key_rd_3 ));
    InMux I__2510 (
            .O(N__15128),
            .I(N__15122));
    InMux I__2509 (
            .O(N__15127),
            .I(N__15122));
    LocalMux I__2508 (
            .O(N__15122),
            .I(N__15119));
    Span4Mux_v I__2507 (
            .O(N__15119),
            .I(N__15116));
    Odrv4 I__2506 (
            .O(N__15116),
            .I(\tok.key_rd_5 ));
    CascadeMux I__2505 (
            .O(N__15113),
            .I(N__15110));
    InMux I__2504 (
            .O(N__15110),
            .I(N__15107));
    LocalMux I__2503 (
            .O(N__15107),
            .I(\tok.n20 ));
    InMux I__2502 (
            .O(N__15104),
            .I(N__15101));
    LocalMux I__2501 (
            .O(N__15101),
            .I(\tok.n18_adj_759 ));
    CascadeMux I__2500 (
            .O(N__15098),
            .I(N__15095));
    InMux I__2499 (
            .O(N__15095),
            .I(N__15089));
    InMux I__2498 (
            .O(N__15094),
            .I(N__15089));
    LocalMux I__2497 (
            .O(N__15089),
            .I(N__15086));
    Span4Mux_h I__2496 (
            .O(N__15086),
            .I(N__15083));
    Odrv4 I__2495 (
            .O(N__15083),
            .I(\tok.key_rd_1 ));
    CascadeMux I__2494 (
            .O(N__15080),
            .I(N__15077));
    InMux I__2493 (
            .O(N__15077),
            .I(N__15071));
    InMux I__2492 (
            .O(N__15076),
            .I(N__15071));
    LocalMux I__2491 (
            .O(N__15071),
            .I(N__15068));
    Span4Mux_h I__2490 (
            .O(N__15068),
            .I(N__15065));
    Odrv4 I__2489 (
            .O(N__15065),
            .I(\tok.key_rd_4 ));
    InMux I__2488 (
            .O(N__15062),
            .I(N__15059));
    LocalMux I__2487 (
            .O(N__15059),
            .I(\tok.n25_adj_758 ));
    InMux I__2486 (
            .O(N__15056),
            .I(N__15050));
    InMux I__2485 (
            .O(N__15055),
            .I(N__15050));
    LocalMux I__2484 (
            .O(N__15050),
            .I(N__15047));
    Span4Mux_h I__2483 (
            .O(N__15047),
            .I(N__15044));
    Odrv4 I__2482 (
            .O(N__15044),
            .I(\tok.key_rd_0 ));
    InMux I__2481 (
            .O(N__15041),
            .I(N__15035));
    InMux I__2480 (
            .O(N__15040),
            .I(N__15035));
    LocalMux I__2479 (
            .O(N__15035),
            .I(N__15032));
    Span4Mux_v I__2478 (
            .O(N__15032),
            .I(N__15029));
    Odrv4 I__2477 (
            .O(N__15029),
            .I(\tok.key_rd_6 ));
    InMux I__2476 (
            .O(N__15026),
            .I(N__15023));
    LocalMux I__2475 (
            .O(N__15023),
            .I(\tok.n5590 ));
    InMux I__2474 (
            .O(N__15020),
            .I(N__15010));
    InMux I__2473 (
            .O(N__15019),
            .I(N__15010));
    InMux I__2472 (
            .O(N__15018),
            .I(N__15010));
    CascadeMux I__2471 (
            .O(N__15017),
            .I(N__15007));
    LocalMux I__2470 (
            .O(N__15010),
            .I(N__15004));
    InMux I__2469 (
            .O(N__15007),
            .I(N__15001));
    Span12Mux_s6_v I__2468 (
            .O(N__15004),
            .I(N__14998));
    LocalMux I__2467 (
            .O(N__15001),
            .I(\tok.c_stk_r_3 ));
    Odrv12 I__2466 (
            .O(N__14998),
            .I(\tok.c_stk_r_3 ));
    CascadeMux I__2465 (
            .O(N__14993),
            .I(\tok.ram.n5580_cascade_ ));
    InMux I__2464 (
            .O(N__14990),
            .I(N__14987));
    LocalMux I__2463 (
            .O(N__14987),
            .I(\tok.n5460 ));
    CascadeMux I__2462 (
            .O(N__14984),
            .I(\tok.n3_adj_659_cascade_ ));
    InMux I__2461 (
            .O(N__14981),
            .I(N__14978));
    LocalMux I__2460 (
            .O(N__14978),
            .I(N__14973));
    InMux I__2459 (
            .O(N__14977),
            .I(N__14968));
    InMux I__2458 (
            .O(N__14976),
            .I(N__14968));
    Span4Mux_v I__2457 (
            .O(N__14973),
            .I(N__14964));
    LocalMux I__2456 (
            .O(N__14968),
            .I(N__14961));
    InMux I__2455 (
            .O(N__14967),
            .I(N__14958));
    Span4Mux_h I__2454 (
            .O(N__14964),
            .I(N__14953));
    Span4Mux_h I__2453 (
            .O(N__14961),
            .I(N__14953));
    LocalMux I__2452 (
            .O(N__14958),
            .I(\tok.tc_plus_1_3 ));
    Odrv4 I__2451 (
            .O(N__14953),
            .I(\tok.tc_plus_1_3 ));
    CascadeMux I__2450 (
            .O(N__14948),
            .I(\tok.n13_adj_660_cascade_ ));
    InMux I__2449 (
            .O(N__14945),
            .I(N__14939));
    InMux I__2448 (
            .O(N__14944),
            .I(N__14939));
    LocalMux I__2447 (
            .O(N__14939),
            .I(N__14936));
    Span4Mux_h I__2446 (
            .O(N__14936),
            .I(N__14933));
    Odrv4 I__2445 (
            .O(N__14933),
            .I(n92_adj_867));
    InMux I__2444 (
            .O(N__14930),
            .I(N__14927));
    LocalMux I__2443 (
            .O(N__14927),
            .I(N__14924));
    Span4Mux_v I__2442 (
            .O(N__14924),
            .I(N__14920));
    InMux I__2441 (
            .O(N__14923),
            .I(N__14917));
    Odrv4 I__2440 (
            .O(N__14920),
            .I(\tok.n17_adj_777 ));
    LocalMux I__2439 (
            .O(N__14917),
            .I(\tok.n17_adj_777 ));
    CascadeMux I__2438 (
            .O(N__14912),
            .I(\tok.n4_adj_778_cascade_ ));
    CascadeMux I__2437 (
            .O(N__14909),
            .I(\tok.n26_adj_760_cascade_ ));
    InMux I__2436 (
            .O(N__14906),
            .I(N__14903));
    LocalMux I__2435 (
            .O(N__14903),
            .I(\tok.n30_adj_761 ));
    CascadeMux I__2434 (
            .O(N__14900),
            .I(\tok.n5587_cascade_ ));
    CascadeMux I__2433 (
            .O(N__14897),
            .I(\tok.n5_cascade_ ));
    InMux I__2432 (
            .O(N__14894),
            .I(N__14891));
    LocalMux I__2431 (
            .O(N__14891),
            .I(\tok.n5 ));
    InMux I__2430 (
            .O(N__14888),
            .I(N__14885));
    LocalMux I__2429 (
            .O(N__14885),
            .I(\tok.n33 ));
    CascadeMux I__2428 (
            .O(N__14882),
            .I(\tok.n27_cascade_ ));
    CascadeMux I__2427 (
            .O(N__14879),
            .I(N__14876));
    CascadeBuf I__2426 (
            .O(N__14876),
            .I(N__14872));
    CascadeMux I__2425 (
            .O(N__14875),
            .I(N__14869));
    CascadeMux I__2424 (
            .O(N__14872),
            .I(N__14866));
    CascadeBuf I__2423 (
            .O(N__14869),
            .I(N__14863));
    InMux I__2422 (
            .O(N__14866),
            .I(N__14860));
    CascadeMux I__2421 (
            .O(N__14863),
            .I(N__14857));
    LocalMux I__2420 (
            .O(N__14860),
            .I(N__14854));
    InMux I__2419 (
            .O(N__14857),
            .I(N__14851));
    Span4Mux_h I__2418 (
            .O(N__14854),
            .I(N__14845));
    LocalMux I__2417 (
            .O(N__14851),
            .I(N__14842));
    InMux I__2416 (
            .O(N__14850),
            .I(N__14839));
    InMux I__2415 (
            .O(N__14849),
            .I(N__14836));
    InMux I__2414 (
            .O(N__14848),
            .I(N__14833));
    Span4Mux_v I__2413 (
            .O(N__14845),
            .I(N__14830));
    Span12Mux_s6_h I__2412 (
            .O(N__14842),
            .I(N__14827));
    LocalMux I__2411 (
            .O(N__14839),
            .I(\tok.idx_0 ));
    LocalMux I__2410 (
            .O(N__14836),
            .I(\tok.idx_0 ));
    LocalMux I__2409 (
            .O(N__14833),
            .I(\tok.idx_0 ));
    Odrv4 I__2408 (
            .O(N__14830),
            .I(\tok.idx_0 ));
    Odrv12 I__2407 (
            .O(N__14827),
            .I(\tok.idx_0 ));
    CascadeMux I__2406 (
            .O(N__14816),
            .I(\tok.n83_adj_652_cascade_ ));
    InMux I__2405 (
            .O(N__14813),
            .I(bfn_6_3_0_));
    InMux I__2404 (
            .O(N__14810),
            .I(\tok.n4747 ));
    InMux I__2403 (
            .O(N__14807),
            .I(\tok.n4748 ));
    InMux I__2402 (
            .O(N__14804),
            .I(\tok.n4749 ));
    CascadeMux I__2401 (
            .O(N__14801),
            .I(N__14798));
    CascadeBuf I__2400 (
            .O(N__14798),
            .I(N__14794));
    CascadeMux I__2399 (
            .O(N__14797),
            .I(N__14791));
    CascadeMux I__2398 (
            .O(N__14794),
            .I(N__14788));
    CascadeBuf I__2397 (
            .O(N__14791),
            .I(N__14785));
    InMux I__2396 (
            .O(N__14788),
            .I(N__14782));
    CascadeMux I__2395 (
            .O(N__14785),
            .I(N__14779));
    LocalMux I__2394 (
            .O(N__14782),
            .I(N__14775));
    InMux I__2393 (
            .O(N__14779),
            .I(N__14772));
    CascadeMux I__2392 (
            .O(N__14778),
            .I(N__14769));
    Span4Mux_h I__2391 (
            .O(N__14775),
            .I(N__14764));
    LocalMux I__2390 (
            .O(N__14772),
            .I(N__14761));
    InMux I__2389 (
            .O(N__14769),
            .I(N__14758));
    InMux I__2388 (
            .O(N__14768),
            .I(N__14755));
    InMux I__2387 (
            .O(N__14767),
            .I(N__14752));
    Span4Mux_v I__2386 (
            .O(N__14764),
            .I(N__14749));
    Span12Mux_s5_h I__2385 (
            .O(N__14761),
            .I(N__14746));
    LocalMux I__2384 (
            .O(N__14758),
            .I(\tok.idx_4 ));
    LocalMux I__2383 (
            .O(N__14755),
            .I(\tok.idx_4 ));
    LocalMux I__2382 (
            .O(N__14752),
            .I(\tok.idx_4 ));
    Odrv4 I__2381 (
            .O(N__14749),
            .I(\tok.idx_4 ));
    Odrv12 I__2380 (
            .O(N__14746),
            .I(\tok.idx_4 ));
    InMux I__2379 (
            .O(N__14735),
            .I(N__14732));
    LocalMux I__2378 (
            .O(N__14732),
            .I(\tok.n33_adj_819 ));
    InMux I__2377 (
            .O(N__14729),
            .I(\tok.n4750 ));
    CascadeMux I__2376 (
            .O(N__14726),
            .I(N__14723));
    CascadeBuf I__2375 (
            .O(N__14723),
            .I(N__14719));
    CascadeMux I__2374 (
            .O(N__14722),
            .I(N__14716));
    CascadeMux I__2373 (
            .O(N__14719),
            .I(N__14713));
    CascadeBuf I__2372 (
            .O(N__14716),
            .I(N__14710));
    InMux I__2371 (
            .O(N__14713),
            .I(N__14707));
    CascadeMux I__2370 (
            .O(N__14710),
            .I(N__14704));
    LocalMux I__2369 (
            .O(N__14707),
            .I(N__14701));
    InMux I__2368 (
            .O(N__14704),
            .I(N__14698));
    Span4Mux_v I__2367 (
            .O(N__14701),
            .I(N__14692));
    LocalMux I__2366 (
            .O(N__14698),
            .I(N__14689));
    InMux I__2365 (
            .O(N__14697),
            .I(N__14686));
    InMux I__2364 (
            .O(N__14696),
            .I(N__14683));
    InMux I__2363 (
            .O(N__14695),
            .I(N__14680));
    Span4Mux_v I__2362 (
            .O(N__14692),
            .I(N__14677));
    Span4Mux_h I__2361 (
            .O(N__14689),
            .I(N__14674));
    LocalMux I__2360 (
            .O(N__14686),
            .I(N__14665));
    LocalMux I__2359 (
            .O(N__14683),
            .I(N__14665));
    LocalMux I__2358 (
            .O(N__14680),
            .I(N__14665));
    Span4Mux_s2_v I__2357 (
            .O(N__14677),
            .I(N__14665));
    Span4Mux_v I__2356 (
            .O(N__14674),
            .I(N__14662));
    Odrv4 I__2355 (
            .O(N__14665),
            .I(\tok.idx_5 ));
    Odrv4 I__2354 (
            .O(N__14662),
            .I(\tok.idx_5 ));
    InMux I__2353 (
            .O(N__14657),
            .I(N__14654));
    LocalMux I__2352 (
            .O(N__14654),
            .I(\tok.n33_adj_811 ));
    InMux I__2351 (
            .O(N__14651),
            .I(\tok.n4751 ));
    CascadeMux I__2350 (
            .O(N__14648),
            .I(N__14644));
    CascadeMux I__2349 (
            .O(N__14647),
            .I(N__14641));
    CascadeBuf I__2348 (
            .O(N__14644),
            .I(N__14638));
    CascadeBuf I__2347 (
            .O(N__14641),
            .I(N__14635));
    CascadeMux I__2346 (
            .O(N__14638),
            .I(N__14632));
    CascadeMux I__2345 (
            .O(N__14635),
            .I(N__14629));
    InMux I__2344 (
            .O(N__14632),
            .I(N__14626));
    InMux I__2343 (
            .O(N__14629),
            .I(N__14623));
    LocalMux I__2342 (
            .O(N__14626),
            .I(N__14619));
    LocalMux I__2341 (
            .O(N__14623),
            .I(N__14616));
    InMux I__2340 (
            .O(N__14622),
            .I(N__14611));
    Span4Mux_v I__2339 (
            .O(N__14619),
            .I(N__14608));
    Span4Mux_h I__2338 (
            .O(N__14616),
            .I(N__14605));
    InMux I__2337 (
            .O(N__14615),
            .I(N__14602));
    InMux I__2336 (
            .O(N__14614),
            .I(N__14599));
    LocalMux I__2335 (
            .O(N__14611),
            .I(N__14594));
    Span4Mux_v I__2334 (
            .O(N__14608),
            .I(N__14594));
    Span4Mux_v I__2333 (
            .O(N__14605),
            .I(N__14591));
    LocalMux I__2332 (
            .O(N__14602),
            .I(\tok.idx_6 ));
    LocalMux I__2331 (
            .O(N__14599),
            .I(\tok.idx_6 ));
    Odrv4 I__2330 (
            .O(N__14594),
            .I(\tok.idx_6 ));
    Odrv4 I__2329 (
            .O(N__14591),
            .I(\tok.idx_6 ));
    InMux I__2328 (
            .O(N__14582),
            .I(N__14579));
    LocalMux I__2327 (
            .O(N__14579),
            .I(\tok.n33_adj_804 ));
    InMux I__2326 (
            .O(N__14576),
            .I(\tok.n4752 ));
    CascadeMux I__2325 (
            .O(N__14573),
            .I(N__14569));
    CascadeMux I__2324 (
            .O(N__14572),
            .I(N__14566));
    CascadeBuf I__2323 (
            .O(N__14569),
            .I(N__14563));
    CascadeBuf I__2322 (
            .O(N__14566),
            .I(N__14560));
    CascadeMux I__2321 (
            .O(N__14563),
            .I(N__14557));
    CascadeMux I__2320 (
            .O(N__14560),
            .I(N__14554));
    InMux I__2319 (
            .O(N__14557),
            .I(N__14549));
    InMux I__2318 (
            .O(N__14554),
            .I(N__14546));
    InMux I__2317 (
            .O(N__14553),
            .I(N__14542));
    InMux I__2316 (
            .O(N__14552),
            .I(N__14539));
    LocalMux I__2315 (
            .O(N__14549),
            .I(N__14534));
    LocalMux I__2314 (
            .O(N__14546),
            .I(N__14534));
    InMux I__2313 (
            .O(N__14545),
            .I(N__14531));
    LocalMux I__2312 (
            .O(N__14542),
            .I(N__14526));
    LocalMux I__2311 (
            .O(N__14539),
            .I(N__14526));
    Span12Mux_s11_v I__2310 (
            .O(N__14534),
            .I(N__14523));
    LocalMux I__2309 (
            .O(N__14531),
            .I(\tok.idx_7 ));
    Odrv4 I__2308 (
            .O(N__14526),
            .I(\tok.idx_7 ));
    Odrv12 I__2307 (
            .O(N__14523),
            .I(\tok.idx_7 ));
    InMux I__2306 (
            .O(N__14516),
            .I(\tok.n4753 ));
    InMux I__2305 (
            .O(N__14513),
            .I(N__14510));
    LocalMux I__2304 (
            .O(N__14510),
            .I(\tok.n33_adj_801 ));
    InMux I__2303 (
            .O(N__14507),
            .I(N__14504));
    LocalMux I__2302 (
            .O(N__14504),
            .I(N__14501));
    Odrv4 I__2301 (
            .O(N__14501),
            .I(reset_c));
    CascadeMux I__2300 (
            .O(N__14498),
            .I(N__14495));
    InMux I__2299 (
            .O(N__14495),
            .I(N__14489));
    InMux I__2298 (
            .O(N__14494),
            .I(N__14489));
    LocalMux I__2297 (
            .O(N__14489),
            .I(\tok.A_stk.tail_16 ));
    InMux I__2296 (
            .O(N__14486),
            .I(N__14480));
    InMux I__2295 (
            .O(N__14485),
            .I(N__14480));
    LocalMux I__2294 (
            .O(N__14480),
            .I(\tok.A_stk.tail_32 ));
    InMux I__2293 (
            .O(N__14477),
            .I(N__14471));
    InMux I__2292 (
            .O(N__14476),
            .I(N__14471));
    LocalMux I__2291 (
            .O(N__14471),
            .I(\tok.A_stk.tail_48 ));
    InMux I__2290 (
            .O(N__14468),
            .I(N__14462));
    InMux I__2289 (
            .O(N__14467),
            .I(N__14462));
    LocalMux I__2288 (
            .O(N__14462),
            .I(\tok.A_stk.tail_64 ));
    CascadeMux I__2287 (
            .O(N__14459),
            .I(N__14455));
    InMux I__2286 (
            .O(N__14458),
            .I(N__14452));
    InMux I__2285 (
            .O(N__14455),
            .I(N__14449));
    LocalMux I__2284 (
            .O(N__14452),
            .I(N__14444));
    LocalMux I__2283 (
            .O(N__14449),
            .I(N__14444));
    Odrv4 I__2282 (
            .O(N__14444),
            .I(tail_112));
    InMux I__2281 (
            .O(N__14441),
            .I(N__14435));
    InMux I__2280 (
            .O(N__14440),
            .I(N__14435));
    LocalMux I__2279 (
            .O(N__14435),
            .I(\tok.A_stk.tail_80 ));
    CascadeMux I__2278 (
            .O(N__14432),
            .I(N__14428));
    InMux I__2277 (
            .O(N__14431),
            .I(N__14425));
    InMux I__2276 (
            .O(N__14428),
            .I(N__14422));
    LocalMux I__2275 (
            .O(N__14425),
            .I(tail_96));
    LocalMux I__2274 (
            .O(N__14422),
            .I(tail_96));
    InMux I__2273 (
            .O(N__14417),
            .I(N__14411));
    InMux I__2272 (
            .O(N__14416),
            .I(N__14411));
    LocalMux I__2271 (
            .O(N__14411),
            .I(\tok.A_stk.tail_0 ));
    InMux I__2270 (
            .O(N__14408),
            .I(N__14405));
    LocalMux I__2269 (
            .O(N__14405),
            .I(N__14402));
    Span4Mux_h I__2268 (
            .O(N__14402),
            .I(N__14398));
    CascadeMux I__2267 (
            .O(N__14401),
            .I(N__14395));
    Span4Mux_v I__2266 (
            .O(N__14398),
            .I(N__14392));
    InMux I__2265 (
            .O(N__14395),
            .I(N__14389));
    Span4Mux_v I__2264 (
            .O(N__14392),
            .I(N__14386));
    LocalMux I__2263 (
            .O(N__14389),
            .I(sender_9));
    Odrv4 I__2262 (
            .O(N__14386),
            .I(sender_9));
    SRMux I__2261 (
            .O(N__14381),
            .I(N__14378));
    LocalMux I__2260 (
            .O(N__14378),
            .I(N__14375));
    Span4Mux_s3_h I__2259 (
            .O(N__14375),
            .I(N__14362));
    InMux I__2258 (
            .O(N__14374),
            .I(N__14357));
    InMux I__2257 (
            .O(N__14373),
            .I(N__14357));
    InMux I__2256 (
            .O(N__14372),
            .I(N__14342));
    InMux I__2255 (
            .O(N__14371),
            .I(N__14342));
    InMux I__2254 (
            .O(N__14370),
            .I(N__14342));
    InMux I__2253 (
            .O(N__14369),
            .I(N__14342));
    InMux I__2252 (
            .O(N__14368),
            .I(N__14342));
    InMux I__2251 (
            .O(N__14367),
            .I(N__14342));
    InMux I__2250 (
            .O(N__14366),
            .I(N__14342));
    InMux I__2249 (
            .O(N__14365),
            .I(N__14339));
    Span4Mux_v I__2248 (
            .O(N__14362),
            .I(N__14336));
    LocalMux I__2247 (
            .O(N__14357),
            .I(N__14333));
    LocalMux I__2246 (
            .O(N__14342),
            .I(N__14329));
    LocalMux I__2245 (
            .O(N__14339),
            .I(N__14326));
    Span4Mux_v I__2244 (
            .O(N__14336),
            .I(N__14321));
    Span4Mux_v I__2243 (
            .O(N__14333),
            .I(N__14321));
    InMux I__2242 (
            .O(N__14332),
            .I(N__14318));
    Span4Mux_v I__2241 (
            .O(N__14329),
            .I(N__14313));
    Span4Mux_h I__2240 (
            .O(N__14326),
            .I(N__14313));
    Odrv4 I__2239 (
            .O(N__14321),
            .I(n23));
    LocalMux I__2238 (
            .O(N__14318),
            .I(n23));
    Odrv4 I__2237 (
            .O(N__14313),
            .I(n23));
    InMux I__2236 (
            .O(N__14306),
            .I(N__14303));
    LocalMux I__2235 (
            .O(N__14303),
            .I(\tok.uart.sender_8 ));
    CEMux I__2234 (
            .O(N__14300),
            .I(N__14297));
    LocalMux I__2233 (
            .O(N__14297),
            .I(N__14294));
    Span4Mux_h I__2232 (
            .O(N__14294),
            .I(N__14290));
    CEMux I__2231 (
            .O(N__14293),
            .I(N__14287));
    Span4Mux_v I__2230 (
            .O(N__14290),
            .I(N__14284));
    LocalMux I__2229 (
            .O(N__14287),
            .I(N__14281));
    Span4Mux_s2_h I__2228 (
            .O(N__14284),
            .I(N__14278));
    Span12Mux_s4_v I__2227 (
            .O(N__14281),
            .I(N__14275));
    Odrv4 I__2226 (
            .O(N__14278),
            .I(\tok.uart.n1017 ));
    Odrv12 I__2225 (
            .O(N__14275),
            .I(\tok.uart.n1017 ));
    InMux I__2224 (
            .O(N__14270),
            .I(N__14266));
    InMux I__2223 (
            .O(N__14269),
            .I(N__14261));
    LocalMux I__2222 (
            .O(N__14266),
            .I(N__14257));
    InMux I__2221 (
            .O(N__14265),
            .I(N__14252));
    InMux I__2220 (
            .O(N__14264),
            .I(N__14248));
    LocalMux I__2219 (
            .O(N__14261),
            .I(N__14245));
    InMux I__2218 (
            .O(N__14260),
            .I(N__14242));
    Span4Mux_s3_v I__2217 (
            .O(N__14257),
            .I(N__14239));
    InMux I__2216 (
            .O(N__14256),
            .I(N__14236));
    InMux I__2215 (
            .O(N__14255),
            .I(N__14233));
    LocalMux I__2214 (
            .O(N__14252),
            .I(N__14230));
    InMux I__2213 (
            .O(N__14251),
            .I(N__14227));
    LocalMux I__2212 (
            .O(N__14248),
            .I(N__14220));
    Span4Mux_h I__2211 (
            .O(N__14245),
            .I(N__14220));
    LocalMux I__2210 (
            .O(N__14242),
            .I(N__14220));
    Span4Mux_h I__2209 (
            .O(N__14239),
            .I(N__14213));
    LocalMux I__2208 (
            .O(N__14236),
            .I(N__14213));
    LocalMux I__2207 (
            .O(N__14233),
            .I(N__14213));
    Odrv4 I__2206 (
            .O(N__14230),
            .I(\tok.C_stk.n602 ));
    LocalMux I__2205 (
            .O(N__14227),
            .I(\tok.C_stk.n602 ));
    Odrv4 I__2204 (
            .O(N__14220),
            .I(\tok.C_stk.n602 ));
    Odrv4 I__2203 (
            .O(N__14213),
            .I(\tok.C_stk.n602 ));
    InMux I__2202 (
            .O(N__14204),
            .I(N__14201));
    LocalMux I__2201 (
            .O(N__14201),
            .I(N__14198));
    IoSpan4Mux I__2200 (
            .O(N__14198),
            .I(N__14192));
    InMux I__2199 (
            .O(N__14197),
            .I(N__14189));
    InMux I__2198 (
            .O(N__14196),
            .I(N__14182));
    CascadeMux I__2197 (
            .O(N__14195),
            .I(N__14179));
    Span4Mux_s3_v I__2196 (
            .O(N__14192),
            .I(N__14174));
    LocalMux I__2195 (
            .O(N__14189),
            .I(N__14174));
    InMux I__2194 (
            .O(N__14188),
            .I(N__14171));
    InMux I__2193 (
            .O(N__14187),
            .I(N__14168));
    InMux I__2192 (
            .O(N__14186),
            .I(N__14165));
    InMux I__2191 (
            .O(N__14185),
            .I(N__14161));
    LocalMux I__2190 (
            .O(N__14182),
            .I(N__14158));
    InMux I__2189 (
            .O(N__14179),
            .I(N__14155));
    Span4Mux_v I__2188 (
            .O(N__14174),
            .I(N__14146));
    LocalMux I__2187 (
            .O(N__14171),
            .I(N__14146));
    LocalMux I__2186 (
            .O(N__14168),
            .I(N__14146));
    LocalMux I__2185 (
            .O(N__14165),
            .I(N__14146));
    InMux I__2184 (
            .O(N__14164),
            .I(N__14143));
    LocalMux I__2183 (
            .O(N__14161),
            .I(N__14140));
    Span4Mux_v I__2182 (
            .O(N__14158),
            .I(N__14135));
    LocalMux I__2181 (
            .O(N__14155),
            .I(N__14135));
    Span4Mux_h I__2180 (
            .O(N__14146),
            .I(N__14132));
    LocalMux I__2179 (
            .O(N__14143),
            .I(N__14129));
    Span4Mux_v I__2178 (
            .O(N__14140),
            .I(N__14124));
    Span4Mux_h I__2177 (
            .O(N__14135),
            .I(N__14124));
    Odrv4 I__2176 (
            .O(N__14132),
            .I(\tok.n241 ));
    Odrv12 I__2175 (
            .O(N__14129),
            .I(\tok.n241 ));
    Odrv4 I__2174 (
            .O(N__14124),
            .I(\tok.n241 ));
    CascadeMux I__2173 (
            .O(N__14117),
            .I(\tok.C_stk.n5438_cascade_ ));
    InMux I__2172 (
            .O(N__14114),
            .I(N__14109));
    CascadeMux I__2171 (
            .O(N__14113),
            .I(N__14106));
    InMux I__2170 (
            .O(N__14112),
            .I(N__14102));
    LocalMux I__2169 (
            .O(N__14109),
            .I(N__14099));
    InMux I__2168 (
            .O(N__14106),
            .I(N__14094));
    InMux I__2167 (
            .O(N__14105),
            .I(N__14094));
    LocalMux I__2166 (
            .O(N__14102),
            .I(N__14091));
    Odrv12 I__2165 (
            .O(N__14099),
            .I(tc_6));
    LocalMux I__2164 (
            .O(N__14094),
            .I(tc_6));
    Odrv4 I__2163 (
            .O(N__14091),
            .I(tc_6));
    CascadeMux I__2162 (
            .O(N__14084),
            .I(N__14080));
    InMux I__2161 (
            .O(N__14083),
            .I(N__14076));
    InMux I__2160 (
            .O(N__14080),
            .I(N__14071));
    InMux I__2159 (
            .O(N__14079),
            .I(N__14071));
    LocalMux I__2158 (
            .O(N__14076),
            .I(N__14065));
    LocalMux I__2157 (
            .O(N__14071),
            .I(N__14065));
    InMux I__2156 (
            .O(N__14070),
            .I(N__14062));
    Span4Mux_v I__2155 (
            .O(N__14065),
            .I(N__14059));
    LocalMux I__2154 (
            .O(N__14062),
            .I(\tok.c_stk_r_6 ));
    Odrv4 I__2153 (
            .O(N__14059),
            .I(\tok.c_stk_r_6 ));
    InMux I__2152 (
            .O(N__14054),
            .I(N__14048));
    InMux I__2151 (
            .O(N__14053),
            .I(N__14048));
    LocalMux I__2150 (
            .O(N__14048),
            .I(\tok.C_stk.tail_6 ));
    CascadeMux I__2149 (
            .O(N__14045),
            .I(N__14041));
    InMux I__2148 (
            .O(N__14044),
            .I(N__13991));
    InMux I__2147 (
            .O(N__14041),
            .I(N__13988));
    InMux I__2146 (
            .O(N__14040),
            .I(N__13983));
    InMux I__2145 (
            .O(N__14039),
            .I(N__13983));
    InMux I__2144 (
            .O(N__14038),
            .I(N__13980));
    InMux I__2143 (
            .O(N__14037),
            .I(N__13963));
    InMux I__2142 (
            .O(N__14036),
            .I(N__13963));
    InMux I__2141 (
            .O(N__14035),
            .I(N__13963));
    InMux I__2140 (
            .O(N__14034),
            .I(N__13963));
    InMux I__2139 (
            .O(N__14033),
            .I(N__13963));
    InMux I__2138 (
            .O(N__14032),
            .I(N__13963));
    InMux I__2137 (
            .O(N__14031),
            .I(N__13950));
    InMux I__2136 (
            .O(N__14030),
            .I(N__13950));
    InMux I__2135 (
            .O(N__14029),
            .I(N__13950));
    InMux I__2134 (
            .O(N__14028),
            .I(N__13950));
    InMux I__2133 (
            .O(N__14027),
            .I(N__13950));
    InMux I__2132 (
            .O(N__14026),
            .I(N__13950));
    InMux I__2131 (
            .O(N__14025),
            .I(N__13943));
    InMux I__2130 (
            .O(N__14024),
            .I(N__13943));
    InMux I__2129 (
            .O(N__14023),
            .I(N__13943));
    InMux I__2128 (
            .O(N__14022),
            .I(N__13930));
    InMux I__2127 (
            .O(N__14021),
            .I(N__13930));
    InMux I__2126 (
            .O(N__14020),
            .I(N__13930));
    InMux I__2125 (
            .O(N__14019),
            .I(N__13930));
    InMux I__2124 (
            .O(N__14018),
            .I(N__13930));
    InMux I__2123 (
            .O(N__14017),
            .I(N__13930));
    InMux I__2122 (
            .O(N__14016),
            .I(N__13921));
    InMux I__2121 (
            .O(N__14015),
            .I(N__13921));
    InMux I__2120 (
            .O(N__14014),
            .I(N__13921));
    InMux I__2119 (
            .O(N__14013),
            .I(N__13921));
    InMux I__2118 (
            .O(N__14012),
            .I(N__13908));
    InMux I__2117 (
            .O(N__14011),
            .I(N__13908));
    InMux I__2116 (
            .O(N__14010),
            .I(N__13908));
    InMux I__2115 (
            .O(N__14009),
            .I(N__13908));
    InMux I__2114 (
            .O(N__14008),
            .I(N__13908));
    InMux I__2113 (
            .O(N__14007),
            .I(N__13908));
    InMux I__2112 (
            .O(N__14006),
            .I(N__13893));
    InMux I__2111 (
            .O(N__14005),
            .I(N__13880));
    InMux I__2110 (
            .O(N__14004),
            .I(N__13880));
    InMux I__2109 (
            .O(N__14003),
            .I(N__13880));
    InMux I__2108 (
            .O(N__14002),
            .I(N__13880));
    InMux I__2107 (
            .O(N__14001),
            .I(N__13880));
    InMux I__2106 (
            .O(N__14000),
            .I(N__13880));
    InMux I__2105 (
            .O(N__13999),
            .I(N__13867));
    InMux I__2104 (
            .O(N__13998),
            .I(N__13867));
    InMux I__2103 (
            .O(N__13997),
            .I(N__13867));
    InMux I__2102 (
            .O(N__13996),
            .I(N__13867));
    InMux I__2101 (
            .O(N__13995),
            .I(N__13867));
    InMux I__2100 (
            .O(N__13994),
            .I(N__13867));
    LocalMux I__2099 (
            .O(N__13991),
            .I(N__13864));
    LocalMux I__2098 (
            .O(N__13988),
            .I(N__13859));
    LocalMux I__2097 (
            .O(N__13983),
            .I(N__13859));
    LocalMux I__2096 (
            .O(N__13980),
            .I(N__13856));
    InMux I__2095 (
            .O(N__13979),
            .I(N__13847));
    InMux I__2094 (
            .O(N__13978),
            .I(N__13847));
    InMux I__2093 (
            .O(N__13977),
            .I(N__13847));
    InMux I__2092 (
            .O(N__13976),
            .I(N__13847));
    LocalMux I__2091 (
            .O(N__13963),
            .I(N__13842));
    LocalMux I__2090 (
            .O(N__13950),
            .I(N__13842));
    LocalMux I__2089 (
            .O(N__13943),
            .I(N__13839));
    LocalMux I__2088 (
            .O(N__13930),
            .I(N__13836));
    LocalMux I__2087 (
            .O(N__13921),
            .I(N__13833));
    LocalMux I__2086 (
            .O(N__13908),
            .I(N__13830));
    InMux I__2085 (
            .O(N__13907),
            .I(N__13817));
    InMux I__2084 (
            .O(N__13906),
            .I(N__13817));
    InMux I__2083 (
            .O(N__13905),
            .I(N__13817));
    InMux I__2082 (
            .O(N__13904),
            .I(N__13817));
    InMux I__2081 (
            .O(N__13903),
            .I(N__13817));
    InMux I__2080 (
            .O(N__13902),
            .I(N__13817));
    InMux I__2079 (
            .O(N__13901),
            .I(N__13804));
    InMux I__2078 (
            .O(N__13900),
            .I(N__13804));
    InMux I__2077 (
            .O(N__13899),
            .I(N__13804));
    InMux I__2076 (
            .O(N__13898),
            .I(N__13804));
    InMux I__2075 (
            .O(N__13897),
            .I(N__13804));
    InMux I__2074 (
            .O(N__13896),
            .I(N__13804));
    LocalMux I__2073 (
            .O(N__13893),
            .I(N__13801));
    LocalMux I__2072 (
            .O(N__13880),
            .I(N__13794));
    LocalMux I__2071 (
            .O(N__13867),
            .I(N__13794));
    Span4Mux_v I__2070 (
            .O(N__13864),
            .I(N__13794));
    Span4Mux_v I__2069 (
            .O(N__13859),
            .I(N__13785));
    Span4Mux_s1_h I__2068 (
            .O(N__13856),
            .I(N__13785));
    LocalMux I__2067 (
            .O(N__13847),
            .I(N__13785));
    Span4Mux_v I__2066 (
            .O(N__13842),
            .I(N__13785));
    Span4Mux_h I__2065 (
            .O(N__13839),
            .I(N__13778));
    Span4Mux_h I__2064 (
            .O(N__13836),
            .I(N__13778));
    Span4Mux_h I__2063 (
            .O(N__13833),
            .I(N__13778));
    Span4Mux_v I__2062 (
            .O(N__13830),
            .I(N__13773));
    LocalMux I__2061 (
            .O(N__13817),
            .I(N__13773));
    LocalMux I__2060 (
            .O(N__13804),
            .I(N__13770));
    Span4Mux_v I__2059 (
            .O(N__13801),
            .I(N__13765));
    Span4Mux_v I__2058 (
            .O(N__13794),
            .I(N__13765));
    Span4Mux_h I__2057 (
            .O(N__13785),
            .I(N__13762));
    Span4Mux_v I__2056 (
            .O(N__13778),
            .I(N__13757));
    Span4Mux_h I__2055 (
            .O(N__13773),
            .I(N__13757));
    Odrv4 I__2054 (
            .O(N__13770),
            .I(\tok.n2515 ));
    Odrv4 I__2053 (
            .O(N__13765),
            .I(\tok.n2515 ));
    Odrv4 I__2052 (
            .O(N__13762),
            .I(\tok.n2515 ));
    Odrv4 I__2051 (
            .O(N__13757),
            .I(\tok.n2515 ));
    InMux I__2050 (
            .O(N__13748),
            .I(N__13742));
    InMux I__2049 (
            .O(N__13747),
            .I(N__13742));
    LocalMux I__2048 (
            .O(N__13742),
            .I(\tok.tail_14 ));
    CascadeMux I__2047 (
            .O(N__13739),
            .I(N__13736));
    InMux I__2046 (
            .O(N__13736),
            .I(N__13733));
    LocalMux I__2045 (
            .O(N__13733),
            .I(N__13729));
    InMux I__2044 (
            .O(N__13732),
            .I(N__13726));
    Odrv4 I__2043 (
            .O(N__13729),
            .I(\tok.tail_30 ));
    LocalMux I__2042 (
            .O(N__13726),
            .I(\tok.tail_30 ));
    CascadeMux I__2041 (
            .O(N__13721),
            .I(N__13717));
    InMux I__2040 (
            .O(N__13720),
            .I(N__13708));
    InMux I__2039 (
            .O(N__13717),
            .I(N__13703));
    InMux I__2038 (
            .O(N__13716),
            .I(N__13703));
    CascadeMux I__2037 (
            .O(N__13715),
            .I(N__13700));
    CascadeMux I__2036 (
            .O(N__13714),
            .I(N__13697));
    CascadeMux I__2035 (
            .O(N__13713),
            .I(N__13678));
    CascadeMux I__2034 (
            .O(N__13712),
            .I(N__13675));
    CascadeMux I__2033 (
            .O(N__13711),
            .I(N__13672));
    LocalMux I__2032 (
            .O(N__13708),
            .I(N__13658));
    LocalMux I__2031 (
            .O(N__13703),
            .I(N__13658));
    InMux I__2030 (
            .O(N__13700),
            .I(N__13649));
    InMux I__2029 (
            .O(N__13697),
            .I(N__13649));
    InMux I__2028 (
            .O(N__13696),
            .I(N__13649));
    InMux I__2027 (
            .O(N__13695),
            .I(N__13649));
    InMux I__2026 (
            .O(N__13694),
            .I(N__13639));
    InMux I__2025 (
            .O(N__13693),
            .I(N__13636));
    CascadeMux I__2024 (
            .O(N__13692),
            .I(N__13628));
    CascadeMux I__2023 (
            .O(N__13691),
            .I(N__13624));
    CascadeMux I__2022 (
            .O(N__13690),
            .I(N__13619));
    CascadeMux I__2021 (
            .O(N__13689),
            .I(N__13616));
    CascadeMux I__2020 (
            .O(N__13688),
            .I(N__13613));
    InMux I__2019 (
            .O(N__13687),
            .I(N__13590));
    InMux I__2018 (
            .O(N__13686),
            .I(N__13590));
    InMux I__2017 (
            .O(N__13685),
            .I(N__13590));
    InMux I__2016 (
            .O(N__13684),
            .I(N__13590));
    InMux I__2015 (
            .O(N__13683),
            .I(N__13583));
    InMux I__2014 (
            .O(N__13682),
            .I(N__13583));
    InMux I__2013 (
            .O(N__13681),
            .I(N__13583));
    InMux I__2012 (
            .O(N__13678),
            .I(N__13570));
    InMux I__2011 (
            .O(N__13675),
            .I(N__13570));
    InMux I__2010 (
            .O(N__13672),
            .I(N__13570));
    InMux I__2009 (
            .O(N__13671),
            .I(N__13570));
    InMux I__2008 (
            .O(N__13670),
            .I(N__13570));
    InMux I__2007 (
            .O(N__13669),
            .I(N__13570));
    InMux I__2006 (
            .O(N__13668),
            .I(N__13557));
    InMux I__2005 (
            .O(N__13667),
            .I(N__13557));
    InMux I__2004 (
            .O(N__13666),
            .I(N__13557));
    InMux I__2003 (
            .O(N__13665),
            .I(N__13557));
    InMux I__2002 (
            .O(N__13664),
            .I(N__13557));
    InMux I__2001 (
            .O(N__13663),
            .I(N__13557));
    Span4Mux_h I__2000 (
            .O(N__13658),
            .I(N__13552));
    LocalMux I__1999 (
            .O(N__13649),
            .I(N__13552));
    InMux I__1998 (
            .O(N__13648),
            .I(N__13546));
    InMux I__1997 (
            .O(N__13647),
            .I(N__13533));
    InMux I__1996 (
            .O(N__13646),
            .I(N__13533));
    InMux I__1995 (
            .O(N__13645),
            .I(N__13533));
    InMux I__1994 (
            .O(N__13644),
            .I(N__13533));
    InMux I__1993 (
            .O(N__13643),
            .I(N__13533));
    InMux I__1992 (
            .O(N__13642),
            .I(N__13533));
    LocalMux I__1991 (
            .O(N__13639),
            .I(N__13530));
    LocalMux I__1990 (
            .O(N__13636),
            .I(N__13527));
    InMux I__1989 (
            .O(N__13635),
            .I(N__13520));
    InMux I__1988 (
            .O(N__13634),
            .I(N__13520));
    InMux I__1987 (
            .O(N__13633),
            .I(N__13520));
    InMux I__1986 (
            .O(N__13632),
            .I(N__13515));
    InMux I__1985 (
            .O(N__13631),
            .I(N__13515));
    InMux I__1984 (
            .O(N__13628),
            .I(N__13512));
    InMux I__1983 (
            .O(N__13627),
            .I(N__13503));
    InMux I__1982 (
            .O(N__13624),
            .I(N__13503));
    InMux I__1981 (
            .O(N__13623),
            .I(N__13503));
    InMux I__1980 (
            .O(N__13622),
            .I(N__13503));
    InMux I__1979 (
            .O(N__13619),
            .I(N__13492));
    InMux I__1978 (
            .O(N__13616),
            .I(N__13492));
    InMux I__1977 (
            .O(N__13613),
            .I(N__13492));
    InMux I__1976 (
            .O(N__13612),
            .I(N__13492));
    InMux I__1975 (
            .O(N__13611),
            .I(N__13492));
    InMux I__1974 (
            .O(N__13610),
            .I(N__13479));
    InMux I__1973 (
            .O(N__13609),
            .I(N__13479));
    InMux I__1972 (
            .O(N__13608),
            .I(N__13479));
    InMux I__1971 (
            .O(N__13607),
            .I(N__13479));
    InMux I__1970 (
            .O(N__13606),
            .I(N__13479));
    InMux I__1969 (
            .O(N__13605),
            .I(N__13479));
    InMux I__1968 (
            .O(N__13604),
            .I(N__13466));
    InMux I__1967 (
            .O(N__13603),
            .I(N__13466));
    InMux I__1966 (
            .O(N__13602),
            .I(N__13466));
    InMux I__1965 (
            .O(N__13601),
            .I(N__13466));
    InMux I__1964 (
            .O(N__13600),
            .I(N__13466));
    InMux I__1963 (
            .O(N__13599),
            .I(N__13466));
    LocalMux I__1962 (
            .O(N__13590),
            .I(N__13463));
    LocalMux I__1961 (
            .O(N__13583),
            .I(N__13454));
    LocalMux I__1960 (
            .O(N__13570),
            .I(N__13454));
    LocalMux I__1959 (
            .O(N__13557),
            .I(N__13454));
    Span4Mux_h I__1958 (
            .O(N__13552),
            .I(N__13454));
    InMux I__1957 (
            .O(N__13551),
            .I(N__13447));
    InMux I__1956 (
            .O(N__13550),
            .I(N__13447));
    InMux I__1955 (
            .O(N__13549),
            .I(N__13447));
    LocalMux I__1954 (
            .O(N__13546),
            .I(N__13444));
    LocalMux I__1953 (
            .O(N__13533),
            .I(N__13439));
    Span4Mux_v I__1952 (
            .O(N__13530),
            .I(N__13439));
    Span4Mux_h I__1951 (
            .O(N__13527),
            .I(N__13436));
    LocalMux I__1950 (
            .O(N__13520),
            .I(N__13415));
    LocalMux I__1949 (
            .O(N__13515),
            .I(N__13415));
    LocalMux I__1948 (
            .O(N__13512),
            .I(N__13415));
    LocalMux I__1947 (
            .O(N__13503),
            .I(N__13415));
    LocalMux I__1946 (
            .O(N__13492),
            .I(N__13415));
    LocalMux I__1945 (
            .O(N__13479),
            .I(N__13415));
    LocalMux I__1944 (
            .O(N__13466),
            .I(N__13415));
    Span4Mux_v I__1943 (
            .O(N__13463),
            .I(N__13415));
    Span4Mux_v I__1942 (
            .O(N__13454),
            .I(N__13415));
    LocalMux I__1941 (
            .O(N__13447),
            .I(N__13415));
    Span4Mux_h I__1940 (
            .O(N__13444),
            .I(N__13412));
    Span4Mux_h I__1939 (
            .O(N__13439),
            .I(N__13407));
    Span4Mux_v I__1938 (
            .O(N__13436),
            .I(N__13407));
    Span4Mux_v I__1937 (
            .O(N__13415),
            .I(N__13404));
    Odrv4 I__1936 (
            .O(N__13412),
            .I(\tok.n29_adj_787 ));
    Odrv4 I__1935 (
            .O(N__13407),
            .I(\tok.n29_adj_787 ));
    Odrv4 I__1934 (
            .O(N__13404),
            .I(\tok.n29_adj_787 ));
    CascadeMux I__1933 (
            .O(N__13397),
            .I(N__13393));
    CascadeMux I__1932 (
            .O(N__13396),
            .I(N__13390));
    InMux I__1931 (
            .O(N__13393),
            .I(N__13387));
    InMux I__1930 (
            .O(N__13390),
            .I(N__13384));
    LocalMux I__1929 (
            .O(N__13387),
            .I(N__13381));
    LocalMux I__1928 (
            .O(N__13384),
            .I(\tok.C_stk.tail_22 ));
    Odrv4 I__1927 (
            .O(N__13381),
            .I(\tok.C_stk.tail_22 ));
    CEMux I__1926 (
            .O(N__13376),
            .I(N__13373));
    LocalMux I__1925 (
            .O(N__13373),
            .I(N__13367));
    CEMux I__1924 (
            .O(N__13372),
            .I(N__13364));
    CEMux I__1923 (
            .O(N__13371),
            .I(N__13357));
    CEMux I__1922 (
            .O(N__13370),
            .I(N__13354));
    Span4Mux_v I__1921 (
            .O(N__13367),
            .I(N__13349));
    LocalMux I__1920 (
            .O(N__13364),
            .I(N__13349));
    CEMux I__1919 (
            .O(N__13363),
            .I(N__13346));
    CEMux I__1918 (
            .O(N__13362),
            .I(N__13342));
    CEMux I__1917 (
            .O(N__13361),
            .I(N__13339));
    CEMux I__1916 (
            .O(N__13360),
            .I(N__13336));
    LocalMux I__1915 (
            .O(N__13357),
            .I(N__13331));
    LocalMux I__1914 (
            .O(N__13354),
            .I(N__13331));
    Span4Mux_v I__1913 (
            .O(N__13349),
            .I(N__13325));
    LocalMux I__1912 (
            .O(N__13346),
            .I(N__13322));
    CEMux I__1911 (
            .O(N__13345),
            .I(N__13319));
    LocalMux I__1910 (
            .O(N__13342),
            .I(N__13316));
    LocalMux I__1909 (
            .O(N__13339),
            .I(N__13313));
    LocalMux I__1908 (
            .O(N__13336),
            .I(N__13310));
    Span4Mux_v I__1907 (
            .O(N__13331),
            .I(N__13307));
    CEMux I__1906 (
            .O(N__13330),
            .I(N__13304));
    CEMux I__1905 (
            .O(N__13329),
            .I(N__13301));
    CEMux I__1904 (
            .O(N__13328),
            .I(N__13298));
    Span4Mux_s2_h I__1903 (
            .O(N__13325),
            .I(N__13295));
    Span4Mux_h I__1902 (
            .O(N__13322),
            .I(N__13290));
    LocalMux I__1901 (
            .O(N__13319),
            .I(N__13290));
    Span4Mux_v I__1900 (
            .O(N__13316),
            .I(N__13285));
    Span4Mux_v I__1899 (
            .O(N__13313),
            .I(N__13285));
    Span4Mux_v I__1898 (
            .O(N__13310),
            .I(N__13276));
    Span4Mux_v I__1897 (
            .O(N__13307),
            .I(N__13276));
    LocalMux I__1896 (
            .O(N__13304),
            .I(N__13276));
    LocalMux I__1895 (
            .O(N__13301),
            .I(N__13276));
    LocalMux I__1894 (
            .O(N__13298),
            .I(N__13273));
    Odrv4 I__1893 (
            .O(N__13295),
            .I(\tok.C_stk_delta_0 ));
    Odrv4 I__1892 (
            .O(N__13290),
            .I(\tok.C_stk_delta_0 ));
    Odrv4 I__1891 (
            .O(N__13285),
            .I(\tok.C_stk_delta_0 ));
    Odrv4 I__1890 (
            .O(N__13276),
            .I(\tok.C_stk_delta_0 ));
    Odrv4 I__1889 (
            .O(N__13273),
            .I(\tok.C_stk_delta_0 ));
    InMux I__1888 (
            .O(N__13262),
            .I(N__13256));
    InMux I__1887 (
            .O(N__13261),
            .I(N__13256));
    LocalMux I__1886 (
            .O(N__13256),
            .I(uart_rx_data_4));
    InMux I__1885 (
            .O(N__13253),
            .I(N__13250));
    LocalMux I__1884 (
            .O(N__13250),
            .I(N__13247));
    Odrv4 I__1883 (
            .O(N__13247),
            .I(\tok.n12_adj_826 ));
    InMux I__1882 (
            .O(N__13244),
            .I(N__13241));
    LocalMux I__1881 (
            .O(N__13241),
            .I(N__13238));
    Span4Mux_h I__1880 (
            .O(N__13238),
            .I(N__13234));
    InMux I__1879 (
            .O(N__13237),
            .I(N__13231));
    Odrv4 I__1878 (
            .O(N__13234),
            .I(\tok.n11_adj_788 ));
    LocalMux I__1877 (
            .O(N__13231),
            .I(\tok.n11_adj_788 ));
    CascadeMux I__1876 (
            .O(N__13226),
            .I(N__13223));
    InMux I__1875 (
            .O(N__13223),
            .I(N__13220));
    LocalMux I__1874 (
            .O(N__13220),
            .I(N__13217));
    Span4Mux_h I__1873 (
            .O(N__13217),
            .I(N__13214));
    Span4Mux_v I__1872 (
            .O(N__13214),
            .I(N__13211));
    Odrv4 I__1871 (
            .O(N__13211),
            .I(sender_2));
    InMux I__1870 (
            .O(N__13208),
            .I(N__13205));
    LocalMux I__1869 (
            .O(N__13205),
            .I(\tok.uart.sender_3 ));
    InMux I__1868 (
            .O(N__13202),
            .I(N__13199));
    LocalMux I__1867 (
            .O(N__13199),
            .I(\tok.uart.sender_4 ));
    InMux I__1866 (
            .O(N__13196),
            .I(N__13193));
    LocalMux I__1865 (
            .O(N__13193),
            .I(\tok.uart.sender_5 ));
    InMux I__1864 (
            .O(N__13190),
            .I(N__13187));
    LocalMux I__1863 (
            .O(N__13187),
            .I(\tok.uart.sender_6 ));
    InMux I__1862 (
            .O(N__13184),
            .I(N__13181));
    LocalMux I__1861 (
            .O(N__13181),
            .I(\tok.uart.sender_7 ));
    InMux I__1860 (
            .O(N__13178),
            .I(N__13175));
    LocalMux I__1859 (
            .O(N__13175),
            .I(N__13172));
    Span4Mux_h I__1858 (
            .O(N__13172),
            .I(N__13169));
    Odrv4 I__1857 (
            .O(N__13169),
            .I(\tok.n5391 ));
    CascadeMux I__1856 (
            .O(N__13166),
            .I(\tok.n14_adj_688_cascade_ ));
    CascadeMux I__1855 (
            .O(N__13163),
            .I(\tok.n2735_cascade_ ));
    CascadeMux I__1854 (
            .O(N__13160),
            .I(\tok.n1_adj_850_cascade_ ));
    InMux I__1853 (
            .O(N__13157),
            .I(N__13154));
    LocalMux I__1852 (
            .O(N__13154),
            .I(\tok.n26_adj_750 ));
    InMux I__1851 (
            .O(N__13151),
            .I(N__13148));
    LocalMux I__1850 (
            .O(N__13148),
            .I(\tok.n5380 ));
    CascadeMux I__1849 (
            .O(N__13145),
            .I(N__13142));
    InMux I__1848 (
            .O(N__13142),
            .I(N__13139));
    LocalMux I__1847 (
            .O(N__13139),
            .I(\tok.n8_adj_805 ));
    InMux I__1846 (
            .O(N__13136),
            .I(N__13133));
    LocalMux I__1845 (
            .O(N__13133),
            .I(N__13130));
    Span4Mux_v I__1844 (
            .O(N__13130),
            .I(N__13125));
    InMux I__1843 (
            .O(N__13129),
            .I(N__13122));
    InMux I__1842 (
            .O(N__13128),
            .I(N__13119));
    Odrv4 I__1841 (
            .O(N__13125),
            .I(\tok.n11_adj_793 ));
    LocalMux I__1840 (
            .O(N__13122),
            .I(\tok.n11_adj_793 ));
    LocalMux I__1839 (
            .O(N__13119),
            .I(\tok.n11_adj_793 ));
    CascadeMux I__1838 (
            .O(N__13112),
            .I(\tok.n5271_cascade_ ));
    InMux I__1837 (
            .O(N__13109),
            .I(N__13106));
    LocalMux I__1836 (
            .O(N__13106),
            .I(\tok.n5318 ));
    InMux I__1835 (
            .O(N__13103),
            .I(N__13100));
    LocalMux I__1834 (
            .O(N__13100),
            .I(\tok.n11_adj_694 ));
    InMux I__1833 (
            .O(N__13097),
            .I(N__13094));
    LocalMux I__1832 (
            .O(N__13094),
            .I(\tok.n15_adj_695 ));
    InMux I__1831 (
            .O(N__13091),
            .I(N__13087));
    CascadeMux I__1830 (
            .O(N__13090),
            .I(N__13083));
    LocalMux I__1829 (
            .O(N__13087),
            .I(N__13080));
    CascadeMux I__1828 (
            .O(N__13086),
            .I(N__13077));
    InMux I__1827 (
            .O(N__13083),
            .I(N__13073));
    Span4Mux_s2_h I__1826 (
            .O(N__13080),
            .I(N__13070));
    InMux I__1825 (
            .O(N__13077),
            .I(N__13065));
    InMux I__1824 (
            .O(N__13076),
            .I(N__13065));
    LocalMux I__1823 (
            .O(N__13073),
            .I(N__13062));
    Odrv4 I__1822 (
            .O(N__13070),
            .I(tc_3));
    LocalMux I__1821 (
            .O(N__13065),
            .I(tc_3));
    Odrv4 I__1820 (
            .O(N__13062),
            .I(tc_3));
    InMux I__1819 (
            .O(N__13055),
            .I(\tok.n4756 ));
    InMux I__1818 (
            .O(N__13052),
            .I(\tok.n4757 ));
    InMux I__1817 (
            .O(N__13049),
            .I(N__13045));
    CascadeMux I__1816 (
            .O(N__13048),
            .I(N__13042));
    LocalMux I__1815 (
            .O(N__13045),
            .I(N__13037));
    InMux I__1814 (
            .O(N__13042),
            .I(N__13032));
    InMux I__1813 (
            .O(N__13041),
            .I(N__13032));
    InMux I__1812 (
            .O(N__13040),
            .I(N__13029));
    Odrv4 I__1811 (
            .O(N__13037),
            .I(tc_5));
    LocalMux I__1810 (
            .O(N__13032),
            .I(tc_5));
    LocalMux I__1809 (
            .O(N__13029),
            .I(tc_5));
    InMux I__1808 (
            .O(N__13022),
            .I(N__13019));
    LocalMux I__1807 (
            .O(N__13019),
            .I(N__13015));
    InMux I__1806 (
            .O(N__13018),
            .I(N__13010));
    Span4Mux_h I__1805 (
            .O(N__13015),
            .I(N__13007));
    InMux I__1804 (
            .O(N__13014),
            .I(N__13002));
    InMux I__1803 (
            .O(N__13013),
            .I(N__13002));
    LocalMux I__1802 (
            .O(N__13010),
            .I(\tok.tc_plus_1_5 ));
    Odrv4 I__1801 (
            .O(N__13007),
            .I(\tok.tc_plus_1_5 ));
    LocalMux I__1800 (
            .O(N__13002),
            .I(\tok.tc_plus_1_5 ));
    InMux I__1799 (
            .O(N__12995),
            .I(\tok.n4758 ));
    InMux I__1798 (
            .O(N__12992),
            .I(\tok.n4759 ));
    InMux I__1797 (
            .O(N__12989),
            .I(N__12984));
    InMux I__1796 (
            .O(N__12988),
            .I(N__12978));
    InMux I__1795 (
            .O(N__12987),
            .I(N__12978));
    LocalMux I__1794 (
            .O(N__12984),
            .I(N__12975));
    InMux I__1793 (
            .O(N__12983),
            .I(N__12972));
    LocalMux I__1792 (
            .O(N__12978),
            .I(N__12967));
    Span4Mux_h I__1791 (
            .O(N__12975),
            .I(N__12967));
    LocalMux I__1790 (
            .O(N__12972),
            .I(tc_7));
    Odrv4 I__1789 (
            .O(N__12967),
            .I(tc_7));
    InMux I__1788 (
            .O(N__12962),
            .I(\tok.n4760 ));
    InMux I__1787 (
            .O(N__12959),
            .I(N__12954));
    InMux I__1786 (
            .O(N__12958),
            .I(N__12949));
    InMux I__1785 (
            .O(N__12957),
            .I(N__12949));
    LocalMux I__1784 (
            .O(N__12954),
            .I(N__12943));
    LocalMux I__1783 (
            .O(N__12949),
            .I(N__12943));
    InMux I__1782 (
            .O(N__12948),
            .I(N__12940));
    Span4Mux_h I__1781 (
            .O(N__12943),
            .I(N__12937));
    LocalMux I__1780 (
            .O(N__12940),
            .I(\tok.tc_plus_1_7 ));
    Odrv4 I__1779 (
            .O(N__12937),
            .I(\tok.tc_plus_1_7 ));
    CascadeMux I__1778 (
            .O(N__12932),
            .I(N__12929));
    InMux I__1777 (
            .O(N__12929),
            .I(N__12920));
    InMux I__1776 (
            .O(N__12928),
            .I(N__12907));
    InMux I__1775 (
            .O(N__12927),
            .I(N__12907));
    InMux I__1774 (
            .O(N__12926),
            .I(N__12907));
    InMux I__1773 (
            .O(N__12925),
            .I(N__12907));
    InMux I__1772 (
            .O(N__12924),
            .I(N__12907));
    InMux I__1771 (
            .O(N__12923),
            .I(N__12907));
    LocalMux I__1770 (
            .O(N__12920),
            .I(N__12904));
    LocalMux I__1769 (
            .O(N__12907),
            .I(N__12901));
    Span4Mux_v I__1768 (
            .O(N__12904),
            .I(N__12898));
    Odrv12 I__1767 (
            .O(N__12901),
            .I(\tok.n9_adj_798 ));
    Odrv4 I__1766 (
            .O(N__12898),
            .I(\tok.n9_adj_798 ));
    InMux I__1765 (
            .O(N__12893),
            .I(N__12890));
    LocalMux I__1764 (
            .O(N__12890),
            .I(\tok.n5293 ));
    InMux I__1763 (
            .O(N__12887),
            .I(N__12881));
    InMux I__1762 (
            .O(N__12886),
            .I(N__12881));
    LocalMux I__1761 (
            .O(N__12881),
            .I(N__12878));
    Span4Mux_v I__1760 (
            .O(N__12878),
            .I(N__12875));
    Odrv4 I__1759 (
            .O(N__12875),
            .I(\tok.key_rd_7 ));
    InMux I__1758 (
            .O(N__12872),
            .I(N__12866));
    InMux I__1757 (
            .O(N__12871),
            .I(N__12866));
    LocalMux I__1756 (
            .O(N__12866),
            .I(N__12863));
    Span4Mux_h I__1755 (
            .O(N__12863),
            .I(N__12860));
    Odrv4 I__1754 (
            .O(N__12860),
            .I(\tok.key_rd_2 ));
    InMux I__1753 (
            .O(N__12857),
            .I(N__12854));
    LocalMux I__1752 (
            .O(N__12854),
            .I(\tok.n22_adj_721 ));
    InMux I__1751 (
            .O(N__12851),
            .I(N__12848));
    LocalMux I__1750 (
            .O(N__12848),
            .I(\tok.n23_adj_731 ));
    InMux I__1749 (
            .O(N__12845),
            .I(N__12842));
    LocalMux I__1748 (
            .O(N__12842),
            .I(\tok.n24_adj_651 ));
    InMux I__1747 (
            .O(N__12839),
            .I(N__12833));
    InMux I__1746 (
            .O(N__12838),
            .I(N__12833));
    LocalMux I__1745 (
            .O(N__12833),
            .I(N__12830));
    Odrv4 I__1744 (
            .O(N__12830),
            .I(\tok.key_rd_14 ));
    InMux I__1743 (
            .O(N__12827),
            .I(N__12821));
    InMux I__1742 (
            .O(N__12826),
            .I(N__12821));
    LocalMux I__1741 (
            .O(N__12821),
            .I(N__12818));
    Span4Mux_h I__1740 (
            .O(N__12818),
            .I(N__12815));
    Odrv4 I__1739 (
            .O(N__12815),
            .I(\tok.key_rd_15 ));
    CascadeMux I__1738 (
            .O(N__12812),
            .I(N__12809));
    InMux I__1737 (
            .O(N__12809),
            .I(N__12803));
    InMux I__1736 (
            .O(N__12808),
            .I(N__12803));
    LocalMux I__1735 (
            .O(N__12803),
            .I(N__12800));
    Odrv4 I__1734 (
            .O(N__12800),
            .I(\tok.key_rd_9 ));
    InMux I__1733 (
            .O(N__12797),
            .I(N__12791));
    InMux I__1732 (
            .O(N__12796),
            .I(N__12791));
    LocalMux I__1731 (
            .O(N__12791),
            .I(N__12788));
    Odrv4 I__1730 (
            .O(N__12788),
            .I(\tok.key_rd_11 ));
    InMux I__1729 (
            .O(N__12785),
            .I(N__12781));
    InMux I__1728 (
            .O(N__12784),
            .I(N__12776));
    LocalMux I__1727 (
            .O(N__12781),
            .I(N__12773));
    InMux I__1726 (
            .O(N__12780),
            .I(N__12768));
    InMux I__1725 (
            .O(N__12779),
            .I(N__12768));
    LocalMux I__1724 (
            .O(N__12776),
            .I(N__12765));
    Odrv4 I__1723 (
            .O(N__12773),
            .I(tc_0));
    LocalMux I__1722 (
            .O(N__12768),
            .I(tc_0));
    Odrv4 I__1721 (
            .O(N__12765),
            .I(tc_0));
    InMux I__1720 (
            .O(N__12758),
            .I(N__12753));
    InMux I__1719 (
            .O(N__12757),
            .I(N__12749));
    CascadeMux I__1718 (
            .O(N__12756),
            .I(N__12746));
    LocalMux I__1717 (
            .O(N__12753),
            .I(N__12743));
    InMux I__1716 (
            .O(N__12752),
            .I(N__12740));
    LocalMux I__1715 (
            .O(N__12749),
            .I(N__12737));
    InMux I__1714 (
            .O(N__12746),
            .I(N__12734));
    Span12Mux_s1_h I__1713 (
            .O(N__12743),
            .I(N__12729));
    LocalMux I__1712 (
            .O(N__12740),
            .I(N__12729));
    Span4Mux_h I__1711 (
            .O(N__12737),
            .I(N__12726));
    LocalMux I__1710 (
            .O(N__12734),
            .I(\tok.tc_plus_1_0 ));
    Odrv12 I__1709 (
            .O(N__12729),
            .I(\tok.tc_plus_1_0 ));
    Odrv4 I__1708 (
            .O(N__12726),
            .I(\tok.tc_plus_1_0 ));
    InMux I__1707 (
            .O(N__12719),
            .I(bfn_5_8_0_));
    InMux I__1706 (
            .O(N__12716),
            .I(N__12713));
    LocalMux I__1705 (
            .O(N__12713),
            .I(N__12707));
    InMux I__1704 (
            .O(N__12712),
            .I(N__12702));
    InMux I__1703 (
            .O(N__12711),
            .I(N__12702));
    InMux I__1702 (
            .O(N__12710),
            .I(N__12699));
    Span4Mux_h I__1701 (
            .O(N__12707),
            .I(N__12696));
    LocalMux I__1700 (
            .O(N__12702),
            .I(N__12693));
    LocalMux I__1699 (
            .O(N__12699),
            .I(\tok.tc_plus_1_1 ));
    Odrv4 I__1698 (
            .O(N__12696),
            .I(\tok.tc_plus_1_1 ));
    Odrv4 I__1697 (
            .O(N__12693),
            .I(\tok.tc_plus_1_1 ));
    InMux I__1696 (
            .O(N__12686),
            .I(\tok.n4754 ));
    InMux I__1695 (
            .O(N__12683),
            .I(N__12677));
    InMux I__1694 (
            .O(N__12682),
            .I(N__12674));
    InMux I__1693 (
            .O(N__12681),
            .I(N__12669));
    InMux I__1692 (
            .O(N__12680),
            .I(N__12669));
    LocalMux I__1691 (
            .O(N__12677),
            .I(N__12666));
    LocalMux I__1690 (
            .O(N__12674),
            .I(tc_2));
    LocalMux I__1689 (
            .O(N__12669),
            .I(tc_2));
    Odrv12 I__1688 (
            .O(N__12666),
            .I(tc_2));
    InMux I__1687 (
            .O(N__12659),
            .I(N__12655));
    InMux I__1686 (
            .O(N__12658),
            .I(N__12651));
    LocalMux I__1685 (
            .O(N__12655),
            .I(N__12647));
    InMux I__1684 (
            .O(N__12654),
            .I(N__12644));
    LocalMux I__1683 (
            .O(N__12651),
            .I(N__12641));
    InMux I__1682 (
            .O(N__12650),
            .I(N__12638));
    Span4Mux_v I__1681 (
            .O(N__12647),
            .I(N__12633));
    LocalMux I__1680 (
            .O(N__12644),
            .I(N__12633));
    Span4Mux_h I__1679 (
            .O(N__12641),
            .I(N__12630));
    LocalMux I__1678 (
            .O(N__12638),
            .I(\tok.tc_plus_1_2 ));
    Odrv4 I__1677 (
            .O(N__12633),
            .I(\tok.tc_plus_1_2 ));
    Odrv4 I__1676 (
            .O(N__12630),
            .I(\tok.tc_plus_1_2 ));
    InMux I__1675 (
            .O(N__12623),
            .I(\tok.n4755 ));
    CascadeMux I__1674 (
            .O(N__12620),
            .I(\tok.n83_adj_848_cascade_ ));
    CascadeMux I__1673 (
            .O(N__12617),
            .I(N__12613));
    InMux I__1672 (
            .O(N__12616),
            .I(N__12606));
    InMux I__1671 (
            .O(N__12613),
            .I(N__12606));
    InMux I__1670 (
            .O(N__12612),
            .I(N__12603));
    InMux I__1669 (
            .O(N__12611),
            .I(N__12600));
    LocalMux I__1668 (
            .O(N__12606),
            .I(N__12595));
    LocalMux I__1667 (
            .O(N__12603),
            .I(N__12595));
    LocalMux I__1666 (
            .O(N__12600),
            .I(\tok.c_stk_r_1 ));
    Odrv12 I__1665 (
            .O(N__12595),
            .I(\tok.c_stk_r_1 ));
    CascadeMux I__1664 (
            .O(N__12590),
            .I(\tok.ram.n5594_cascade_ ));
    InMux I__1663 (
            .O(N__12587),
            .I(N__12584));
    LocalMux I__1662 (
            .O(N__12584),
            .I(\tok.n5610 ));
    CascadeMux I__1661 (
            .O(N__12581),
            .I(\tok.n3_cascade_ ));
    CascadeMux I__1660 (
            .O(N__12578),
            .I(\tok.n13_cascade_ ));
    InMux I__1659 (
            .O(N__12575),
            .I(N__12572));
    LocalMux I__1658 (
            .O(N__12572),
            .I(N__12569));
    Span4Mux_h I__1657 (
            .O(N__12569),
            .I(N__12566));
    Span4Mux_s3_h I__1656 (
            .O(N__12566),
            .I(N__12563));
    Odrv4 I__1655 (
            .O(N__12563),
            .I(\tok.uart.n5 ));
    InMux I__1654 (
            .O(N__12560),
            .I(N__12554));
    InMux I__1653 (
            .O(N__12559),
            .I(N__12554));
    LocalMux I__1652 (
            .O(N__12554),
            .I(N__12551));
    Odrv4 I__1651 (
            .O(N__12551),
            .I(\tok.key_rd_10 ));
    CascadeMux I__1650 (
            .O(N__12548),
            .I(N__12545));
    InMux I__1649 (
            .O(N__12545),
            .I(N__12539));
    InMux I__1648 (
            .O(N__12544),
            .I(N__12539));
    LocalMux I__1647 (
            .O(N__12539),
            .I(N__12536));
    Odrv4 I__1646 (
            .O(N__12536),
            .I(\tok.key_rd_12 ));
    CascadeMux I__1645 (
            .O(N__12533),
            .I(\tok.n21_adj_733_cascade_ ));
    CascadeMux I__1644 (
            .O(N__12530),
            .I(\tok.n13_adj_691_cascade_ ));
    CascadeMux I__1643 (
            .O(N__12527),
            .I(n10_adj_871_cascade_));
    CascadeMux I__1642 (
            .O(N__12524),
            .I(N__12521));
    InMux I__1641 (
            .O(N__12521),
            .I(N__12518));
    LocalMux I__1640 (
            .O(N__12518),
            .I(N__12515));
    Span4Mux_h I__1639 (
            .O(N__12515),
            .I(N__12512));
    Sp12to4 I__1638 (
            .O(N__12512),
            .I(N__12509));
    Odrv12 I__1637 (
            .O(N__12509),
            .I(\tok.tc_6 ));
    CascadeMux I__1636 (
            .O(N__12506),
            .I(\tok.ram.n5605_cascade_ ));
    InMux I__1635 (
            .O(N__12503),
            .I(N__12500));
    LocalMux I__1634 (
            .O(N__12500),
            .I(\tok.n3_adj_690 ));
    CascadeMux I__1633 (
            .O(N__12497),
            .I(\tok.n83_adj_687_cascade_ ));
    CascadeMux I__1632 (
            .O(N__12494),
            .I(N__12491));
    InMux I__1631 (
            .O(N__12491),
            .I(N__12488));
    LocalMux I__1630 (
            .O(N__12488),
            .I(\tok.n5505 ));
    InMux I__1629 (
            .O(N__12485),
            .I(N__12482));
    LocalMux I__1628 (
            .O(N__12482),
            .I(n10_adj_871));
    InMux I__1627 (
            .O(N__12479),
            .I(N__12476));
    LocalMux I__1626 (
            .O(N__12476),
            .I(\tok.n27_adj_825 ));
    CascadeMux I__1625 (
            .O(N__12473),
            .I(\tok.n5285_cascade_ ));
    CascadeMux I__1624 (
            .O(N__12470),
            .I(\tok.n1_adj_715_cascade_ ));
    InMux I__1623 (
            .O(N__12467),
            .I(N__12455));
    InMux I__1622 (
            .O(N__12466),
            .I(N__12455));
    InMux I__1621 (
            .O(N__12465),
            .I(N__12455));
    InMux I__1620 (
            .O(N__12464),
            .I(N__12455));
    LocalMux I__1619 (
            .O(N__12455),
            .I(\tok.n190 ));
    InMux I__1618 (
            .O(N__12452),
            .I(N__12447));
    InMux I__1617 (
            .O(N__12451),
            .I(N__12441));
    InMux I__1616 (
            .O(N__12450),
            .I(N__12441));
    LocalMux I__1615 (
            .O(N__12447),
            .I(N__12438));
    InMux I__1614 (
            .O(N__12446),
            .I(N__12435));
    LocalMux I__1613 (
            .O(N__12441),
            .I(N__12432));
    Odrv4 I__1612 (
            .O(N__12438),
            .I(\tok.n890 ));
    LocalMux I__1611 (
            .O(N__12435),
            .I(\tok.n890 ));
    Odrv4 I__1610 (
            .O(N__12432),
            .I(\tok.n890 ));
    CascadeMux I__1609 (
            .O(N__12425),
            .I(\tok.n10_adj_763_cascade_ ));
    InMux I__1608 (
            .O(N__12422),
            .I(N__12416));
    CascadeMux I__1607 (
            .O(N__12421),
            .I(N__12412));
    InMux I__1606 (
            .O(N__12420),
            .I(N__12409));
    InMux I__1605 (
            .O(N__12419),
            .I(N__12406));
    LocalMux I__1604 (
            .O(N__12416),
            .I(N__12403));
    InMux I__1603 (
            .O(N__12415),
            .I(N__12398));
    InMux I__1602 (
            .O(N__12412),
            .I(N__12398));
    LocalMux I__1601 (
            .O(N__12409),
            .I(\tok.n5338 ));
    LocalMux I__1600 (
            .O(N__12406),
            .I(\tok.n5338 ));
    Odrv4 I__1599 (
            .O(N__12403),
            .I(\tok.n5338 ));
    LocalMux I__1598 (
            .O(N__12398),
            .I(\tok.n5338 ));
    InMux I__1597 (
            .O(N__12389),
            .I(N__12383));
    InMux I__1596 (
            .O(N__12388),
            .I(N__12383));
    LocalMux I__1595 (
            .O(N__12383),
            .I(\tok.n5340 ));
    CascadeMux I__1594 (
            .O(N__12380),
            .I(N__12374));
    InMux I__1593 (
            .O(N__12379),
            .I(N__12371));
    InMux I__1592 (
            .O(N__12378),
            .I(N__12364));
    InMux I__1591 (
            .O(N__12377),
            .I(N__12364));
    InMux I__1590 (
            .O(N__12374),
            .I(N__12364));
    LocalMux I__1589 (
            .O(N__12371),
            .I(\tok.A_stk_delta_1__N_4 ));
    LocalMux I__1588 (
            .O(N__12364),
            .I(\tok.A_stk_delta_1__N_4 ));
    InMux I__1587 (
            .O(N__12359),
            .I(N__12348));
    InMux I__1586 (
            .O(N__12358),
            .I(N__12348));
    InMux I__1585 (
            .O(N__12357),
            .I(N__12345));
    InMux I__1584 (
            .O(N__12356),
            .I(N__12336));
    InMux I__1583 (
            .O(N__12355),
            .I(N__12336));
    InMux I__1582 (
            .O(N__12354),
            .I(N__12336));
    InMux I__1581 (
            .O(N__12353),
            .I(N__12336));
    LocalMux I__1580 (
            .O(N__12348),
            .I(\tok.n61 ));
    LocalMux I__1579 (
            .O(N__12345),
            .I(\tok.n61 ));
    LocalMux I__1578 (
            .O(N__12336),
            .I(\tok.n61 ));
    InMux I__1577 (
            .O(N__12329),
            .I(N__12317));
    InMux I__1576 (
            .O(N__12328),
            .I(N__12317));
    InMux I__1575 (
            .O(N__12327),
            .I(N__12317));
    InMux I__1574 (
            .O(N__12326),
            .I(N__12317));
    LocalMux I__1573 (
            .O(N__12317),
            .I(\tok.n4_adj_813 ));
    InMux I__1572 (
            .O(N__12314),
            .I(N__12310));
    InMux I__1571 (
            .O(N__12313),
            .I(N__12307));
    LocalMux I__1570 (
            .O(N__12310),
            .I(tail_97));
    LocalMux I__1569 (
            .O(N__12307),
            .I(tail_97));
    InMux I__1568 (
            .O(N__12302),
            .I(N__12299));
    LocalMux I__1567 (
            .O(N__12299),
            .I(N__12295));
    InMux I__1566 (
            .O(N__12298),
            .I(N__12292));
    Odrv12 I__1565 (
            .O(N__12295),
            .I(tail_113));
    LocalMux I__1564 (
            .O(N__12292),
            .I(tail_113));
    CascadeMux I__1563 (
            .O(N__12287),
            .I(\tok.n27_adj_828_cascade_ ));
    CascadeMux I__1562 (
            .O(N__12284),
            .I(\tok.n27_adj_831_cascade_ ));
    CascadeMux I__1561 (
            .O(N__12281),
            .I(\tok.n27_adj_833_cascade_ ));
    InMux I__1560 (
            .O(N__12278),
            .I(N__12275));
    LocalMux I__1559 (
            .O(N__12275),
            .I(N__12272));
    Odrv12 I__1558 (
            .O(N__12272),
            .I(\tok.n7_adj_785 ));
    CascadeMux I__1557 (
            .O(N__12269),
            .I(\tok.n14_adj_644_cascade_ ));
    InMux I__1556 (
            .O(N__12266),
            .I(N__12263));
    LocalMux I__1555 (
            .O(N__12263),
            .I(N__12260));
    Odrv4 I__1554 (
            .O(N__12260),
            .I(\tok.table_wr_data_11 ));
    InMux I__1553 (
            .O(N__12257),
            .I(N__12254));
    LocalMux I__1552 (
            .O(N__12254),
            .I(\tok.table_wr_data_10 ));
    InMux I__1551 (
            .O(N__12251),
            .I(N__12248));
    LocalMux I__1550 (
            .O(N__12248),
            .I(\tok.table_wr_data_9 ));
    InMux I__1549 (
            .O(N__12245),
            .I(N__12242));
    LocalMux I__1548 (
            .O(N__12242),
            .I(\tok.table_wr_data_8 ));
    InMux I__1547 (
            .O(N__12239),
            .I(N__12236));
    LocalMux I__1546 (
            .O(N__12236),
            .I(\tok.table_wr_data_0 ));
    InMux I__1545 (
            .O(N__12233),
            .I(N__12230));
    LocalMux I__1544 (
            .O(N__12230),
            .I(N__12227));
    Odrv12 I__1543 (
            .O(N__12227),
            .I(\tok.n8_adj_790 ));
    InMux I__1542 (
            .O(N__12224),
            .I(N__12221));
    LocalMux I__1541 (
            .O(N__12221),
            .I(N__12218));
    Span12Mux_s4_h I__1540 (
            .O(N__12218),
            .I(N__12215));
    Odrv12 I__1539 (
            .O(N__12215),
            .I(\tok.table_wr_data_15 ));
    InMux I__1538 (
            .O(N__12212),
            .I(N__12209));
    LocalMux I__1537 (
            .O(N__12209),
            .I(\tok.table_wr_data_14 ));
    InMux I__1536 (
            .O(N__12206),
            .I(N__12203));
    LocalMux I__1535 (
            .O(N__12203),
            .I(N__12200));
    Span4Mux_v I__1534 (
            .O(N__12200),
            .I(N__12197));
    Odrv4 I__1533 (
            .O(N__12197),
            .I(\tok.table_wr_data_3 ));
    InMux I__1532 (
            .O(N__12194),
            .I(N__12191));
    LocalMux I__1531 (
            .O(N__12191),
            .I(N__12188));
    Span4Mux_v I__1530 (
            .O(N__12188),
            .I(N__12185));
    Span4Mux_h I__1529 (
            .O(N__12185),
            .I(N__12182));
    Odrv4 I__1528 (
            .O(N__12182),
            .I(\tok.table_wr_data_2 ));
    InMux I__1527 (
            .O(N__12179),
            .I(N__12176));
    LocalMux I__1526 (
            .O(N__12176),
            .I(N__12173));
    Odrv4 I__1525 (
            .O(N__12173),
            .I(\tok.table_wr_data_1 ));
    InMux I__1524 (
            .O(N__12170),
            .I(N__12167));
    LocalMux I__1523 (
            .O(N__12167),
            .I(N__12164));
    Odrv4 I__1522 (
            .O(N__12164),
            .I(\tok.table_wr_data_5 ));
    InMux I__1521 (
            .O(N__12161),
            .I(N__12158));
    LocalMux I__1520 (
            .O(N__12158),
            .I(N__12155));
    Odrv4 I__1519 (
            .O(N__12155),
            .I(\tok.table_wr_data_7 ));
    InMux I__1518 (
            .O(N__12152),
            .I(N__12149));
    LocalMux I__1517 (
            .O(N__12149),
            .I(N__12146));
    Odrv4 I__1516 (
            .O(N__12146),
            .I(\tok.table_wr_data_13 ));
    InMux I__1515 (
            .O(N__12143),
            .I(N__12140));
    LocalMux I__1514 (
            .O(N__12140),
            .I(\tok.table_wr_data_12 ));
    CascadeMux I__1513 (
            .O(N__12137),
            .I(\tok.ram.n5608_cascade_ ));
    CascadeMux I__1512 (
            .O(N__12134),
            .I(N__12129));
    InMux I__1511 (
            .O(N__12133),
            .I(N__12121));
    InMux I__1510 (
            .O(N__12132),
            .I(N__12121));
    InMux I__1509 (
            .O(N__12129),
            .I(N__12121));
    CascadeMux I__1508 (
            .O(N__12128),
            .I(N__12118));
    LocalMux I__1507 (
            .O(N__12121),
            .I(N__12115));
    InMux I__1506 (
            .O(N__12118),
            .I(N__12112));
    Span4Mux_h I__1505 (
            .O(N__12115),
            .I(N__12109));
    LocalMux I__1504 (
            .O(N__12112),
            .I(\tok.c_stk_r_5 ));
    Odrv4 I__1503 (
            .O(N__12109),
            .I(\tok.c_stk_r_5 ));
    CascadeMux I__1502 (
            .O(N__12104),
            .I(\tok.n83_adj_678_cascade_ ));
    InMux I__1501 (
            .O(N__12101),
            .I(N__12098));
    LocalMux I__1500 (
            .O(N__12098),
            .I(\tok.n3_adj_683 ));
    CascadeMux I__1499 (
            .O(N__12095),
            .I(\tok.n5483_cascade_ ));
    CascadeMux I__1498 (
            .O(N__12092),
            .I(\tok.n5_adj_684_cascade_ ));
    CascadeMux I__1497 (
            .O(N__12089),
            .I(n92_adj_868_cascade_));
    CascadeMux I__1496 (
            .O(N__12086),
            .I(N__12083));
    InMux I__1495 (
            .O(N__12083),
            .I(N__12080));
    LocalMux I__1494 (
            .O(N__12080),
            .I(N__12077));
    Span4Mux_v I__1493 (
            .O(N__12077),
            .I(N__12074));
    Odrv4 I__1492 (
            .O(N__12074),
            .I(\tok.tc_5 ));
    InMux I__1491 (
            .O(N__12071),
            .I(N__12068));
    LocalMux I__1490 (
            .O(N__12068),
            .I(n92_adj_868));
    InMux I__1489 (
            .O(N__12065),
            .I(N__12062));
    LocalMux I__1488 (
            .O(N__12062),
            .I(N__12059));
    Odrv4 I__1487 (
            .O(N__12059),
            .I(\tok.table_wr_data_4 ));
    CascadeMux I__1486 (
            .O(N__12056),
            .I(N__12052));
    CascadeMux I__1485 (
            .O(N__12055),
            .I(N__12049));
    InMux I__1484 (
            .O(N__12052),
            .I(N__12041));
    InMux I__1483 (
            .O(N__12049),
            .I(N__12041));
    InMux I__1482 (
            .O(N__12048),
            .I(N__12041));
    LocalMux I__1481 (
            .O(N__12041),
            .I(N__12036));
    InMux I__1480 (
            .O(N__12040),
            .I(N__12031));
    InMux I__1479 (
            .O(N__12039),
            .I(N__12031));
    Span4Mux_h I__1478 (
            .O(N__12036),
            .I(N__12028));
    LocalMux I__1477 (
            .O(N__12031),
            .I(\tok.uart.sentbits_0 ));
    Odrv4 I__1476 (
            .O(N__12028),
            .I(\tok.uart.sentbits_0 ));
    InMux I__1475 (
            .O(N__12023),
            .I(N__12014));
    InMux I__1474 (
            .O(N__12022),
            .I(N__12014));
    InMux I__1473 (
            .O(N__12021),
            .I(N__12014));
    LocalMux I__1472 (
            .O(N__12014),
            .I(N__12010));
    InMux I__1471 (
            .O(N__12013),
            .I(N__12007));
    Span4Mux_h I__1470 (
            .O(N__12010),
            .I(N__12004));
    LocalMux I__1469 (
            .O(N__12007),
            .I(\tok.uart.sentbits_1 ));
    Odrv4 I__1468 (
            .O(N__12004),
            .I(\tok.uart.sentbits_1 ));
    CEMux I__1467 (
            .O(N__11999),
            .I(N__11996));
    LocalMux I__1466 (
            .O(N__11996),
            .I(N__11992));
    CEMux I__1465 (
            .O(N__11995),
            .I(N__11989));
    Span4Mux_v I__1464 (
            .O(N__11992),
            .I(N__11984));
    LocalMux I__1463 (
            .O(N__11989),
            .I(N__11984));
    Odrv4 I__1462 (
            .O(N__11984),
            .I(\tok.uart.n1023 ));
    SRMux I__1461 (
            .O(N__11981),
            .I(N__11977));
    SRMux I__1460 (
            .O(N__11980),
            .I(N__11974));
    LocalMux I__1459 (
            .O(N__11977),
            .I(N__11971));
    LocalMux I__1458 (
            .O(N__11974),
            .I(N__11968));
    Span4Mux_h I__1457 (
            .O(N__11971),
            .I(N__11965));
    Span4Mux_h I__1456 (
            .O(N__11968),
            .I(N__11962));
    Odrv4 I__1455 (
            .O(N__11965),
            .I(\tok.uart.n1093 ));
    Odrv4 I__1454 (
            .O(N__11962),
            .I(\tok.uart.n1093 ));
    CascadeMux I__1453 (
            .O(N__11957),
            .I(N__11954));
    InMux I__1452 (
            .O(N__11954),
            .I(N__11951));
    LocalMux I__1451 (
            .O(N__11951),
            .I(N__11948));
    Span4Mux_v I__1450 (
            .O(N__11948),
            .I(N__11945));
    Odrv4 I__1449 (
            .O(N__11945),
            .I(\tok.n4_adj_707 ));
    InMux I__1448 (
            .O(N__11942),
            .I(N__11939));
    LocalMux I__1447 (
            .O(N__11939),
            .I(N__11936));
    Span4Mux_h I__1446 (
            .O(N__11936),
            .I(N__11933));
    Odrv4 I__1445 (
            .O(N__11933),
            .I(\tok.n42 ));
    InMux I__1444 (
            .O(N__11930),
            .I(N__11927));
    LocalMux I__1443 (
            .O(N__11927),
            .I(\tok.n5287 ));
    CascadeMux I__1442 (
            .O(N__11924),
            .I(\tok.n5287_cascade_ ));
    InMux I__1441 (
            .O(N__11921),
            .I(N__11918));
    LocalMux I__1440 (
            .O(N__11918),
            .I(N__11915));
    Span4Mux_h I__1439 (
            .O(N__11915),
            .I(N__11912));
    Odrv4 I__1438 (
            .O(N__11912),
            .I(\tok.n7 ));
    CascadeMux I__1437 (
            .O(N__11909),
            .I(\tok.n5312_cascade_ ));
    CascadeMux I__1436 (
            .O(N__11906),
            .I(\tok.n15_adj_817_cascade_ ));
    InMux I__1435 (
            .O(N__11903),
            .I(N__11900));
    LocalMux I__1434 (
            .O(N__11900),
            .I(\tok.n898 ));
    CascadeMux I__1433 (
            .O(N__11897),
            .I(\tok.n898_cascade_ ));
    InMux I__1432 (
            .O(N__11894),
            .I(N__11891));
    LocalMux I__1431 (
            .O(N__11891),
            .I(\tok.uart.n6 ));
    CascadeMux I__1430 (
            .O(N__11888),
            .I(N__11883));
    InMux I__1429 (
            .O(N__11887),
            .I(N__11876));
    InMux I__1428 (
            .O(N__11886),
            .I(N__11876));
    InMux I__1427 (
            .O(N__11883),
            .I(N__11871));
    InMux I__1426 (
            .O(N__11882),
            .I(N__11871));
    InMux I__1425 (
            .O(N__11881),
            .I(N__11868));
    LocalMux I__1424 (
            .O(N__11876),
            .I(\tok.n59 ));
    LocalMux I__1423 (
            .O(N__11871),
            .I(\tok.n59 ));
    LocalMux I__1422 (
            .O(N__11868),
            .I(\tok.n59 ));
    InMux I__1421 (
            .O(N__11861),
            .I(N__11858));
    LocalMux I__1420 (
            .O(N__11858),
            .I(\tok.depth_3 ));
    CascadeMux I__1419 (
            .O(N__11855),
            .I(N__11850));
    CascadeMux I__1418 (
            .O(N__11854),
            .I(N__11847));
    InMux I__1417 (
            .O(N__11853),
            .I(N__11830));
    InMux I__1416 (
            .O(N__11850),
            .I(N__11830));
    InMux I__1415 (
            .O(N__11847),
            .I(N__11830));
    InMux I__1414 (
            .O(N__11846),
            .I(N__11830));
    InMux I__1413 (
            .O(N__11845),
            .I(N__11830));
    InMux I__1412 (
            .O(N__11844),
            .I(N__11830));
    InMux I__1411 (
            .O(N__11843),
            .I(N__11827));
    LocalMux I__1410 (
            .O(N__11830),
            .I(\tok.n60 ));
    LocalMux I__1409 (
            .O(N__11827),
            .I(\tok.n60 ));
    InMux I__1408 (
            .O(N__11822),
            .I(N__11819));
    LocalMux I__1407 (
            .O(N__11819),
            .I(\tok.depth_2 ));
    CascadeMux I__1406 (
            .O(N__11816),
            .I(N__11813));
    InMux I__1405 (
            .O(N__11813),
            .I(N__11810));
    LocalMux I__1404 (
            .O(N__11810),
            .I(N__11807));
    Odrv4 I__1403 (
            .O(N__11807),
            .I(\tok.n807 ));
    CascadeMux I__1402 (
            .O(N__11804),
            .I(n23_cascade_));
    InMux I__1401 (
            .O(N__11801),
            .I(N__11795));
    InMux I__1400 (
            .O(N__11800),
            .I(N__11795));
    LocalMux I__1399 (
            .O(N__11795),
            .I(N__11788));
    SRMux I__1398 (
            .O(N__11794),
            .I(N__11785));
    SRMux I__1397 (
            .O(N__11793),
            .I(N__11782));
    InMux I__1396 (
            .O(N__11792),
            .I(N__11777));
    InMux I__1395 (
            .O(N__11791),
            .I(N__11777));
    Span4Mux_v I__1394 (
            .O(N__11788),
            .I(N__11774));
    LocalMux I__1393 (
            .O(N__11785),
            .I(txtick));
    LocalMux I__1392 (
            .O(N__11782),
            .I(txtick));
    LocalMux I__1391 (
            .O(N__11777),
            .I(txtick));
    Odrv4 I__1390 (
            .O(N__11774),
            .I(txtick));
    CascadeMux I__1389 (
            .O(N__11765),
            .I(\tok.A_stk_delta_1__N_4_cascade_ ));
    CascadeMux I__1388 (
            .O(N__11762),
            .I(\tok.depth_1_cascade_ ));
    InMux I__1387 (
            .O(N__11759),
            .I(N__11756));
    LocalMux I__1386 (
            .O(N__11756),
            .I(N__11753));
    Span4Mux_h I__1385 (
            .O(N__11753),
            .I(N__11750));
    Odrv4 I__1384 (
            .O(N__11750),
            .I(\tok.n37 ));
    CascadeMux I__1383 (
            .O(N__11747),
            .I(\tok.n2585_cascade_ ));
    InMux I__1382 (
            .O(N__11744),
            .I(N__11738));
    InMux I__1381 (
            .O(N__11743),
            .I(N__11738));
    LocalMux I__1380 (
            .O(N__11738),
            .I(\tok.A_stk.tail_33 ));
    InMux I__1379 (
            .O(N__11735),
            .I(N__11729));
    InMux I__1378 (
            .O(N__11734),
            .I(N__11729));
    LocalMux I__1377 (
            .O(N__11729),
            .I(\tok.A_stk.tail_49 ));
    InMux I__1376 (
            .O(N__11726),
            .I(N__11720));
    InMux I__1375 (
            .O(N__11725),
            .I(N__11720));
    LocalMux I__1374 (
            .O(N__11720),
            .I(\tok.A_stk.tail_65 ));
    InMux I__1373 (
            .O(N__11717),
            .I(N__11711));
    InMux I__1372 (
            .O(N__11716),
            .I(N__11711));
    LocalMux I__1371 (
            .O(N__11711),
            .I(\tok.A_stk.tail_81 ));
    InMux I__1370 (
            .O(N__11708),
            .I(N__11702));
    InMux I__1369 (
            .O(N__11707),
            .I(N__11702));
    LocalMux I__1368 (
            .O(N__11702),
            .I(\tok.A_stk.tail_1 ));
    CascadeMux I__1367 (
            .O(N__11699),
            .I(N__11696));
    InMux I__1366 (
            .O(N__11696),
            .I(N__11693));
    LocalMux I__1365 (
            .O(N__11693),
            .I(N__11689));
    InMux I__1364 (
            .O(N__11692),
            .I(N__11686));
    Odrv4 I__1363 (
            .O(N__11689),
            .I(\tok.tail_62 ));
    LocalMux I__1362 (
            .O(N__11686),
            .I(\tok.tail_62 ));
    CascadeMux I__1361 (
            .O(N__11681),
            .I(N__11678));
    InMux I__1360 (
            .O(N__11678),
            .I(N__11675));
    LocalMux I__1359 (
            .O(N__11675),
            .I(\tok.C_stk.n5444 ));
    CascadeMux I__1358 (
            .O(N__11672),
            .I(N__11669));
    InMux I__1357 (
            .O(N__11669),
            .I(N__11665));
    InMux I__1356 (
            .O(N__11668),
            .I(N__11662));
    LocalMux I__1355 (
            .O(N__11665),
            .I(\tok.tail_54 ));
    LocalMux I__1354 (
            .O(N__11662),
            .I(\tok.tail_54 ));
    InMux I__1353 (
            .O(N__11657),
            .I(N__11651));
    InMux I__1352 (
            .O(N__11656),
            .I(N__11651));
    LocalMux I__1351 (
            .O(N__11651),
            .I(\tok.C_stk.tail_38 ));
    InMux I__1350 (
            .O(N__11648),
            .I(N__11642));
    InMux I__1349 (
            .O(N__11647),
            .I(N__11642));
    LocalMux I__1348 (
            .O(N__11642),
            .I(\tok.tail_46 ));
    InMux I__1347 (
            .O(N__11639),
            .I(N__11636));
    LocalMux I__1346 (
            .O(N__11636),
            .I(N__11633));
    Span12Mux_s6_v I__1345 (
            .O(N__11633),
            .I(N__11629));
    InMux I__1344 (
            .O(N__11632),
            .I(N__11626));
    Odrv12 I__1343 (
            .O(N__11629),
            .I(sender_1));
    LocalMux I__1342 (
            .O(N__11626),
            .I(sender_1));
    IoInMux I__1341 (
            .O(N__11621),
            .I(N__11618));
    LocalMux I__1340 (
            .O(N__11618),
            .I(N__11615));
    Span4Mux_s1_v I__1339 (
            .O(N__11615),
            .I(N__11612));
    Odrv4 I__1338 (
            .O(N__11612),
            .I(tx_c));
    CascadeMux I__1337 (
            .O(N__11609),
            .I(N__11606));
    InMux I__1336 (
            .O(N__11606),
            .I(N__11600));
    InMux I__1335 (
            .O(N__11605),
            .I(N__11600));
    LocalMux I__1334 (
            .O(N__11600),
            .I(\tok.A_stk.tail_17 ));
    CascadeMux I__1333 (
            .O(N__11597),
            .I(N__11594));
    InMux I__1332 (
            .O(N__11594),
            .I(N__11591));
    LocalMux I__1331 (
            .O(N__11591),
            .I(\tok.tc_7 ));
    CascadeMux I__1330 (
            .O(N__11588),
            .I(\tok.ram.n5600_cascade_ ));
    CascadeMux I__1329 (
            .O(N__11585),
            .I(N__11580));
    InMux I__1328 (
            .O(N__11584),
            .I(N__11576));
    InMux I__1327 (
            .O(N__11583),
            .I(N__11571));
    InMux I__1326 (
            .O(N__11580),
            .I(N__11571));
    InMux I__1325 (
            .O(N__11579),
            .I(N__11568));
    LocalMux I__1324 (
            .O(N__11576),
            .I(\tok.c_stk_r_7 ));
    LocalMux I__1323 (
            .O(N__11571),
            .I(\tok.c_stk_r_7 ));
    LocalMux I__1322 (
            .O(N__11568),
            .I(\tok.c_stk_r_7 ));
    InMux I__1321 (
            .O(N__11561),
            .I(N__11558));
    LocalMux I__1320 (
            .O(N__11558),
            .I(\tok.n5511 ));
    CascadeMux I__1319 (
            .O(N__11555),
            .I(\tok.n3_adj_719_cascade_ ));
    CascadeMux I__1318 (
            .O(N__11552),
            .I(\tok.n5_adj_720_cascade_ ));
    InMux I__1317 (
            .O(N__11549),
            .I(N__11546));
    LocalMux I__1316 (
            .O(N__11546),
            .I(n92_adj_869));
    CascadeMux I__1315 (
            .O(N__11543),
            .I(n92_adj_869_cascade_));
    InMux I__1314 (
            .O(N__11540),
            .I(N__11537));
    LocalMux I__1313 (
            .O(N__11537),
            .I(N__11534));
    Odrv4 I__1312 (
            .O(N__11534),
            .I(\tok.n5507 ));
    InMux I__1311 (
            .O(N__11531),
            .I(N__11527));
    InMux I__1310 (
            .O(N__11530),
            .I(N__11524));
    LocalMux I__1309 (
            .O(N__11527),
            .I(\tok.C_stk.tail_4 ));
    LocalMux I__1308 (
            .O(N__11524),
            .I(\tok.C_stk.tail_4 ));
    InMux I__1307 (
            .O(N__11519),
            .I(N__11516));
    LocalMux I__1306 (
            .O(N__11516),
            .I(n10));
    CascadeMux I__1305 (
            .O(N__11513),
            .I(\tok.n36_cascade_ ));
    CascadeMux I__1304 (
            .O(N__11510),
            .I(\tok.n83_adj_842_cascade_ ));
    CascadeMux I__1303 (
            .O(N__11507),
            .I(\tok.ram.n5597_cascade_ ));
    CascadeMux I__1302 (
            .O(N__11504),
            .I(N__11500));
    InMux I__1301 (
            .O(N__11503),
            .I(N__11492));
    InMux I__1300 (
            .O(N__11500),
            .I(N__11492));
    InMux I__1299 (
            .O(N__11499),
            .I(N__11492));
    LocalMux I__1298 (
            .O(N__11492),
            .I(N__11488));
    InMux I__1297 (
            .O(N__11491),
            .I(N__11485));
    Span4Mux_h I__1296 (
            .O(N__11488),
            .I(N__11482));
    LocalMux I__1295 (
            .O(N__11485),
            .I(\tok.c_stk_r_0 ));
    Odrv4 I__1294 (
            .O(N__11482),
            .I(\tok.c_stk_r_0 ));
    InMux I__1293 (
            .O(N__11477),
            .I(N__11474));
    LocalMux I__1292 (
            .O(N__11474),
            .I(\tok.n5583 ));
    CascadeMux I__1291 (
            .O(N__11471),
            .I(\tok.n3_adj_863_cascade_ ));
    InMux I__1290 (
            .O(N__11468),
            .I(N__11465));
    LocalMux I__1289 (
            .O(N__11465),
            .I(\tok.n5_adj_864 ));
    CascadeMux I__1288 (
            .O(N__11462),
            .I(\tok.n83_adj_714_cascade_ ));
    CascadeMux I__1287 (
            .O(N__11459),
            .I(N__11456));
    InMux I__1286 (
            .O(N__11456),
            .I(N__11452));
    InMux I__1285 (
            .O(N__11455),
            .I(N__11449));
    LocalMux I__1284 (
            .O(N__11452),
            .I(\tok.tail_29 ));
    LocalMux I__1283 (
            .O(N__11449),
            .I(\tok.tail_29 ));
    InMux I__1282 (
            .O(N__11444),
            .I(N__11438));
    InMux I__1281 (
            .O(N__11443),
            .I(N__11438));
    LocalMux I__1280 (
            .O(N__11438),
            .I(\tok.C_stk.tail_37 ));
    CascadeMux I__1279 (
            .O(N__11435),
            .I(N__11432));
    InMux I__1278 (
            .O(N__11432),
            .I(N__11428));
    CascadeMux I__1277 (
            .O(N__11431),
            .I(N__11425));
    LocalMux I__1276 (
            .O(N__11428),
            .I(N__11422));
    InMux I__1275 (
            .O(N__11425),
            .I(N__11419));
    Span4Mux_v I__1274 (
            .O(N__11422),
            .I(N__11416));
    LocalMux I__1273 (
            .O(N__11419),
            .I(N__11413));
    Odrv4 I__1272 (
            .O(N__11416),
            .I(\tok.tail_53 ));
    Odrv4 I__1271 (
            .O(N__11413),
            .I(\tok.tail_53 ));
    CascadeMux I__1270 (
            .O(N__11408),
            .I(N__11404));
    InMux I__1269 (
            .O(N__11407),
            .I(N__11401));
    InMux I__1268 (
            .O(N__11404),
            .I(N__11398));
    LocalMux I__1267 (
            .O(N__11401),
            .I(N__11395));
    LocalMux I__1266 (
            .O(N__11398),
            .I(\tok.tail_45 ));
    Odrv4 I__1265 (
            .O(N__11395),
            .I(\tok.tail_45 ));
    CascadeMux I__1264 (
            .O(N__11390),
            .I(N__11387));
    InMux I__1263 (
            .O(N__11387),
            .I(N__11384));
    LocalMux I__1262 (
            .O(N__11384),
            .I(N__11381));
    Span4Mux_v I__1261 (
            .O(N__11381),
            .I(N__11378));
    Odrv4 I__1260 (
            .O(N__11378),
            .I(\tok.tc_0 ));
    InMux I__1259 (
            .O(N__11375),
            .I(N__11372));
    LocalMux I__1258 (
            .O(N__11372),
            .I(n92));
    CascadeMux I__1257 (
            .O(N__11369),
            .I(n92_cascade_));
    CascadeMux I__1256 (
            .O(N__11366),
            .I(N__11363));
    InMux I__1255 (
            .O(N__11363),
            .I(N__11360));
    LocalMux I__1254 (
            .O(N__11360),
            .I(N__11357));
    Odrv4 I__1253 (
            .O(N__11357),
            .I(\tok.tc_3 ));
    InMux I__1252 (
            .O(N__11354),
            .I(N__11351));
    LocalMux I__1251 (
            .O(N__11351),
            .I(N__11348));
    Odrv4 I__1250 (
            .O(N__11348),
            .I(\tok.n13_adj_646 ));
    CascadeMux I__1249 (
            .O(N__11345),
            .I(n10_cascade_));
    CascadeMux I__1248 (
            .O(N__11342),
            .I(N__11339));
    InMux I__1247 (
            .O(N__11339),
            .I(N__11336));
    LocalMux I__1246 (
            .O(N__11336),
            .I(N__11333));
    Odrv4 I__1245 (
            .O(N__11333),
            .I(\tok.tc_2 ));
    CascadeMux I__1244 (
            .O(N__11330),
            .I(\tok.n31_adj_795_cascade_ ));
    InMux I__1243 (
            .O(N__11327),
            .I(N__11324));
    LocalMux I__1242 (
            .O(N__11324),
            .I(\tok.n5473 ));
    CascadeMux I__1241 (
            .O(N__11321),
            .I(\tok.C_stk.n5441_cascade_ ));
    CascadeMux I__1240 (
            .O(N__11318),
            .I(N__11315));
    InMux I__1239 (
            .O(N__11315),
            .I(N__11309));
    InMux I__1238 (
            .O(N__11314),
            .I(N__11309));
    LocalMux I__1237 (
            .O(N__11309),
            .I(\tok.C_stk.tail_5 ));
    InMux I__1236 (
            .O(N__11306),
            .I(N__11300));
    InMux I__1235 (
            .O(N__11305),
            .I(N__11300));
    LocalMux I__1234 (
            .O(N__11300),
            .I(\tok.tail_13 ));
    CascadeMux I__1233 (
            .O(N__11297),
            .I(N__11293));
    InMux I__1232 (
            .O(N__11296),
            .I(N__11290));
    InMux I__1231 (
            .O(N__11293),
            .I(N__11287));
    LocalMux I__1230 (
            .O(N__11290),
            .I(\tok.C_stk.tail_21 ));
    LocalMux I__1229 (
            .O(N__11287),
            .I(\tok.C_stk.tail_21 ));
    CascadeMux I__1228 (
            .O(N__11282),
            .I(\tok.uart.n2_cascade_ ));
    SRMux I__1227 (
            .O(N__11279),
            .I(N__11276));
    LocalMux I__1226 (
            .O(N__11276),
            .I(N__11273));
    Span4Mux_s2_h I__1225 (
            .O(N__11273),
            .I(N__11270));
    Odrv4 I__1224 (
            .O(N__11270),
            .I(\tok.uart.rxclkcounter_6__N_477 ));
    InMux I__1223 (
            .O(N__11267),
            .I(N__11257));
    InMux I__1222 (
            .O(N__11266),
            .I(N__11257));
    InMux I__1221 (
            .O(N__11265),
            .I(N__11257));
    InMux I__1220 (
            .O(N__11264),
            .I(N__11254));
    LocalMux I__1219 (
            .O(N__11257),
            .I(N__11251));
    LocalMux I__1218 (
            .O(N__11254),
            .I(\tok.uart.bytephase_2 ));
    Odrv4 I__1217 (
            .O(N__11251),
            .I(\tok.uart.bytephase_2 ));
    CascadeMux I__1216 (
            .O(N__11246),
            .I(\tok.uart.n13_cascade_ ));
    InMux I__1215 (
            .O(N__11243),
            .I(N__11233));
    InMux I__1214 (
            .O(N__11242),
            .I(N__11233));
    InMux I__1213 (
            .O(N__11241),
            .I(N__11233));
    InMux I__1212 (
            .O(N__11240),
            .I(N__11230));
    LocalMux I__1211 (
            .O(N__11233),
            .I(N__11227));
    LocalMux I__1210 (
            .O(N__11230),
            .I(\tok.uart.bytephase_4 ));
    Odrv4 I__1209 (
            .O(N__11227),
            .I(\tok.uart.bytephase_4 ));
    SRMux I__1208 (
            .O(N__11222),
            .I(N__11219));
    LocalMux I__1207 (
            .O(N__11219),
            .I(N__11215));
    InMux I__1206 (
            .O(N__11218),
            .I(N__11212));
    Span4Mux_s1_v I__1205 (
            .O(N__11215),
            .I(N__11207));
    LocalMux I__1204 (
            .O(N__11212),
            .I(N__11207));
    Odrv4 I__1203 (
            .O(N__11207),
            .I(bytephase_5__N_510));
    CascadeMux I__1202 (
            .O(N__11204),
            .I(N__11198));
    InMux I__1201 (
            .O(N__11203),
            .I(N__11195));
    InMux I__1200 (
            .O(N__11202),
            .I(N__11188));
    InMux I__1199 (
            .O(N__11201),
            .I(N__11188));
    InMux I__1198 (
            .O(N__11198),
            .I(N__11188));
    LocalMux I__1197 (
            .O(N__11195),
            .I(N__11182));
    LocalMux I__1196 (
            .O(N__11188),
            .I(N__11182));
    InMux I__1195 (
            .O(N__11187),
            .I(N__11179));
    Span4Mux_v I__1194 (
            .O(N__11182),
            .I(N__11176));
    LocalMux I__1193 (
            .O(N__11179),
            .I(\tok.uart.bytephase_0 ));
    Odrv4 I__1192 (
            .O(N__11176),
            .I(\tok.uart.bytephase_0 ));
    InMux I__1191 (
            .O(N__11171),
            .I(N__11165));
    InMux I__1190 (
            .O(N__11170),
            .I(N__11165));
    LocalMux I__1189 (
            .O(N__11165),
            .I(N__11162));
    Odrv4 I__1188 (
            .O(N__11162),
            .I(n813));
    InMux I__1187 (
            .O(N__11159),
            .I(N__11146));
    InMux I__1186 (
            .O(N__11158),
            .I(N__11146));
    InMux I__1185 (
            .O(N__11157),
            .I(N__11146));
    InMux I__1184 (
            .O(N__11156),
            .I(N__11146));
    InMux I__1183 (
            .O(N__11155),
            .I(N__11143));
    LocalMux I__1182 (
            .O(N__11146),
            .I(N__11140));
    LocalMux I__1181 (
            .O(N__11143),
            .I(\tok.uart.bytephase_1 ));
    Odrv12 I__1180 (
            .O(N__11140),
            .I(\tok.uart.bytephase_1 ));
    CascadeMux I__1179 (
            .O(N__11135),
            .I(N__11132));
    InMux I__1178 (
            .O(N__11132),
            .I(N__11127));
    InMux I__1177 (
            .O(N__11131),
            .I(N__11123));
    InMux I__1176 (
            .O(N__11130),
            .I(N__11120));
    LocalMux I__1175 (
            .O(N__11127),
            .I(N__11117));
    InMux I__1174 (
            .O(N__11126),
            .I(N__11114));
    LocalMux I__1173 (
            .O(N__11123),
            .I(\tok.c_stk_r_2 ));
    LocalMux I__1172 (
            .O(N__11120),
            .I(\tok.c_stk_r_2 ));
    Odrv4 I__1171 (
            .O(N__11117),
            .I(\tok.c_stk_r_2 ));
    LocalMux I__1170 (
            .O(N__11114),
            .I(\tok.c_stk_r_2 ));
    InMux I__1169 (
            .O(N__11105),
            .I(N__11102));
    LocalMux I__1168 (
            .O(N__11102),
            .I(\tok.ram.n5585 ));
    CascadeMux I__1167 (
            .O(N__11099),
            .I(\tok.n3_adj_645_cascade_ ));
    InMux I__1166 (
            .O(N__11096),
            .I(N__11093));
    LocalMux I__1165 (
            .O(N__11093),
            .I(\tok.n83 ));
    InMux I__1164 (
            .O(N__11090),
            .I(N__11087));
    LocalMux I__1163 (
            .O(N__11087),
            .I(\tok.n5603 ));
    InMux I__1162 (
            .O(N__11084),
            .I(N__11080));
    InMux I__1161 (
            .O(N__11083),
            .I(N__11077));
    LocalMux I__1160 (
            .O(N__11080),
            .I(N__11074));
    LocalMux I__1159 (
            .O(N__11077),
            .I(\tok.uart.txclkcounter_5 ));
    Odrv4 I__1158 (
            .O(N__11074),
            .I(\tok.uart.txclkcounter_5 ));
    InMux I__1157 (
            .O(N__11069),
            .I(N__11065));
    InMux I__1156 (
            .O(N__11068),
            .I(N__11062));
    LocalMux I__1155 (
            .O(N__11065),
            .I(\tok.uart.txclkcounter_2 ));
    LocalMux I__1154 (
            .O(N__11062),
            .I(\tok.uart.txclkcounter_2 ));
    CascadeMux I__1153 (
            .O(N__11057),
            .I(N__11053));
    InMux I__1152 (
            .O(N__11056),
            .I(N__11050));
    InMux I__1151 (
            .O(N__11053),
            .I(N__11047));
    LocalMux I__1150 (
            .O(N__11050),
            .I(\tok.uart.txclkcounter_8 ));
    LocalMux I__1149 (
            .O(N__11047),
            .I(\tok.uart.txclkcounter_8 ));
    InMux I__1148 (
            .O(N__11042),
            .I(N__11038));
    InMux I__1147 (
            .O(N__11041),
            .I(N__11035));
    LocalMux I__1146 (
            .O(N__11038),
            .I(\tok.uart.txclkcounter_3 ));
    LocalMux I__1145 (
            .O(N__11035),
            .I(\tok.uart.txclkcounter_3 ));
    CascadeMux I__1144 (
            .O(N__11030),
            .I(N__11025));
    InMux I__1143 (
            .O(N__11029),
            .I(N__11018));
    InMux I__1142 (
            .O(N__11028),
            .I(N__11018));
    InMux I__1141 (
            .O(N__11025),
            .I(N__11018));
    LocalMux I__1140 (
            .O(N__11018),
            .I(\tok.uart.sentbits_2 ));
    InMux I__1139 (
            .O(N__11015),
            .I(N__11011));
    InMux I__1138 (
            .O(N__11014),
            .I(N__11008));
    LocalMux I__1137 (
            .O(N__11011),
            .I(\tok.uart.txclkcounter_4 ));
    LocalMux I__1136 (
            .O(N__11008),
            .I(\tok.uart.txclkcounter_4 ));
    InMux I__1135 (
            .O(N__11003),
            .I(N__10999));
    InMux I__1134 (
            .O(N__11002),
            .I(N__10996));
    LocalMux I__1133 (
            .O(N__10999),
            .I(\tok.uart.txclkcounter_7 ));
    LocalMux I__1132 (
            .O(N__10996),
            .I(\tok.uart.txclkcounter_7 ));
    InMux I__1131 (
            .O(N__10991),
            .I(N__10987));
    InMux I__1130 (
            .O(N__10990),
            .I(N__10984));
    LocalMux I__1129 (
            .O(N__10987),
            .I(\tok.uart.txclkcounter_6 ));
    LocalMux I__1128 (
            .O(N__10984),
            .I(\tok.uart.txclkcounter_6 ));
    InMux I__1127 (
            .O(N__10979),
            .I(N__10975));
    InMux I__1126 (
            .O(N__10978),
            .I(N__10972));
    LocalMux I__1125 (
            .O(N__10975),
            .I(\tok.uart.txclkcounter_0 ));
    LocalMux I__1124 (
            .O(N__10972),
            .I(\tok.uart.txclkcounter_0 ));
    InMux I__1123 (
            .O(N__10967),
            .I(N__10963));
    InMux I__1122 (
            .O(N__10966),
            .I(N__10960));
    LocalMux I__1121 (
            .O(N__10963),
            .I(\tok.uart.txclkcounter_1 ));
    LocalMux I__1120 (
            .O(N__10960),
            .I(\tok.uart.txclkcounter_1 ));
    CascadeMux I__1119 (
            .O(N__10955),
            .I(\tok.uart.n5418_cascade_ ));
    InMux I__1118 (
            .O(N__10952),
            .I(N__10949));
    LocalMux I__1117 (
            .O(N__10949),
            .I(\tok.uart.n12 ));
    CascadeMux I__1116 (
            .O(N__10946),
            .I(txtick_cascade_));
    CascadeMux I__1115 (
            .O(N__10943),
            .I(N__10940));
    InMux I__1114 (
            .O(N__10940),
            .I(N__10937));
    LocalMux I__1113 (
            .O(N__10937),
            .I(N__10934));
    Span4Mux_v I__1112 (
            .O(N__10934),
            .I(N__10930));
    InMux I__1111 (
            .O(N__10933),
            .I(N__10927));
    Odrv4 I__1110 (
            .O(N__10930),
            .I(\tok.tail_61 ));
    LocalMux I__1109 (
            .O(N__10927),
            .I(\tok.tail_61 ));
    InMux I__1108 (
            .O(N__10922),
            .I(\tok.uart.n4826 ));
    InMux I__1107 (
            .O(N__10919),
            .I(N__10915));
    InMux I__1106 (
            .O(N__10918),
            .I(N__10912));
    LocalMux I__1105 (
            .O(N__10915),
            .I(\tok.uart.rxclkcounter_5 ));
    LocalMux I__1104 (
            .O(N__10912),
            .I(\tok.uart.rxclkcounter_5 ));
    InMux I__1103 (
            .O(N__10907),
            .I(N__10903));
    InMux I__1102 (
            .O(N__10906),
            .I(N__10900));
    LocalMux I__1101 (
            .O(N__10903),
            .I(\tok.uart.rxclkcounter_3 ));
    LocalMux I__1100 (
            .O(N__10900),
            .I(\tok.uart.rxclkcounter_3 ));
    CascadeMux I__1099 (
            .O(N__10895),
            .I(N__10891));
    InMux I__1098 (
            .O(N__10894),
            .I(N__10888));
    InMux I__1097 (
            .O(N__10891),
            .I(N__10885));
    LocalMux I__1096 (
            .O(N__10888),
            .I(N__10880));
    LocalMux I__1095 (
            .O(N__10885),
            .I(N__10880));
    Odrv4 I__1094 (
            .O(N__10880),
            .I(\tok.uart.rxclkcounter_2 ));
    CascadeMux I__1093 (
            .O(N__10877),
            .I(n813_cascade_));
    CEMux I__1092 (
            .O(N__10874),
            .I(N__10871));
    LocalMux I__1091 (
            .O(N__10871),
            .I(N__10868));
    Span4Mux_s2_v I__1090 (
            .O(N__10868),
            .I(N__10865));
    Odrv4 I__1089 (
            .O(N__10865),
            .I(n971));
    InMux I__1088 (
            .O(N__10862),
            .I(N__10858));
    InMux I__1087 (
            .O(N__10861),
            .I(N__10855));
    LocalMux I__1086 (
            .O(N__10858),
            .I(\tok.uart.rxclkcounter_6 ));
    LocalMux I__1085 (
            .O(N__10855),
            .I(\tok.uart.rxclkcounter_6 ));
    InMux I__1084 (
            .O(N__10850),
            .I(N__10846));
    InMux I__1083 (
            .O(N__10849),
            .I(N__10843));
    LocalMux I__1082 (
            .O(N__10846),
            .I(\tok.uart.rxclkcounter_0 ));
    LocalMux I__1081 (
            .O(N__10843),
            .I(\tok.uart.rxclkcounter_0 ));
    CascadeMux I__1080 (
            .O(N__10838),
            .I(N__10834));
    InMux I__1079 (
            .O(N__10837),
            .I(N__10831));
    InMux I__1078 (
            .O(N__10834),
            .I(N__10828));
    LocalMux I__1077 (
            .O(N__10831),
            .I(\tok.uart.rxclkcounter_4 ));
    LocalMux I__1076 (
            .O(N__10828),
            .I(\tok.uart.rxclkcounter_4 ));
    InMux I__1075 (
            .O(N__10823),
            .I(N__10819));
    InMux I__1074 (
            .O(N__10822),
            .I(N__10816));
    LocalMux I__1073 (
            .O(N__10819),
            .I(\tok.uart.rxclkcounter_1 ));
    LocalMux I__1072 (
            .O(N__10816),
            .I(\tok.uart.rxclkcounter_1 ));
    InMux I__1071 (
            .O(N__10811),
            .I(N__10808));
    LocalMux I__1070 (
            .O(N__10808),
            .I(\tok.uart.n12_adj_640 ));
    InMux I__1069 (
            .O(N__10805),
            .I(N__10799));
    InMux I__1068 (
            .O(N__10804),
            .I(N__10799));
    LocalMux I__1067 (
            .O(N__10799),
            .I(\tok.uart.sentbits_3 ));
    CascadeMux I__1066 (
            .O(N__10796),
            .I(N__10793));
    InMux I__1065 (
            .O(N__10793),
            .I(N__10789));
    InMux I__1064 (
            .O(N__10792),
            .I(N__10786));
    LocalMux I__1063 (
            .O(N__10789),
            .I(N__10783));
    LocalMux I__1062 (
            .O(N__10786),
            .I(\tok.tail_12 ));
    Odrv4 I__1061 (
            .O(N__10783),
            .I(\tok.tail_12 ));
    CascadeMux I__1060 (
            .O(N__10778),
            .I(N__10774));
    CascadeMux I__1059 (
            .O(N__10777),
            .I(N__10771));
    InMux I__1058 (
            .O(N__10774),
            .I(N__10766));
    InMux I__1057 (
            .O(N__10771),
            .I(N__10766));
    LocalMux I__1056 (
            .O(N__10766),
            .I(\tok.C_stk.tail_20 ));
    InMux I__1055 (
            .O(N__10763),
            .I(N__10757));
    InMux I__1054 (
            .O(N__10762),
            .I(N__10757));
    LocalMux I__1053 (
            .O(N__10757),
            .I(\tok.tail_28 ));
    InMux I__1052 (
            .O(N__10754),
            .I(N__10748));
    InMux I__1051 (
            .O(N__10753),
            .I(N__10748));
    LocalMux I__1050 (
            .O(N__10748),
            .I(\tok.C_stk.tail_36 ));
    CascadeMux I__1049 (
            .O(N__10745),
            .I(N__10741));
    CascadeMux I__1048 (
            .O(N__10744),
            .I(N__10738));
    InMux I__1047 (
            .O(N__10741),
            .I(N__10735));
    InMux I__1046 (
            .O(N__10738),
            .I(N__10732));
    LocalMux I__1045 (
            .O(N__10735),
            .I(N__10727));
    LocalMux I__1044 (
            .O(N__10732),
            .I(N__10727));
    Odrv4 I__1043 (
            .O(N__10727),
            .I(\tok.tail_52 ));
    CascadeMux I__1042 (
            .O(N__10724),
            .I(N__10720));
    InMux I__1041 (
            .O(N__10723),
            .I(N__10717));
    InMux I__1040 (
            .O(N__10720),
            .I(N__10714));
    LocalMux I__1039 (
            .O(N__10717),
            .I(N__10711));
    LocalMux I__1038 (
            .O(N__10714),
            .I(\tok.tail_44 ));
    Odrv4 I__1037 (
            .O(N__10711),
            .I(\tok.tail_44 ));
    InMux I__1036 (
            .O(N__10706),
            .I(bfn_2_2_0_));
    InMux I__1035 (
            .O(N__10703),
            .I(\tok.uart.n4822 ));
    InMux I__1034 (
            .O(N__10700),
            .I(\tok.uart.n4823 ));
    InMux I__1033 (
            .O(N__10697),
            .I(\tok.uart.n4824 ));
    InMux I__1032 (
            .O(N__10694),
            .I(\tok.uart.n4825 ));
    CascadeMux I__1031 (
            .O(N__10691),
            .I(\tok.C_stk.n5435_cascade_ ));
    InMux I__1030 (
            .O(N__10688),
            .I(N__10684));
    InMux I__1029 (
            .O(N__10687),
            .I(N__10681));
    LocalMux I__1028 (
            .O(N__10684),
            .I(\tok.C_stk.tail_7 ));
    LocalMux I__1027 (
            .O(N__10681),
            .I(\tok.C_stk.tail_7 ));
    InMux I__1026 (
            .O(N__10676),
            .I(N__10670));
    InMux I__1025 (
            .O(N__10675),
            .I(N__10670));
    LocalMux I__1024 (
            .O(N__10670),
            .I(\tok.tail_15 ));
    CascadeMux I__1023 (
            .O(N__10667),
            .I(N__10663));
    CascadeMux I__1022 (
            .O(N__10666),
            .I(N__10660));
    InMux I__1021 (
            .O(N__10663),
            .I(N__10655));
    InMux I__1020 (
            .O(N__10660),
            .I(N__10655));
    LocalMux I__1019 (
            .O(N__10655),
            .I(\tok.C_stk.tail_23 ));
    InMux I__1018 (
            .O(N__10652),
            .I(N__10646));
    InMux I__1017 (
            .O(N__10651),
            .I(N__10646));
    LocalMux I__1016 (
            .O(N__10646),
            .I(\tok.tail_31 ));
    InMux I__1015 (
            .O(N__10643),
            .I(N__10637));
    InMux I__1014 (
            .O(N__10642),
            .I(N__10637));
    LocalMux I__1013 (
            .O(N__10637),
            .I(\tok.C_stk.tail_39 ));
    CascadeMux I__1012 (
            .O(N__10634),
            .I(N__10630));
    CascadeMux I__1011 (
            .O(N__10633),
            .I(N__10627));
    InMux I__1010 (
            .O(N__10630),
            .I(N__10624));
    InMux I__1009 (
            .O(N__10627),
            .I(N__10621));
    LocalMux I__1008 (
            .O(N__10624),
            .I(N__10618));
    LocalMux I__1007 (
            .O(N__10621),
            .I(\tok.tail_55 ));
    Odrv4 I__1006 (
            .O(N__10618),
            .I(\tok.tail_55 ));
    CascadeMux I__1005 (
            .O(N__10613),
            .I(N__10610));
    InMux I__1004 (
            .O(N__10610),
            .I(N__10606));
    InMux I__1003 (
            .O(N__10609),
            .I(N__10603));
    LocalMux I__1002 (
            .O(N__10606),
            .I(N__10600));
    LocalMux I__1001 (
            .O(N__10603),
            .I(\tok.tail_47 ));
    Odrv4 I__1000 (
            .O(N__10600),
            .I(\tok.tail_47 ));
    CascadeMux I__999 (
            .O(N__10595),
            .I(N__10592));
    InMux I__998 (
            .O(N__10592),
            .I(N__10588));
    InMux I__997 (
            .O(N__10591),
            .I(N__10585));
    LocalMux I__996 (
            .O(N__10588),
            .I(\tok.tail_60 ));
    LocalMux I__995 (
            .O(N__10585),
            .I(\tok.tail_60 ));
    CascadeMux I__994 (
            .O(N__10580),
            .I(N__10576));
    CascadeMux I__993 (
            .O(N__10579),
            .I(N__10573));
    InMux I__992 (
            .O(N__10576),
            .I(N__10570));
    InMux I__991 (
            .O(N__10573),
            .I(N__10567));
    LocalMux I__990 (
            .O(N__10570),
            .I(N__10564));
    LocalMux I__989 (
            .O(N__10567),
            .I(\tok.tail_51 ));
    Odrv4 I__988 (
            .O(N__10564),
            .I(\tok.tail_51 ));
    CascadeMux I__987 (
            .O(N__10559),
            .I(N__10556));
    InMux I__986 (
            .O(N__10556),
            .I(N__10552));
    InMux I__985 (
            .O(N__10555),
            .I(N__10549));
    LocalMux I__984 (
            .O(N__10552),
            .I(\tok.tail_59 ));
    LocalMux I__983 (
            .O(N__10549),
            .I(\tok.tail_59 ));
    CascadeMux I__982 (
            .O(N__10544),
            .I(N__10541));
    InMux I__981 (
            .O(N__10541),
            .I(N__10537));
    InMux I__980 (
            .O(N__10540),
            .I(N__10534));
    LocalMux I__979 (
            .O(N__10537),
            .I(N__10531));
    LocalMux I__978 (
            .O(N__10534),
            .I(\tok.tail_50 ));
    Odrv4 I__977 (
            .O(N__10531),
            .I(\tok.tail_50 ));
    CascadeMux I__976 (
            .O(N__10526),
            .I(N__10523));
    InMux I__975 (
            .O(N__10523),
            .I(N__10519));
    InMux I__974 (
            .O(N__10522),
            .I(N__10516));
    LocalMux I__973 (
            .O(N__10519),
            .I(\tok.tail_58 ));
    LocalMux I__972 (
            .O(N__10516),
            .I(\tok.tail_58 ));
    InMux I__971 (
            .O(N__10511),
            .I(N__10507));
    CascadeMux I__970 (
            .O(N__10510),
            .I(N__10504));
    LocalMux I__969 (
            .O(N__10507),
            .I(N__10501));
    InMux I__968 (
            .O(N__10504),
            .I(N__10498));
    Odrv4 I__967 (
            .O(N__10501),
            .I(\tok.tail_49 ));
    LocalMux I__966 (
            .O(N__10498),
            .I(\tok.tail_49 ));
    CascadeMux I__965 (
            .O(N__10493),
            .I(N__10490));
    InMux I__964 (
            .O(N__10490),
            .I(N__10487));
    LocalMux I__963 (
            .O(N__10487),
            .I(N__10483));
    InMux I__962 (
            .O(N__10486),
            .I(N__10480));
    Odrv4 I__961 (
            .O(N__10483),
            .I(\tok.tail_57 ));
    LocalMux I__960 (
            .O(N__10480),
            .I(\tok.tail_57 ));
    CascadeMux I__959 (
            .O(N__10475),
            .I(N__10471));
    CascadeMux I__958 (
            .O(N__10474),
            .I(N__10468));
    InMux I__957 (
            .O(N__10471),
            .I(N__10465));
    InMux I__956 (
            .O(N__10468),
            .I(N__10462));
    LocalMux I__955 (
            .O(N__10465),
            .I(N__10459));
    LocalMux I__954 (
            .O(N__10462),
            .I(\tok.tail_48 ));
    Odrv4 I__953 (
            .O(N__10459),
            .I(\tok.tail_48 ));
    CascadeMux I__952 (
            .O(N__10454),
            .I(N__10451));
    InMux I__951 (
            .O(N__10451),
            .I(N__10447));
    InMux I__950 (
            .O(N__10450),
            .I(N__10444));
    LocalMux I__949 (
            .O(N__10447),
            .I(\tok.tail_56 ));
    LocalMux I__948 (
            .O(N__10444),
            .I(\tok.tail_56 ));
    InMux I__947 (
            .O(N__10439),
            .I(N__10435));
    InMux I__946 (
            .O(N__10438),
            .I(N__10432));
    LocalMux I__945 (
            .O(N__10435),
            .I(\tok.tail_63 ));
    LocalMux I__944 (
            .O(N__10432),
            .I(\tok.tail_63 ));
    CascadeMux I__943 (
            .O(N__10427),
            .I(N__10423));
    CascadeMux I__942 (
            .O(N__10426),
            .I(N__10420));
    InMux I__941 (
            .O(N__10423),
            .I(N__10415));
    InMux I__940 (
            .O(N__10420),
            .I(N__10415));
    LocalMux I__939 (
            .O(N__10415),
            .I(\tok.C_stk.tail_18 ));
    CascadeMux I__938 (
            .O(N__10412),
            .I(N__10408));
    CascadeMux I__937 (
            .O(N__10411),
            .I(N__10405));
    InMux I__936 (
            .O(N__10408),
            .I(N__10400));
    InMux I__935 (
            .O(N__10405),
            .I(N__10400));
    LocalMux I__934 (
            .O(N__10400),
            .I(\tok.tail_26 ));
    InMux I__933 (
            .O(N__10397),
            .I(N__10391));
    InMux I__932 (
            .O(N__10396),
            .I(N__10391));
    LocalMux I__931 (
            .O(N__10391),
            .I(\tok.C_stk.tail_34 ));
    CascadeMux I__930 (
            .O(N__10388),
            .I(N__10385));
    InMux I__929 (
            .O(N__10385),
            .I(N__10381));
    InMux I__928 (
            .O(N__10384),
            .I(N__10378));
    LocalMux I__927 (
            .O(N__10381),
            .I(\tok.tail_43 ));
    LocalMux I__926 (
            .O(N__10378),
            .I(\tok.tail_43 ));
    InMux I__925 (
            .O(N__10373),
            .I(N__10369));
    InMux I__924 (
            .O(N__10372),
            .I(N__10366));
    LocalMux I__923 (
            .O(N__10369),
            .I(\tok.tail_42 ));
    LocalMux I__922 (
            .O(N__10366),
            .I(\tok.tail_42 ));
    CascadeMux I__921 (
            .O(N__10361),
            .I(N__10357));
    InMux I__920 (
            .O(N__10360),
            .I(N__10354));
    InMux I__919 (
            .O(N__10357),
            .I(N__10351));
    LocalMux I__918 (
            .O(N__10354),
            .I(N__10348));
    LocalMux I__917 (
            .O(N__10351),
            .I(\tok.tail_41 ));
    Odrv4 I__916 (
            .O(N__10348),
            .I(\tok.tail_41 ));
    CascadeMux I__915 (
            .O(N__10343),
            .I(N__10339));
    InMux I__914 (
            .O(N__10342),
            .I(N__10336));
    InMux I__913 (
            .O(N__10339),
            .I(N__10333));
    LocalMux I__912 (
            .O(N__10336),
            .I(N__10330));
    LocalMux I__911 (
            .O(N__10333),
            .I(\tok.tail_40 ));
    Odrv4 I__910 (
            .O(N__10330),
            .I(\tok.tail_40 ));
    InMux I__909 (
            .O(N__10325),
            .I(N__10321));
    InMux I__908 (
            .O(N__10324),
            .I(N__10318));
    LocalMux I__907 (
            .O(N__10321),
            .I(\tok.C_stk.tail_1 ));
    LocalMux I__906 (
            .O(N__10318),
            .I(\tok.C_stk.tail_1 ));
    CascadeMux I__905 (
            .O(N__10313),
            .I(N__10309));
    InMux I__904 (
            .O(N__10312),
            .I(N__10304));
    InMux I__903 (
            .O(N__10309),
            .I(N__10304));
    LocalMux I__902 (
            .O(N__10304),
            .I(\tok.tail_9 ));
    InMux I__901 (
            .O(N__10301),
            .I(N__10295));
    InMux I__900 (
            .O(N__10300),
            .I(N__10295));
    LocalMux I__899 (
            .O(N__10295),
            .I(\tok.C_stk.tail_17 ));
    InMux I__898 (
            .O(N__10292),
            .I(N__10286));
    InMux I__897 (
            .O(N__10291),
            .I(N__10286));
    LocalMux I__896 (
            .O(N__10286),
            .I(\tok.tail_25 ));
    InMux I__895 (
            .O(N__10283),
            .I(N__10277));
    InMux I__894 (
            .O(N__10282),
            .I(N__10277));
    LocalMux I__893 (
            .O(N__10277),
            .I(\tok.C_stk.tail_33 ));
    CascadeMux I__892 (
            .O(N__10274),
            .I(\tok.C_stk.n5450_cascade_ ));
    InMux I__891 (
            .O(N__10271),
            .I(N__10267));
    InMux I__890 (
            .O(N__10270),
            .I(N__10264));
    LocalMux I__889 (
            .O(N__10267),
            .I(\tok.C_stk.tail_2 ));
    LocalMux I__888 (
            .O(N__10264),
            .I(\tok.C_stk.tail_2 ));
    InMux I__887 (
            .O(N__10259),
            .I(N__10253));
    InMux I__886 (
            .O(N__10258),
            .I(N__10253));
    LocalMux I__885 (
            .O(N__10253),
            .I(\tok.tail_10 ));
    InMux I__884 (
            .O(N__10250),
            .I(\tok.uart.n4816 ));
    InMux I__883 (
            .O(N__10247),
            .I(\tok.uart.n4817 ));
    InMux I__882 (
            .O(N__10244),
            .I(\tok.uart.n4818 ));
    InMux I__881 (
            .O(N__10241),
            .I(\tok.uart.n4819 ));
    InMux I__880 (
            .O(N__10238),
            .I(\tok.uart.n4820 ));
    InMux I__879 (
            .O(N__10235),
            .I(bfn_1_5_0_));
    CascadeMux I__878 (
            .O(N__10232),
            .I(\tok.C_stk.n5453_cascade_ ));
    InMux I__877 (
            .O(N__10229),
            .I(\tok.uart.n4827 ));
    InMux I__876 (
            .O(N__10226),
            .I(\tok.uart.n4828 ));
    InMux I__875 (
            .O(N__10223),
            .I(\tok.uart.n4829 ));
    InMux I__874 (
            .O(N__10220),
            .I(\tok.uart.n4830 ));
    InMux I__873 (
            .O(N__10217),
            .I(\tok.uart.n4831 ));
    InMux I__872 (
            .O(N__10214),
            .I(\tok.uart.n4832 ));
    InMux I__871 (
            .O(N__10211),
            .I(bfn_1_4_0_));
    InMux I__870 (
            .O(N__10208),
            .I(\tok.uart.n4814 ));
    InMux I__869 (
            .O(N__10205),
            .I(\tok.uart.n4815 ));
    CascadeMux I__868 (
            .O(N__10202),
            .I(\tok.C_stk.n5456_cascade_ ));
    CascadeMux I__867 (
            .O(N__10199),
            .I(N__10196));
    InMux I__866 (
            .O(N__10196),
            .I(N__10190));
    InMux I__865 (
            .O(N__10195),
            .I(N__10190));
    LocalMux I__864 (
            .O(N__10190),
            .I(\tok.C_stk.tail_0 ));
    CascadeMux I__863 (
            .O(N__10187),
            .I(N__10183));
    CascadeMux I__862 (
            .O(N__10186),
            .I(N__10180));
    InMux I__861 (
            .O(N__10183),
            .I(N__10175));
    InMux I__860 (
            .O(N__10180),
            .I(N__10175));
    LocalMux I__859 (
            .O(N__10175),
            .I(\tok.tail_8 ));
    CascadeMux I__858 (
            .O(N__10172),
            .I(N__10168));
    InMux I__857 (
            .O(N__10171),
            .I(N__10165));
    InMux I__856 (
            .O(N__10168),
            .I(N__10162));
    LocalMux I__855 (
            .O(N__10165),
            .I(N__10157));
    LocalMux I__854 (
            .O(N__10162),
            .I(N__10157));
    Odrv4 I__853 (
            .O(N__10157),
            .I(\tok.C_stk.tail_16 ));
    InMux I__852 (
            .O(N__10154),
            .I(N__10148));
    InMux I__851 (
            .O(N__10153),
            .I(N__10148));
    LocalMux I__850 (
            .O(N__10148),
            .I(\tok.tail_24 ));
    InMux I__849 (
            .O(N__10145),
            .I(N__10139));
    InMux I__848 (
            .O(N__10144),
            .I(N__10139));
    LocalMux I__847 (
            .O(N__10139),
            .I(\tok.C_stk.tail_32 ));
    InMux I__846 (
            .O(N__10136),
            .I(bfn_1_3_0_));
    CascadeMux I__845 (
            .O(N__10133),
            .I(\tok.C_stk.n5447_cascade_ ));
    CascadeMux I__844 (
            .O(N__10130),
            .I(N__10127));
    InMux I__843 (
            .O(N__10127),
            .I(N__10121));
    InMux I__842 (
            .O(N__10126),
            .I(N__10121));
    LocalMux I__841 (
            .O(N__10121),
            .I(\tok.C_stk.tail_3 ));
    CascadeMux I__840 (
            .O(N__10118),
            .I(N__10114));
    InMux I__839 (
            .O(N__10117),
            .I(N__10111));
    InMux I__838 (
            .O(N__10114),
            .I(N__10108));
    LocalMux I__837 (
            .O(N__10111),
            .I(\tok.tail_11 ));
    LocalMux I__836 (
            .O(N__10108),
            .I(\tok.tail_11 ));
    InMux I__835 (
            .O(N__10103),
            .I(N__10097));
    InMux I__834 (
            .O(N__10102),
            .I(N__10097));
    LocalMux I__833 (
            .O(N__10097),
            .I(\tok.C_stk.tail_19 ));
    InMux I__832 (
            .O(N__10094),
            .I(N__10088));
    InMux I__831 (
            .O(N__10093),
            .I(N__10088));
    LocalMux I__830 (
            .O(N__10088),
            .I(\tok.tail_27 ));
    CascadeMux I__829 (
            .O(N__10085),
            .I(N__10082));
    InMux I__828 (
            .O(N__10082),
            .I(N__10078));
    InMux I__827 (
            .O(N__10081),
            .I(N__10075));
    LocalMux I__826 (
            .O(N__10078),
            .I(\tok.C_stk.tail_35 ));
    LocalMux I__825 (
            .O(N__10075),
            .I(\tok.C_stk.tail_35 ));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(\tok.uart.n4821 ),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_2_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_2_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\tok.n4776 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\tok.n4783_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\tok.n4768 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\tok.n4806 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\tok.n4791 ),
            .carryinitout(bfn_8_8_0_));
    GND GND (
            .Y(GNDG0));
    defparam OSCInst0.CLKHF_DIV="0b01";
    SB_HFOSC OSCInst0 (
            .CLKHFPU(N__24259),
            .CLKHFEN(N__24258),
            .CLKHF(clk));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i3_LC_0_7_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i3_LC_0_7_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i3_LC_0_7_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.tail_i0_i3_LC_0_7_0  (
            .in0(N__13601),
            .in1(N__14010),
            .in2(N__15017),
            .in3(N__10117),
            .lcout(\tok.C_stk.tail_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28473),
            .ce(N__13370),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i5274_3_lut_LC_0_7_1 .C_ON=1'b0;
    defparam \tok.C_stk.i5274_3_lut_LC_0_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i5274_3_lut_LC_0_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i5274_3_lut_LC_0_7_1  (
            .in0(N__10126),
            .in1(N__14264),
            .in2(_gnd_net_),
            .in3(N__14981),
            .lcout(),
            .ltout(\tok.C_stk.n5447_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i3_LC_0_7_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i3_LC_0_7_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i3_LC_0_7_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i3_LC_0_7_2  (
            .in0(N__14188),
            .in1(N__15543),
            .in2(N__10133),
            .in3(N__13091),
            .lcout(\tok.c_stk_r_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28473),
            .ce(N__13370),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i11_LC_0_7_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i11_LC_0_7_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i11_LC_0_7_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i11_LC_0_7_3  (
            .in0(N__14007),
            .in1(N__10103),
            .in2(N__10130),
            .in3(N__13602),
            .lcout(\tok.tail_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28473),
            .ce(N__13370),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i19_LC_0_7_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i19_LC_0_7_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i19_LC_0_7_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i19_LC_0_7_4  (
            .in0(N__13599),
            .in1(N__10094),
            .in2(N__10118),
            .in3(N__14011),
            .lcout(\tok.C_stk.tail_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28473),
            .ce(N__13370),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i27_LC_0_7_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i27_LC_0_7_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i27_LC_0_7_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i27_LC_0_7_5  (
            .in0(N__14008),
            .in1(N__10102),
            .in2(N__10085),
            .in3(N__13603),
            .lcout(\tok.tail_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28473),
            .ce(N__13370),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i35_LC_0_7_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i35_LC_0_7_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i35_LC_0_7_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i35_LC_0_7_6  (
            .in0(N__13600),
            .in1(N__10093),
            .in2(N__10388),
            .in3(N__14012),
            .lcout(\tok.C_stk.tail_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28473),
            .ce(N__13370),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i43_LC_0_7_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i43_LC_0_7_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i43_LC_0_7_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i43_LC_0_7_7  (
            .in0(N__14009),
            .in1(N__10081),
            .in2(N__10579),
            .in3(N__13604),
            .lcout(\tok.tail_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28473),
            .ce(N__13370),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i0_LC_0_8_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i0_LC_0_8_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i0_LC_0_8_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tok.C_stk.tail_i0_i0_LC_0_8_0  (
            .in0(N__13605),
            .in1(N__14020),
            .in2(N__10187),
            .in3(N__11491),
            .lcout(\tok.C_stk.tail_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28478),
            .ce(N__13329),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i5283_3_lut_LC_0_8_1 .C_ON=1'b0;
    defparam \tok.C_stk.i5283_3_lut_LC_0_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i5283_3_lut_LC_0_8_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i5283_3_lut_LC_0_8_1  (
            .in0(N__10195),
            .in1(N__14251),
            .in2(_gnd_net_),
            .in3(N__12758),
            .lcout(),
            .ltout(\tok.C_stk.n5456_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i0_LC_0_8_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i0_LC_0_8_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i0_LC_0_8_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i0_LC_0_8_2  (
            .in0(N__14197),
            .in1(N__15544),
            .in2(N__10202),
            .in3(N__12785),
            .lcout(\tok.c_stk_r_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28478),
            .ce(N__13329),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i8_LC_0_8_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i8_LC_0_8_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i8_LC_0_8_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i8_LC_0_8_3  (
            .in0(N__14019),
            .in1(N__10171),
            .in2(N__10199),
            .in3(N__13610),
            .lcout(\tok.tail_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28478),
            .ce(N__13329),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i16_LC_0_8_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i16_LC_0_8_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i16_LC_0_8_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i16_LC_0_8_4  (
            .in0(N__13606),
            .in1(N__10154),
            .in2(N__10186),
            .in3(N__14021),
            .lcout(\tok.C_stk.tail_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28478),
            .ce(N__13329),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i24_LC_0_8_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i24_LC_0_8_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i24_LC_0_8_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i24_LC_0_8_5  (
            .in0(N__14017),
            .in1(N__10145),
            .in2(N__10172),
            .in3(N__13608),
            .lcout(\tok.tail_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28478),
            .ce(N__13329),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i32_LC_0_8_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i32_LC_0_8_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i32_LC_0_8_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i32_LC_0_8_6  (
            .in0(N__13607),
            .in1(N__10153),
            .in2(N__10343),
            .in3(N__14022),
            .lcout(\tok.C_stk.tail_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28478),
            .ce(N__13329),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i40_LC_0_8_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i40_LC_0_8_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i40_LC_0_8_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i40_LC_0_8_7  (
            .in0(N__14018),
            .in1(N__10144),
            .in2(N__10475),
            .in3(N__13609),
            .lcout(\tok.tail_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28478),
            .ce(N__13329),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i52_LC_0_9_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i52_LC_0_9_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i52_LC_0_9_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i52_LC_0_9_7  (
            .in0(N__14038),
            .in1(N__10723),
            .in2(N__10595),
            .in3(N__13694),
            .lcout(\tok.tail_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28483),
            .ce(N__13371),
            .sr(_gnd_net_));
    defparam \tok.uart.rxclkcounter_148__i0_LC_1_3_0 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_148__i0_LC_1_3_0 .SEQ_MODE=4'b1001;
    defparam \tok.uart.rxclkcounter_148__i0_LC_1_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_148__i0_LC_1_3_0  (
            .in0(_gnd_net_),
            .in1(N__10850),
            .in2(_gnd_net_),
            .in3(N__10136),
            .lcout(\tok.uart.rxclkcounter_0 ),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\tok.uart.n4827 ),
            .clk(N__28466),
            .ce(),
            .sr(N__11279));
    defparam \tok.uart.rxclkcounter_148__i1_LC_1_3_1 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_148__i1_LC_1_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_148__i1_LC_1_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_148__i1_LC_1_3_1  (
            .in0(_gnd_net_),
            .in1(N__10823),
            .in2(_gnd_net_),
            .in3(N__10229),
            .lcout(\tok.uart.rxclkcounter_1 ),
            .ltout(),
            .carryin(\tok.uart.n4827 ),
            .carryout(\tok.uart.n4828 ),
            .clk(N__28466),
            .ce(),
            .sr(N__11279));
    defparam \tok.uart.rxclkcounter_148__i2_LC_1_3_2 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_148__i2_LC_1_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_148__i2_LC_1_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_148__i2_LC_1_3_2  (
            .in0(_gnd_net_),
            .in1(N__10894),
            .in2(_gnd_net_),
            .in3(N__10226),
            .lcout(\tok.uart.rxclkcounter_2 ),
            .ltout(),
            .carryin(\tok.uart.n4828 ),
            .carryout(\tok.uart.n4829 ),
            .clk(N__28466),
            .ce(),
            .sr(N__11279));
    defparam \tok.uart.rxclkcounter_148__i3_LC_1_3_3 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_148__i3_LC_1_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_148__i3_LC_1_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_148__i3_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__10907),
            .in2(_gnd_net_),
            .in3(N__10223),
            .lcout(\tok.uart.rxclkcounter_3 ),
            .ltout(),
            .carryin(\tok.uart.n4829 ),
            .carryout(\tok.uart.n4830 ),
            .clk(N__28466),
            .ce(),
            .sr(N__11279));
    defparam \tok.uart.rxclkcounter_148__i4_LC_1_3_4 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_148__i4_LC_1_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_148__i4_LC_1_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_148__i4_LC_1_3_4  (
            .in0(_gnd_net_),
            .in1(N__10837),
            .in2(_gnd_net_),
            .in3(N__10220),
            .lcout(\tok.uart.rxclkcounter_4 ),
            .ltout(),
            .carryin(\tok.uart.n4830 ),
            .carryout(\tok.uart.n4831 ),
            .clk(N__28466),
            .ce(),
            .sr(N__11279));
    defparam \tok.uart.rxclkcounter_148__i5_LC_1_3_5 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_148__i5_LC_1_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_148__i5_LC_1_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_148__i5_LC_1_3_5  (
            .in0(_gnd_net_),
            .in1(N__10919),
            .in2(_gnd_net_),
            .in3(N__10217),
            .lcout(\tok.uart.rxclkcounter_5 ),
            .ltout(),
            .carryin(\tok.uart.n4831 ),
            .carryout(\tok.uart.n4832 ),
            .clk(N__28466),
            .ce(),
            .sr(N__11279));
    defparam \tok.uart.rxclkcounter_148__i6_LC_1_3_6 .C_ON=1'b0;
    defparam \tok.uart.rxclkcounter_148__i6_LC_1_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_148__i6_LC_1_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_148__i6_LC_1_3_6  (
            .in0(_gnd_net_),
            .in1(N__10862),
            .in2(_gnd_net_),
            .in3(N__10214),
            .lcout(\tok.uart.rxclkcounter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28466),
            .ce(),
            .sr(N__11279));
    defparam \tok.uart.txclkcounter_145__i0_LC_1_4_0 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_145__i0_LC_1_4_0 .SEQ_MODE=4'b1001;
    defparam \tok.uart.txclkcounter_145__i0_LC_1_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_145__i0_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(N__10979),
            .in2(_gnd_net_),
            .in3(N__10211),
            .lcout(\tok.uart.txclkcounter_0 ),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(\tok.uart.n4814 ),
            .clk(N__28468),
            .ce(),
            .sr(N__11793));
    defparam \tok.uart.txclkcounter_145__i1_LC_1_4_1 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_145__i1_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_145__i1_LC_1_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_145__i1_LC_1_4_1  (
            .in0(_gnd_net_),
            .in1(N__10967),
            .in2(_gnd_net_),
            .in3(N__10208),
            .lcout(\tok.uart.txclkcounter_1 ),
            .ltout(),
            .carryin(\tok.uart.n4814 ),
            .carryout(\tok.uart.n4815 ),
            .clk(N__28468),
            .ce(),
            .sr(N__11793));
    defparam \tok.uart.txclkcounter_145__i2_LC_1_4_2 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_145__i2_LC_1_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_145__i2_LC_1_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_145__i2_LC_1_4_2  (
            .in0(_gnd_net_),
            .in1(N__11069),
            .in2(_gnd_net_),
            .in3(N__10205),
            .lcout(\tok.uart.txclkcounter_2 ),
            .ltout(),
            .carryin(\tok.uart.n4815 ),
            .carryout(\tok.uart.n4816 ),
            .clk(N__28468),
            .ce(),
            .sr(N__11793));
    defparam \tok.uart.txclkcounter_145__i3_LC_1_4_3 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_145__i3_LC_1_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_145__i3_LC_1_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_145__i3_LC_1_4_3  (
            .in0(_gnd_net_),
            .in1(N__11042),
            .in2(_gnd_net_),
            .in3(N__10250),
            .lcout(\tok.uart.txclkcounter_3 ),
            .ltout(),
            .carryin(\tok.uart.n4816 ),
            .carryout(\tok.uart.n4817 ),
            .clk(N__28468),
            .ce(),
            .sr(N__11793));
    defparam \tok.uart.txclkcounter_145__i4_LC_1_4_4 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_145__i4_LC_1_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_145__i4_LC_1_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_145__i4_LC_1_4_4  (
            .in0(_gnd_net_),
            .in1(N__11015),
            .in2(_gnd_net_),
            .in3(N__10247),
            .lcout(\tok.uart.txclkcounter_4 ),
            .ltout(),
            .carryin(\tok.uart.n4817 ),
            .carryout(\tok.uart.n4818 ),
            .clk(N__28468),
            .ce(),
            .sr(N__11793));
    defparam \tok.uart.txclkcounter_145__i5_LC_1_4_5 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_145__i5_LC_1_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_145__i5_LC_1_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_145__i5_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(N__11083),
            .in2(_gnd_net_),
            .in3(N__10244),
            .lcout(\tok.uart.txclkcounter_5 ),
            .ltout(),
            .carryin(\tok.uart.n4818 ),
            .carryout(\tok.uart.n4819 ),
            .clk(N__28468),
            .ce(),
            .sr(N__11793));
    defparam \tok.uart.txclkcounter_145__i6_LC_1_4_6 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_145__i6_LC_1_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_145__i6_LC_1_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_145__i6_LC_1_4_6  (
            .in0(_gnd_net_),
            .in1(N__10991),
            .in2(_gnd_net_),
            .in3(N__10241),
            .lcout(\tok.uart.txclkcounter_6 ),
            .ltout(),
            .carryin(\tok.uart.n4819 ),
            .carryout(\tok.uart.n4820 ),
            .clk(N__28468),
            .ce(),
            .sr(N__11793));
    defparam \tok.uart.txclkcounter_145__i7_LC_1_4_7 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_145__i7_LC_1_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_145__i7_LC_1_4_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_145__i7_LC_1_4_7  (
            .in0(_gnd_net_),
            .in1(N__11003),
            .in2(_gnd_net_),
            .in3(N__10238),
            .lcout(\tok.uart.txclkcounter_7 ),
            .ltout(),
            .carryin(\tok.uart.n4820 ),
            .carryout(\tok.uart.n4821 ),
            .clk(N__28468),
            .ce(),
            .sr(N__11793));
    defparam \tok.uart.txclkcounter_145__i8_LC_1_5_0 .C_ON=1'b0;
    defparam \tok.uart.txclkcounter_145__i8_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_145__i8_LC_1_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_145__i8_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(N__11056),
            .in2(_gnd_net_),
            .in3(N__10235),
            .lcout(\tok.uart.txclkcounter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28470),
            .ce(),
            .sr(N__11794));
    defparam \tok.C_stk.tail_i0_i1_LC_1_6_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i1_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i1_LC_1_6_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \tok.C_stk.tail_i0_i1_LC_1_6_0  (
            .in0(N__10312),
            .in1(N__13899),
            .in2(N__13692),
            .in3(N__12611),
            .lcout(\tok.C_stk.tail_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28474),
            .ce(N__13345),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i5280_3_lut_LC_1_6_1 .C_ON=1'b0;
    defparam \tok.C_stk.i5280_3_lut_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i5280_3_lut_LC_1_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i5280_3_lut_LC_1_6_1  (
            .in0(N__10324),
            .in1(N__14269),
            .in2(_gnd_net_),
            .in3(N__12716),
            .lcout(),
            .ltout(\tok.C_stk.n5453_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i1_LC_1_6_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i1_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i1_LC_1_6_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i1_LC_1_6_2  (
            .in0(N__14164),
            .in1(N__15545),
            .in2(N__10232),
            .in3(N__15731),
            .lcout(\tok.c_stk_r_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28474),
            .ce(N__13345),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i9_LC_1_6_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i9_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i9_LC_1_6_3 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.C_stk.tail_i0_i9_LC_1_6_3  (
            .in0(N__13898),
            .in1(N__10301),
            .in2(N__13690),
            .in3(N__10325),
            .lcout(\tok.tail_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28474),
            .ce(N__13345),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i17_LC_1_6_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i17_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i17_LC_1_6_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i17_LC_1_6_4  (
            .in0(N__10292),
            .in1(N__13611),
            .in2(N__10313),
            .in3(N__13900),
            .lcout(\tok.C_stk.tail_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28474),
            .ce(N__13345),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i25_LC_1_6_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i25_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i25_LC_1_6_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.C_stk.tail_i0_i25_LC_1_6_5  (
            .in0(N__13896),
            .in1(N__10300),
            .in2(N__13688),
            .in3(N__10283),
            .lcout(\tok.tail_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28474),
            .ce(N__13345),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i33_LC_1_6_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i33_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i33_LC_1_6_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i33_LC_1_6_6  (
            .in0(N__10291),
            .in1(N__13612),
            .in2(N__10361),
            .in3(N__13901),
            .lcout(\tok.C_stk.tail_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28474),
            .ce(N__13345),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i41_LC_1_6_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i41_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i41_LC_1_6_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.C_stk.tail_i0_i41_LC_1_6_7  (
            .in0(N__13897),
            .in1(N__10511),
            .in2(N__13689),
            .in3(N__10282),
            .lcout(\tok.tail_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28474),
            .ce(N__13345),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i2_LC_1_7_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i2_LC_1_7_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i2_LC_1_7_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.C_stk.tail_i0_i2_LC_1_7_0  (
            .in0(N__14001),
            .in1(N__11131),
            .in2(N__13691),
            .in3(N__10259),
            .lcout(\tok.C_stk.tail_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28479),
            .ce(N__13361),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i5277_3_lut_LC_1_7_1 .C_ON=1'b0;
    defparam \tok.C_stk.i5277_3_lut_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i5277_3_lut_LC_1_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.C_stk.i5277_3_lut_LC_1_7_1  (
            .in0(N__14260),
            .in1(N__10270),
            .in2(_gnd_net_),
            .in3(N__12659),
            .lcout(),
            .ltout(\tok.C_stk.n5450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i2_LC_1_7_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i2_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i2_LC_1_7_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i2_LC_1_7_2  (
            .in0(N__14187),
            .in1(N__15542),
            .in2(N__10274),
            .in3(N__12682),
            .lcout(\tok.c_stk_r_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28479),
            .ce(N__13361),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i10_LC_1_7_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i10_LC_1_7_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i10_LC_1_7_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i10_LC_1_7_3  (
            .in0(N__10271),
            .in1(N__13622),
            .in2(N__10427),
            .in3(N__14003),
            .lcout(\tok.tail_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28479),
            .ce(N__13361),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i18_LC_1_7_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i18_LC_1_7_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i18_LC_1_7_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i18_LC_1_7_4  (
            .in0(N__14000),
            .in1(N__10258),
            .in2(N__10412),
            .in3(N__13631),
            .lcout(\tok.C_stk.tail_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28479),
            .ce(N__13361),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i26_LC_1_7_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i26_LC_1_7_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i26_LC_1_7_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i26_LC_1_7_5  (
            .in0(N__10397),
            .in1(N__13623),
            .in2(N__10426),
            .in3(N__14004),
            .lcout(\tok.tail_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28479),
            .ce(N__13361),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i34_LC_1_7_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i34_LC_1_7_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i34_LC_1_7_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i34_LC_1_7_6  (
            .in0(N__14002),
            .in1(N__10373),
            .in2(N__10411),
            .in3(N__13632),
            .lcout(\tok.C_stk.tail_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28479),
            .ce(N__13361),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i42_LC_1_7_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i42_LC_1_7_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i42_LC_1_7_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i42_LC_1_7_7  (
            .in0(N__10396),
            .in1(N__13627),
            .in2(N__10544),
            .in3(N__14005),
            .lcout(\tok.tail_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28479),
            .ce(N__13361),
            .sr(_gnd_net_));
    defparam \tok.i2454_2_lut_LC_1_8_1 .C_ON=1'b0;
    defparam \tok.i2454_2_lut_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2454_2_lut_LC_1_8_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \tok.i2454_2_lut_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(N__13549),
            .in2(_gnd_net_),
            .in3(N__13902),
            .lcout(\tok.C_stk_delta_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i51_LC_1_8_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i51_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i51_LC_1_8_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i51_LC_1_8_2  (
            .in0(N__13904),
            .in1(N__10384),
            .in2(N__10559),
            .in3(N__13634),
            .lcout(\tok.tail_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28484),
            .ce(N__13328),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i50_LC_1_8_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i50_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i50_LC_1_8_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i50_LC_1_8_3  (
            .in0(N__10372),
            .in1(N__13551),
            .in2(N__10526),
            .in3(N__13907),
            .lcout(\tok.tail_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28484),
            .ce(N__13328),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i49_LC_1_8_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i49_LC_1_8_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i49_LC_1_8_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i49_LC_1_8_4  (
            .in0(N__13903),
            .in1(N__10360),
            .in2(N__10493),
            .in3(N__13633),
            .lcout(\tok.tail_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28484),
            .ce(N__13328),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i48_LC_1_8_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i48_LC_1_8_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i48_LC_1_8_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i48_LC_1_8_5  (
            .in0(N__10342),
            .in1(N__13550),
            .in2(N__10454),
            .in3(N__13906),
            .lcout(\tok.tail_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28484),
            .ce(N__13328),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i55_LC_1_8_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i55_LC_1_8_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i55_LC_1_8_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i55_LC_1_8_6  (
            .in0(N__13905),
            .in1(N__10439),
            .in2(N__10613),
            .in3(N__13635),
            .lcout(\tok.tail_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28484),
            .ce(N__13328),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i60_LC_1_9_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i60_LC_1_9_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i60_LC_1_9_0 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.C_stk.tail_i0_i60_LC_1_9_0  (
            .in0(N__10591),
            .in1(N__13683),
            .in2(N__10744),
            .in3(N__14040),
            .lcout(\tok.tail_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i59_LC_1_9_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i59_LC_1_9_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i59_LC_1_9_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \tok.C_stk.tail_i0_i59_LC_1_9_1  (
            .in0(N__13977),
            .in1(N__10555),
            .in2(N__10580),
            .in3(N__13685),
            .lcout(\tok.tail_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i58_LC_1_9_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i58_LC_1_9_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i58_LC_1_9_2 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \tok.C_stk.tail_i0_i58_LC_1_9_2  (
            .in0(N__10522),
            .in1(N__13682),
            .in2(N__14045),
            .in3(N__10540),
            .lcout(\tok.tail_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i57_LC_1_9_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i57_LC_1_9_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i57_LC_1_9_3 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \tok.C_stk.tail_i0_i57_LC_1_9_3  (
            .in0(N__13976),
            .in1(N__10486),
            .in2(N__10510),
            .in3(N__13684),
            .lcout(\tok.tail_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i56_LC_1_9_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i56_LC_1_9_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i56_LC_1_9_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.C_stk.tail_i0_i56_LC_1_9_4  (
            .in0(N__10450),
            .in1(N__13681),
            .in2(N__10474),
            .in3(N__14039),
            .lcout(\tok.tail_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i63_LC_1_9_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i63_LC_1_9_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i63_LC_1_9_5 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \tok.C_stk.tail_i0_i63_LC_1_9_5  (
            .in0(N__13979),
            .in1(N__10438),
            .in2(N__10633),
            .in3(N__13687),
            .lcout(\tok.tail_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i547_4_lut_LC_1_9_6 .C_ON=1'b0;
    defparam \tok.C_stk.i547_4_lut_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i547_4_lut_LC_1_9_6 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \tok.C_stk.i547_4_lut_LC_1_9_6  (
            .in0(N__13244),
            .in1(N__17498),
            .in2(N__14195),
            .in3(N__13136),
            .lcout(\tok.C_stk.n602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i61_LC_1_9_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i61_LC_1_9_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i61_LC_1_9_7 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \tok.C_stk.tail_i0_i61_LC_1_9_7  (
            .in0(N__13978),
            .in1(N__10933),
            .in2(N__11435),
            .in3(N__13686),
            .lcout(\tok.tail_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i7_LC_1_10_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i7_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i7_LC_1_10_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.C_stk.tail_i0_i7_LC_1_10_0  (
            .in0(N__14034),
            .in1(N__10676),
            .in2(N__13713),
            .in3(N__11584),
            .lcout(\tok.C_stk.tail_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28496),
            .ce(N__13330),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i5262_3_lut_LC_1_10_1 .C_ON=1'b0;
    defparam \tok.C_stk.i5262_3_lut_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i5262_3_lut_LC_1_10_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.C_stk.i5262_3_lut_LC_1_10_1  (
            .in0(N__14256),
            .in1(N__10687),
            .in2(_gnd_net_),
            .in3(N__12959),
            .lcout(),
            .ltout(\tok.C_stk.n5435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i7_LC_1_10_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i7_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i7_LC_1_10_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.head_i0_i7_LC_1_10_2  (
            .in0(N__14196),
            .in1(N__12983),
            .in2(N__10691),
            .in3(N__15527),
            .lcout(\tok.c_stk_r_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28496),
            .ce(N__13330),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i15_LC_1_10_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i15_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i15_LC_1_10_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i15_LC_1_10_3  (
            .in0(N__10688),
            .in1(N__13669),
            .in2(N__10667),
            .in3(N__14035),
            .lcout(\tok.tail_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28496),
            .ce(N__13330),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i23_LC_1_10_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i23_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i23_LC_1_10_4 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.C_stk.tail_i0_i23_LC_1_10_4  (
            .in0(N__14032),
            .in1(N__10652),
            .in2(N__13711),
            .in3(N__10675),
            .lcout(\tok.C_stk.tail_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28496),
            .ce(N__13330),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i31_LC_1_10_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i31_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i31_LC_1_10_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i31_LC_1_10_5  (
            .in0(N__10643),
            .in1(N__13670),
            .in2(N__10666),
            .in3(N__14036),
            .lcout(\tok.tail_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28496),
            .ce(N__13330),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i39_LC_1_10_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i39_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i39_LC_1_10_6 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.C_stk.tail_i0_i39_LC_1_10_6  (
            .in0(N__14033),
            .in1(N__10609),
            .in2(N__13712),
            .in3(N__10651),
            .lcout(\tok.C_stk.tail_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28496),
            .ce(N__13330),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i47_LC_1_10_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i47_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i47_LC_1_10_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i47_LC_1_10_7  (
            .in0(N__10642),
            .in1(N__13671),
            .in2(N__10634),
            .in3(N__14037),
            .lcout(\tok.tail_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28496),
            .ce(N__13330),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i4_LC_1_11_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i4_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i4_LC_1_11_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.tail_i0_i4_LC_1_11_2  (
            .in0(N__13665),
            .in1(N__14029),
            .in2(N__16071),
            .in3(N__10792),
            .lcout(\tok.C_stk.tail_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28501),
            .ce(N__13360),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i12_LC_1_11_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i12_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i12_LC_1_11_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i12_LC_1_11_3  (
            .in0(N__14026),
            .in1(N__11531),
            .in2(N__10778),
            .in3(N__13666),
            .lcout(\tok.tail_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28501),
            .ce(N__13360),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i20_LC_1_11_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i20_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i20_LC_1_11_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i20_LC_1_11_4  (
            .in0(N__13663),
            .in1(N__10763),
            .in2(N__10796),
            .in3(N__14030),
            .lcout(\tok.C_stk.tail_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28501),
            .ce(N__13360),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i28_LC_1_11_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i28_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i28_LC_1_11_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i28_LC_1_11_5  (
            .in0(N__14027),
            .in1(N__10754),
            .in2(N__10777),
            .in3(N__13667),
            .lcout(\tok.tail_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28501),
            .ce(N__13360),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i36_LC_1_11_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i36_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i36_LC_1_11_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i36_LC_1_11_6  (
            .in0(N__13664),
            .in1(N__10762),
            .in2(N__10724),
            .in3(N__14031),
            .lcout(\tok.C_stk.tail_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28501),
            .ce(N__13360),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i44_LC_1_11_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i44_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i44_LC_1_11_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i44_LC_1_11_7  (
            .in0(N__14028),
            .in1(N__10753),
            .in2(N__10745),
            .in3(N__13668),
            .lcout(\tok.tail_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28501),
            .ce(N__13360),
            .sr(_gnd_net_));
    defparam \tok.uart.bytephase__i0_LC_2_2_0 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i0_LC_2_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i0_LC_2_2_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i0_LC_2_2_0  (
            .in0(_gnd_net_),
            .in1(N__11187),
            .in2(_gnd_net_),
            .in3(N__10706),
            .lcout(\tok.uart.bytephase_0 ),
            .ltout(),
            .carryin(bfn_2_2_0_),
            .carryout(\tok.uart.n4822 ),
            .clk(N__28467),
            .ce(N__10874),
            .sr(N__11222));
    defparam \tok.uart.bytephase__i1_LC_2_2_1 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i1_LC_2_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i1_LC_2_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i1_LC_2_2_1  (
            .in0(_gnd_net_),
            .in1(N__11155),
            .in2(_gnd_net_),
            .in3(N__10703),
            .lcout(\tok.uart.bytephase_1 ),
            .ltout(),
            .carryin(\tok.uart.n4822 ),
            .carryout(\tok.uart.n4823 ),
            .clk(N__28467),
            .ce(N__10874),
            .sr(N__11222));
    defparam \tok.uart.bytephase__i2_LC_2_2_2 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i2_LC_2_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i2_LC_2_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i2_LC_2_2_2  (
            .in0(_gnd_net_),
            .in1(N__11264),
            .in2(_gnd_net_),
            .in3(N__10700),
            .lcout(\tok.uart.bytephase_2 ),
            .ltout(),
            .carryin(\tok.uart.n4823 ),
            .carryout(\tok.uart.n4824 ),
            .clk(N__28467),
            .ce(N__10874),
            .sr(N__11222));
    defparam \tok.uart.bytephase__i3_LC_2_2_3 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i3_LC_2_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i3_LC_2_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i3_LC_2_2_3  (
            .in0(_gnd_net_),
            .in1(N__17067),
            .in2(_gnd_net_),
            .in3(N__10697),
            .lcout(\tok.uart.bytephase_3 ),
            .ltout(),
            .carryin(\tok.uart.n4824 ),
            .carryout(\tok.uart.n4825 ),
            .clk(N__28467),
            .ce(N__10874),
            .sr(N__11222));
    defparam \tok.uart.bytephase__i4_LC_2_2_4 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i4_LC_2_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i4_LC_2_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i4_LC_2_2_4  (
            .in0(_gnd_net_),
            .in1(N__11240),
            .in2(_gnd_net_),
            .in3(N__10694),
            .lcout(\tok.uart.bytephase_4 ),
            .ltout(),
            .carryin(\tok.uart.n4825 ),
            .carryout(\tok.uart.n4826 ),
            .clk(N__28467),
            .ce(N__10874),
            .sr(N__11222));
    defparam \tok.uart.bytephase__i5_LC_2_2_5 .C_ON=1'b0;
    defparam \tok.uart.bytephase__i5_LC_2_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i5_LC_2_2_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i5_LC_2_2_5  (
            .in0(_gnd_net_),
            .in1(N__17097),
            .in2(_gnd_net_),
            .in3(N__10922),
            .lcout(\tok.uart.bytephase_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28467),
            .ce(N__10874),
            .sr(N__11222));
    defparam \tok.uart.i6_4_lut_LC_2_3_0 .C_ON=1'b0;
    defparam \tok.uart.i6_4_lut_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i6_4_lut_LC_2_3_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \tok.uart.i6_4_lut_LC_2_3_0  (
            .in0(N__10918),
            .in1(N__10906),
            .in2(N__10895),
            .in3(N__10811),
            .lcout(n813),
            .ltout(n813_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_2_3_1.C_ON=1'b0;
    defparam i1_2_lut_LC_2_3_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_2_3_1.LUT_INIT=16'b1111111100001111;
    LogicCell40 i1_2_lut_LC_2_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10877),
            .in3(N__11218),
            .lcout(n971),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i10_LC_2_3_4 .C_ON=1'b0;
    defparam \tok.uart.sender_i10_LC_2_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i10_LC_2_3_4 .LUT_INIT=16'b1111111001010100;
    LogicCell40 \tok.uart.sender_i10_LC_2_3_4  (
            .in0(N__14374),
            .in1(N__11791),
            .in2(N__14401),
            .in3(N__22326),
            .lcout(sender_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28469),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i2_LC_2_3_5 .C_ON=1'b0;
    defparam \tok.uart.sender_i2_LC_2_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i2_LC_2_3_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \tok.uart.sender_i2_LC_2_3_5  (
            .in0(N__11792),
            .in1(N__11632),
            .in2(N__13226),
            .in3(N__14373),
            .lcout(sender_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28469),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i127_LC_2_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i127_LC_2_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i127_LC_2_3_6 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \tok.A_stk.tail_i0_i127_LC_2_3_6  (
            .in0(N__16516),
            .in1(N__26057),
            .in2(N__17186),
            .in3(N__26581),
            .lcout(tail_127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28469),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i5_4_lut_adj_27_LC_2_3_7 .C_ON=1'b0;
    defparam \tok.uart.i5_4_lut_adj_27_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5_4_lut_adj_27_LC_2_3_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.uart.i5_4_lut_adj_27_LC_2_3_7  (
            .in0(N__10861),
            .in1(N__10849),
            .in2(N__10838),
            .in3(N__10822),
            .lcout(\tok.uart.n12_adj_640 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i2_4_lut_LC_2_4_0 .C_ON=1'b0;
    defparam \tok.uart.i2_4_lut_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_4_lut_LC_2_4_0 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \tok.uart.i2_4_lut_LC_2_4_0  (
            .in0(N__10804),
            .in1(N__12048),
            .in2(N__11030),
            .in3(N__12021),
            .lcout(\tok.uart_tx_busy ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sentbits_147__i3_LC_2_4_1 .C_ON=1'b0;
    defparam \tok.uart.sentbits_147__i3_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_147__i3_LC_2_4_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \tok.uart.sentbits_147__i3_LC_2_4_1  (
            .in0(N__12023),
            .in1(N__11029),
            .in2(N__12056),
            .in3(N__10805),
            .lcout(\tok.uart.sentbits_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28471),
            .ce(N__11999),
            .sr(N__11981));
    defparam \tok.uart.i5_4_lut_LC_2_4_2 .C_ON=1'b0;
    defparam \tok.uart.i5_4_lut_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5_4_lut_LC_2_4_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.uart.i5_4_lut_LC_2_4_2  (
            .in0(N__11084),
            .in1(N__11068),
            .in2(N__11057),
            .in3(N__11041),
            .lcout(\tok.uart.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sentbits_147__i2_LC_2_4_3 .C_ON=1'b0;
    defparam \tok.uart.sentbits_147__i2_LC_2_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_147__i2_LC_2_4_3 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \tok.uart.sentbits_147__i2_LC_2_4_3  (
            .in0(N__12022),
            .in1(_gnd_net_),
            .in2(N__12055),
            .in3(N__11028),
            .lcout(\tok.uart.sentbits_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28471),
            .ce(N__11999),
            .sr(N__11981));
    defparam \tok.uart.i5246_3_lut_LC_2_4_4 .C_ON=1'b0;
    defparam \tok.uart.i5246_3_lut_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5246_3_lut_LC_2_4_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.uart.i5246_3_lut_LC_2_4_4  (
            .in0(N__11014),
            .in1(N__11002),
            .in2(_gnd_net_),
            .in3(N__10990),
            .lcout(),
            .ltout(\tok.uart.n5418_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i5618_4_lut_LC_2_4_5 .C_ON=1'b0;
    defparam \tok.uart.i5618_4_lut_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5618_4_lut_LC_2_4_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \tok.uart.i5618_4_lut_LC_2_4_5  (
            .in0(N__10978),
            .in1(N__10966),
            .in2(N__10955),
            .in3(N__10952),
            .lcout(txtick),
            .ltout(txtick_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i5612_2_lut_LC_2_4_6 .C_ON=1'b0;
    defparam \tok.uart.i5612_2_lut_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5612_2_lut_LC_2_4_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \tok.uart.i5612_2_lut_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10946),
            .in3(N__14365),
            .lcout(\tok.uart.n1017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i53_LC_2_5_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i53_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i53_LC_2_5_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i53_LC_2_5_0  (
            .in0(N__11407),
            .in1(N__13648),
            .in2(N__10943),
            .in3(N__14006),
            .lcout(\tok.tail_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28475),
            .ce(N__13363),
            .sr(_gnd_net_));
    defparam \tok.ram.i5523_4_lut_LC_2_5_1 .C_ON=1'b0;
    defparam \tok.ram.i5523_4_lut_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5523_4_lut_LC_2_5_1 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.ram.i5523_4_lut_LC_2_5_1  (
            .in0(N__15963),
            .in1(N__12658),
            .in2(N__11135),
            .in3(N__19903),
            .lcout(\tok.ram.n5585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_4_lut_LC_2_5_2 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_4_lut_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_4_lut_LC_2_5_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.uart.i1_2_lut_4_lut_LC_2_5_2  (
            .in0(N__11156),
            .in1(N__11265),
            .in2(N__11204),
            .in3(N__11241),
            .lcout(\tok.uart.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i2_2_lut_3_lut_LC_2_5_3 .C_ON=1'b0;
    defparam \tok.uart.i2_2_lut_3_lut_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_2_lut_3_lut_LC_2_5_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.uart.i2_2_lut_3_lut_LC_2_5_3  (
            .in0(N__11266),
            .in1(N__11159),
            .in2(_gnd_net_),
            .in3(N__11202),
            .lcout(),
            .ltout(\tok.uart.n2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rxrst_I_0_4_lut_LC_2_5_4 .C_ON=1'b0;
    defparam \tok.uart.rxrst_I_0_4_lut_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.uart.rxrst_I_0_4_lut_LC_2_5_4 .LUT_INIT=16'b0101010101011101;
    LogicCell40 \tok.uart.rxrst_I_0_4_lut_LC_2_5_4  (
            .in0(N__11171),
            .in1(N__17123),
            .in2(N__11282),
            .in3(N__11243),
            .lcout(\tok.uart.rxclkcounter_6__N_477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i24_3_lut_4_lut_LC_2_5_5 .C_ON=1'b0;
    defparam \tok.uart.i24_3_lut_4_lut_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i24_3_lut_4_lut_LC_2_5_5 .LUT_INIT=16'b0000010010100000;
    LogicCell40 \tok.uart.i24_3_lut_4_lut_LC_2_5_5  (
            .in0(N__17101),
            .in1(N__17159),
            .in2(N__17078),
            .in3(N__11157),
            .lcout(),
            .ltout(\tok.uart.n13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_3_lut_4_lut_LC_2_5_6 .C_ON=1'b0;
    defparam \tok.uart.i1_3_lut_4_lut_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_3_lut_4_lut_LC_2_5_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \tok.uart.i1_3_lut_4_lut_LC_2_5_6  (
            .in0(N__11201),
            .in1(N__11267),
            .in2(N__11246),
            .in3(N__11242),
            .lcout(bytephase_5__N_510),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i2_3_lut_LC_2_5_7 .C_ON=1'b0;
    defparam \tok.uart.i2_3_lut_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_3_lut_LC_2_5_7 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \tok.uart.i2_3_lut_LC_2_5_7  (
            .in0(N__11203),
            .in1(N__11170),
            .in2(_gnd_net_),
            .in3(N__11158),
            .lcout(n4858),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_LC_2_6_0 .C_ON=1'b0;
    defparam \tok.i125_4_lut_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_LC_2_6_0 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_LC_2_6_0  (
            .in0(N__11126),
            .in1(N__18340),
            .in2(N__17719),
            .in3(N__20292),
            .lcout(\tok.n83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6_4_lut_adj_20_LC_2_6_1 .C_ON=1'b0;
    defparam \tok.ram.i6_4_lut_adj_20_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6_4_lut_adj_20_LC_2_6_1 .LUT_INIT=16'b1100110000001010;
    LogicCell40 \tok.ram.i6_4_lut_adj_20_LC_2_6_1  (
            .in0(N__11130),
            .in1(N__11105),
            .in2(N__15889),
            .in3(N__29997),
            .lcout(),
            .ltout(\tok.n3_adj_645_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_29_LC_2_6_2 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_29_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_29_LC_2_6_2 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \tok.i27_4_lut_adj_29_LC_2_6_2  (
            .in0(N__19236),
            .in1(N__11090),
            .in2(N__11099),
            .in3(N__20295),
            .lcout(\tok.n13_adj_646 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5540_2_lut_3_lut_LC_2_6_3 .C_ON=1'b0;
    defparam \tok.i5540_2_lut_3_lut_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5540_2_lut_3_lut_LC_2_6_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.i5540_2_lut_3_lut_LC_2_6_3  (
            .in0(N__11096),
            .in1(N__19056),
            .in2(_gnd_net_),
            .in3(N__29996),
            .lcout(\tok.n5603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_LC_2_6_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_LC_2_6_4 .LUT_INIT=16'b1011111101111111;
    LogicCell40 \tok.i1_4_lut_4_lut_LC_2_6_4  (
            .in0(N__29995),
            .in1(N__18341),
            .in2(N__19255),
            .in3(N__20294),
            .lcout(\tok.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i59_3_lut_adj_127_LC_2_6_5 .C_ON=1'b0;
    defparam \tok.i59_3_lut_adj_127_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i59_3_lut_adj_127_LC_2_6_5 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \tok.i59_3_lut_adj_127_LC_2_6_5  (
            .in0(N__18339),
            .in1(N__19055),
            .in2(_gnd_net_),
            .in3(N__29994),
            .lcout(),
            .ltout(\tok.n31_adj_795_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i58_4_lut_LC_2_6_6 .C_ON=1'b0;
    defparam \tok.i58_4_lut_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i58_4_lut_LC_2_6_6 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \tok.i58_4_lut_LC_2_6_6  (
            .in0(N__19232),
            .in1(N__11327),
            .in2(N__11330),
            .in3(N__20293),
            .lcout(\tok.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5450_4_lut_LC_2_6_7 .C_ON=1'b0;
    defparam \tok.i5450_4_lut_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.i5450_4_lut_LC_2_6_7 .LUT_INIT=16'b0100100010000000;
    LogicCell40 \tok.i5450_4_lut_LC_2_6_7  (
            .in0(N__20291),
            .in1(N__19054),
            .in2(N__18359),
            .in3(N__29993),
            .lcout(\tok.n5473 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i5_LC_2_7_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i5_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i5_LC_2_7_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.tail_i0_i5_LC_2_7_0  (
            .in0(N__13644),
            .in1(N__13997),
            .in2(N__12128),
            .in3(N__11306),
            .lcout(\tok.C_stk.tail_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28485),
            .ce(N__13372),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i5268_3_lut_LC_2_7_1 .C_ON=1'b0;
    defparam \tok.C_stk.i5268_3_lut_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i5268_3_lut_LC_2_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i5268_3_lut_LC_2_7_1  (
            .in0(N__11314),
            .in1(N__14265),
            .in2(_gnd_net_),
            .in3(N__13022),
            .lcout(),
            .ltout(\tok.C_stk.n5441_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i5_LC_2_7_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i5_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i5_LC_2_7_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i5_LC_2_7_2  (
            .in0(N__14186),
            .in1(N__15528),
            .in2(N__11321),
            .in3(N__13049),
            .lcout(\tok.c_stk_r_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28485),
            .ce(N__13372),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i13_LC_2_7_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i13_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i13_LC_2_7_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i13_LC_2_7_3  (
            .in0(N__13994),
            .in1(N__11296),
            .in2(N__11318),
            .in3(N__13645),
            .lcout(\tok.tail_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28485),
            .ce(N__13372),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i21_LC_2_7_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i21_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i21_LC_2_7_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i21_LC_2_7_4  (
            .in0(N__13642),
            .in1(N__11305),
            .in2(N__11459),
            .in3(N__13998),
            .lcout(\tok.C_stk.tail_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28485),
            .ce(N__13372),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i29_LC_2_7_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i29_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i29_LC_2_7_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i29_LC_2_7_5  (
            .in0(N__13995),
            .in1(N__11444),
            .in2(N__11297),
            .in3(N__13646),
            .lcout(\tok.tail_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28485),
            .ce(N__13372),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i37_LC_2_7_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i37_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i37_LC_2_7_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i37_LC_2_7_6  (
            .in0(N__13643),
            .in1(N__11455),
            .in2(N__11408),
            .in3(N__13999),
            .lcout(\tok.C_stk.tail_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28485),
            .ce(N__13372),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i45_LC_2_7_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i45_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i45_LC_2_7_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i45_LC_2_7_7  (
            .in0(N__13996),
            .in1(N__11443),
            .in2(N__11431),
            .in3(N__13647),
            .lcout(\tok.tail_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28485),
            .ce(N__13372),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_89_LC_2_8_0 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_89_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_89_LC_2_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.i26_3_lut_adj_89_LC_2_8_0  (
            .in0(N__11375),
            .in1(N__16196),
            .in2(_gnd_net_),
            .in3(N__12779),
            .lcout(\tok.tc_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_197_LC_2_8_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_197_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_197_LC_2_8_1 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \tok.i1_4_lut_adj_197_LC_2_8_1  (
            .in0(N__16310),
            .in1(N__12752),
            .in2(N__16382),
            .in3(N__11468),
            .lcout(n92),
            .ltout(n92_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i0_LC_2_8_2 .C_ON=1'b0;
    defparam \tok.tc_i0_LC_2_8_2 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i0_LC_2_8_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \tok.tc_i0_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__16197),
            .in2(N__11369),
            .in3(N__12780),
            .lcout(tc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28489),
            .ce(),
            .sr(N__28238));
    defparam \tok.tc_i3_LC_2_8_3 .C_ON=1'b0;
    defparam \tok.tc_i3_LC_2_8_3 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i3_LC_2_8_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \tok.tc_i3_LC_2_8_3  (
            .in0(N__16201),
            .in1(N__14945),
            .in2(N__13086),
            .in3(_gnd_net_),
            .lcout(tc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28489),
            .ce(),
            .sr(N__28238));
    defparam \tok.i26_3_lut_adj_86_LC_2_8_4 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_86_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_86_LC_2_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.i26_3_lut_adj_86_LC_2_8_4  (
            .in0(N__14944),
            .in1(N__13076),
            .in2(_gnd_net_),
            .in3(N__16194),
            .lcout(\tok.tc_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_32_LC_2_8_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_32_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_32_LC_2_8_5 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \tok.i1_4_lut_adj_32_LC_2_8_5  (
            .in0(N__16311),
            .in1(N__12654),
            .in2(N__16383),
            .in3(N__11354),
            .lcout(n10),
            .ltout(n10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_87_LC_2_8_6 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_87_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_87_LC_2_8_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \tok.i26_3_lut_adj_87_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__16195),
            .in2(N__11345),
            .in3(N__12680),
            .lcout(\tok.tc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i2_LC_2_8_7 .C_ON=1'b0;
    defparam \tok.tc_i2_LC_2_8_7 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i2_LC_2_8_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \tok.tc_i2_LC_2_8_7  (
            .in0(N__12681),
            .in1(_gnd_net_),
            .in2(N__16205),
            .in3(N__11519),
            .lcout(tc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28489),
            .ce(),
            .sr(N__28238));
    defparam \tok.i57_3_lut_3_lut_LC_2_9_1 .C_ON=1'b0;
    defparam \tok.i57_3_lut_3_lut_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i57_3_lut_3_lut_LC_2_9_1 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \tok.i57_3_lut_3_lut_LC_2_9_1  (
            .in0(N__19017),
            .in1(N__18293),
            .in2(_gnd_net_),
            .in3(N__29942),
            .lcout(),
            .ltout(\tok.n36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i59_4_lut_LC_2_9_2 .C_ON=1'b0;
    defparam \tok.i59_4_lut_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i59_4_lut_LC_2_9_2 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \tok.i59_4_lut_LC_2_9_2  (
            .in0(N__20265),
            .in1(N__11540),
            .in2(N__11513),
            .in3(N__19198),
            .lcout(\tok.n42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_194_LC_2_9_3 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_194_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_194_LC_2_9_3 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_194_LC_2_9_3  (
            .in0(N__11499),
            .in1(N__18294),
            .in2(N__17560),
            .in3(N__20266),
            .lcout(),
            .ltout(\tok.n83_adj_842_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5522_2_lut_3_lut_LC_2_9_4 .C_ON=1'b0;
    defparam \tok.i5522_2_lut_3_lut_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5522_2_lut_3_lut_LC_2_9_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \tok.i5522_2_lut_3_lut_LC_2_9_4  (
            .in0(N__29943),
            .in1(_gnd_net_),
            .in2(N__11510),
            .in3(N__19018),
            .lcout(\tok.n5583 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5531_4_lut_LC_2_9_5 .C_ON=1'b0;
    defparam \tok.ram.i5531_4_lut_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5531_4_lut_LC_2_9_5 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.ram.i5531_4_lut_LC_2_9_5  (
            .in0(N__15961),
            .in1(N__12757),
            .in2(N__11504),
            .in3(N__19896),
            .lcout(),
            .ltout(\tok.ram.n5597_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6_4_lut_adj_26_LC_2_9_6 .C_ON=1'b0;
    defparam \tok.ram.i6_4_lut_adj_26_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6_4_lut_adj_26_LC_2_9_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \tok.ram.i6_4_lut_adj_26_LC_2_9_6  (
            .in0(N__29944),
            .in1(N__15875),
            .in2(N__11507),
            .in3(N__11503),
            .lcout(),
            .ltout(\tok.n3_adj_863_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i18_4_lut_adj_196_LC_2_9_7 .C_ON=1'b0;
    defparam \tok.i18_4_lut_adj_196_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i18_4_lut_adj_196_LC_2_9_7 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \tok.i18_4_lut_adj_196_LC_2_9_7  (
            .in0(N__19199),
            .in1(N__11477),
            .in2(N__11471),
            .in3(N__20267),
            .lcout(\tok.n5_adj_864 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_68_LC_2_10_0 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_68_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_68_LC_2_10_0 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_68_LC_2_10_0  (
            .in0(N__11579),
            .in1(N__18295),
            .in2(N__19300),
            .in3(N__20268),
            .lcout(),
            .ltout(\tok.n83_adj_714_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5495_2_lut_3_lut_LC_2_10_1 .C_ON=1'b0;
    defparam \tok.i5495_2_lut_3_lut_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5495_2_lut_3_lut_LC_2_10_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i5495_2_lut_3_lut_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__18924),
            .in2(N__11462),
            .in3(N__29945),
            .lcout(\tok.n5511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_LC_2_10_2 .C_ON=1'b0;
    defparam \tok.i26_3_lut_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_LC_2_10_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.i26_3_lut_LC_2_10_2  (
            .in0(N__12987),
            .in1(N__16202),
            .in2(_gnd_net_),
            .in3(N__11549),
            .lcout(\tok.tc_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5535_4_lut_LC_2_10_3 .C_ON=1'b0;
    defparam \tok.ram.i5535_4_lut_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5535_4_lut_LC_2_10_3 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \tok.ram.i5535_4_lut_LC_2_10_3  (
            .in0(N__15962),
            .in1(N__19902),
            .in2(N__11585),
            .in3(N__12957),
            .lcout(),
            .ltout(\tok.ram.n5600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6_4_lut_adj_25_LC_2_10_4 .C_ON=1'b0;
    defparam \tok.ram.i6_4_lut_adj_25_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6_4_lut_adj_25_LC_2_10_4 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \tok.ram.i6_4_lut_adj_25_LC_2_10_4  (
            .in0(N__29946),
            .in1(N__15890),
            .in2(N__11588),
            .in3(N__11583),
            .lcout(),
            .ltout(\tok.n3_adj_719_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i18_4_lut_adj_70_LC_2_10_5 .C_ON=1'b0;
    defparam \tok.i18_4_lut_adj_70_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i18_4_lut_adj_70_LC_2_10_5 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \tok.i18_4_lut_adj_70_LC_2_10_5  (
            .in0(N__20269),
            .in1(N__11561),
            .in2(N__11555),
            .in3(N__19166),
            .lcout(),
            .ltout(\tok.n5_adj_720_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_77_LC_2_10_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_77_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_77_LC_2_10_6 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \tok.i1_4_lut_adj_77_LC_2_10_6  (
            .in0(N__12958),
            .in1(N__16390),
            .in2(N__11552),
            .in3(N__16312),
            .lcout(n92_adj_869),
            .ltout(n92_adj_869_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i7_LC_2_10_7 .C_ON=1'b0;
    defparam \tok.tc_i7_LC_2_10_7 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i7_LC_2_10_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.tc_i7_LC_2_10_7  (
            .in0(N__16203),
            .in1(_gnd_net_),
            .in2(N__11543),
            .in3(N__12988),
            .lcout(tc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28502),
            .ce(),
            .sr(N__28226));
    defparam \tok.i5492_3_lut_4_lut_LC_2_11_4 .C_ON=1'b0;
    defparam \tok.i5492_3_lut_4_lut_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5492_3_lut_4_lut_LC_2_11_4 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \tok.i5492_3_lut_4_lut_LC_2_11_4  (
            .in0(N__18214),
            .in1(N__20145),
            .in2(N__18963),
            .in3(N__29878),
            .lcout(\tok.n5507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i62_LC_2_11_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i62_LC_2_11_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i62_LC_2_11_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.C_stk.tail_i0_i62_LC_2_11_6  (
            .in0(N__11692),
            .in1(N__13693),
            .in2(N__11672),
            .in3(N__14044),
            .lcout(\tok.tail_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28509),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i5271_3_lut_LC_2_11_7 .C_ON=1'b0;
    defparam \tok.C_stk.i5271_3_lut_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i5271_3_lut_LC_2_11_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i5271_3_lut_LC_2_11_7  (
            .in0(N__11530),
            .in1(N__14255),
            .in2(_gnd_net_),
            .in3(N__16253),
            .lcout(\tok.C_stk.n5444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i30_LC_2_12_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i30_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i30_LC_2_12_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.C_stk.tail_i0_i30_LC_2_12_0  (
            .in0(N__11657),
            .in1(N__13695),
            .in2(N__13397),
            .in3(N__14015),
            .lcout(\tok.tail_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28514),
            .ce(N__13376),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i38_LC_2_12_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i38_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i38_LC_2_12_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.C_stk.tail_i0_i38_LC_2_12_1  (
            .in0(N__14013),
            .in1(N__11648),
            .in2(N__13714),
            .in3(N__13732),
            .lcout(\tok.C_stk.tail_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28514),
            .ce(N__13376),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i54_LC_2_12_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i54_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i54_LC_2_12_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i54_LC_2_12_2  (
            .in0(N__11647),
            .in1(N__13696),
            .in2(N__11699),
            .in3(N__14016),
            .lcout(\tok.tail_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28514),
            .ce(N__13376),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i4_LC_2_12_5 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i4_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i4_LC_2_12_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i4_LC_2_12_5  (
            .in0(N__14204),
            .in1(N__15535),
            .in2(N__11681),
            .in3(N__16105),
            .lcout(\tok.c_stk_r_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28514),
            .ce(N__13376),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i46_LC_2_12_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i46_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i46_LC_2_12_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.C_stk.tail_i0_i46_LC_2_12_7  (
            .in0(N__14014),
            .in1(N__11668),
            .in2(N__13715),
            .in3(N__11656),
            .lcout(\tok.tail_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28514),
            .ce(N__13376),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i1_LC_2_13_0 .C_ON=1'b0;
    defparam \tok.uart.sender_i1_LC_2_13_0 .SEQ_MODE=4'b1001;
    defparam \tok.uart.sender_i1_LC_2_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tok.uart.sender_i1_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11639),
            .lcout(tx_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28522),
            .ce(N__14293),
            .sr(N__14381));
    defparam \tok.A_stk.tail_i0_i17_LC_4_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i17_LC_4_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i17_LC_4_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i17_LC_4_2_0  (
            .in0(N__11744),
            .in1(N__11708),
            .in2(_gnd_net_),
            .in3(N__26553),
            .lcout(\tok.A_stk.tail_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28472),
            .ce(N__26072),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i1_LC_4_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i1_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i1_LC_4_2_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i1_LC_4_2_1  (
            .in0(N__26554),
            .in1(_gnd_net_),
            .in2(N__11609),
            .in3(N__23980),
            .lcout(\tok.A_stk.tail_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28472),
            .ce(N__26072),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i33_LC_4_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i33_LC_4_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i33_LC_4_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i33_LC_4_2_2  (
            .in0(N__11735),
            .in1(N__11605),
            .in2(_gnd_net_),
            .in3(N__26555),
            .lcout(\tok.A_stk.tail_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28472),
            .ce(N__26072),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i49_LC_4_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i49_LC_4_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i49_LC_4_2_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i49_LC_4_2_3  (
            .in0(N__26556),
            .in1(N__11743),
            .in2(_gnd_net_),
            .in3(N__11726),
            .lcout(\tok.A_stk.tail_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28472),
            .ce(N__26072),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i65_LC_4_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i65_LC_4_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i65_LC_4_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i65_LC_4_2_4  (
            .in0(N__11734),
            .in1(N__11717),
            .in2(_gnd_net_),
            .in3(N__26557),
            .lcout(\tok.A_stk.tail_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28472),
            .ce(N__26072),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i81_LC_4_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i81_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i81_LC_4_2_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i81_LC_4_2_5  (
            .in0(N__26558),
            .in1(N__12313),
            .in2(_gnd_net_),
            .in3(N__11725),
            .lcout(\tok.A_stk.tail_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28472),
            .ce(N__26072),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i97_LC_4_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i97_LC_4_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i97_LC_4_2_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i97_LC_4_2_6  (
            .in0(N__12302),
            .in1(N__11716),
            .in2(_gnd_net_),
            .in3(N__26559),
            .lcout(tail_97),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28472),
            .ce(N__26072),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i1_LC_4_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i1_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i1_LC_4_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i1_LC_4_2_7  (
            .in0(N__11707),
            .in1(N__25467),
            .in2(_gnd_net_),
            .in3(N__21142),
            .lcout(\tok.S_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28472),
            .ce(N__26072),
            .sr(_gnd_net_));
    defparam \tok.depth_i1_LC_4_3_0 .C_ON=1'b0;
    defparam \tok.depth_i1_LC_4_3_0 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i1_LC_4_3_0 .LUT_INIT=16'b1001011010101010;
    LogicCell40 \tok.depth_i1_LC_4_3_0  (
            .in0(N__12359),
            .in1(N__12379),
            .in2(N__16497),
            .in3(N__16435),
            .lcout(\tok.n61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28476),
            .ce(),
            .sr(N__28235));
    defparam \tok.i1_2_lut_3_lut_adj_156_LC_4_3_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_156_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_156_LC_4_3_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_156_LC_4_3_1  (
            .in0(N__12355),
            .in1(_gnd_net_),
            .in2(N__16493),
            .in3(N__18833),
            .lcout(\tok.n4_adj_707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_4_lut_adj_167_LC_4_3_2 .C_ON=1'b0;
    defparam \tok.i2_3_lut_4_lut_adj_167_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_4_lut_adj_167_LC_4_3_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.i2_3_lut_4_lut_adj_167_LC_4_3_2  (
            .in0(N__12358),
            .in1(N__22150),
            .in2(N__18058),
            .in3(N__16480),
            .lcout(\tok.n807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_i0_LC_4_3_3 .C_ON=1'b0;
    defparam \tok.depth_i0_LC_4_3_3 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i0_LC_4_3_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \tok.depth_i0_LC_4_3_3  (
            .in0(N__16434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16488),
            .lcout(\tok.n62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28476),
            .ce(),
            .sr(N__28235));
    defparam \tok.i1_2_lut_adj_147_LC_4_3_4 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_147_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_147_LC_4_3_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_147_LC_4_3_4  (
            .in0(_gnd_net_),
            .in1(N__16476),
            .in2(_gnd_net_),
            .in3(N__12354),
            .lcout(\tok.n890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_4_lut_LC_4_3_5 .C_ON=1'b0;
    defparam \tok.i1_2_lut_4_lut_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_4_lut_LC_4_3_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i1_2_lut_4_lut_LC_4_3_5  (
            .in0(N__12353),
            .in1(N__11881),
            .in2(N__16492),
            .in3(N__11843),
            .lcout(\tok.A_stk_delta_1__N_4 ),
            .ltout(\tok.A_stk_delta_1__N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_4_lut_LC_4_3_6 .C_ON=1'b0;
    defparam \tok.i2_4_lut_4_lut_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_4_lut_LC_4_3_6 .LUT_INIT=16'b1001011011001100;
    LogicCell40 \tok.i2_4_lut_4_lut_LC_4_3_6  (
            .in0(N__16484),
            .in1(N__12356),
            .in2(N__11765),
            .in3(N__16433),
            .lcout(),
            .ltout(\tok.depth_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5236_3_lut_LC_4_3_7 .C_ON=1'b0;
    defparam \tok.i5236_3_lut_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \tok.i5236_3_lut_LC_4_3_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \tok.i5236_3_lut_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(N__11861),
            .in2(N__11762),
            .in3(N__11822),
            .lcout(\tok.n5408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_4_lut_LC_4_4_0 .C_ON=1'b0;
    defparam \tok.i2_3_lut_4_lut_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_4_lut_LC_4_4_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \tok.i2_3_lut_4_lut_LC_4_4_0  (
            .in0(N__12419),
            .in1(N__12451),
            .in2(N__19334),
            .in3(N__18053),
            .lcout(\tok.n820 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5173_2_lut_LC_4_4_1 .C_ON=1'b0;
    defparam \tok.i5173_2_lut_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5173_2_lut_LC_4_4_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i5173_2_lut_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(N__11882),
            .in2(_gnd_net_),
            .in3(N__11844),
            .lcout(\tok.n5338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2525_2_lut_3_lut_4_lut_LC_4_4_2 .C_ON=1'b0;
    defparam \tok.i2525_2_lut_3_lut_4_lut_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2525_2_lut_3_lut_4_lut_LC_4_4_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i2525_2_lut_3_lut_4_lut_LC_4_4_2  (
            .in0(N__11845),
            .in1(N__12450),
            .in2(N__11888),
            .in3(N__16944),
            .lcout(\tok.n2585 ),
            .ltout(\tok.n2585_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_4_lut_LC_4_4_3 .C_ON=1'b0;
    defparam \tok.i3_3_lut_4_lut_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_4_lut_LC_4_4_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \tok.i3_3_lut_4_lut_LC_4_4_3  (
            .in0(N__18054),
            .in1(N__11759),
            .in2(N__11747),
            .in3(N__19333),
            .lcout(\tok.n29_adj_787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_i3_LC_4_4_4 .C_ON=1'b0;
    defparam \tok.depth_i3_LC_4_4_4 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i3_LC_4_4_4 .LUT_INIT=16'b1101101100100100;
    LogicCell40 \tok.depth_i3_LC_4_4_4  (
            .in0(N__12329),
            .in1(N__12467),
            .in2(N__11855),
            .in3(N__11887),
            .lcout(\tok.n59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28480),
            .ce(),
            .sr(N__28236));
    defparam \tok.depth_i2_LC_4_4_5 .C_ON=1'b0;
    defparam \tok.depth_i2_LC_4_4_5 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i2_LC_4_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \tok.depth_i2_LC_4_4_5  (
            .in0(N__12466),
            .in1(N__11853),
            .in2(_gnd_net_),
            .in3(N__12328),
            .lcout(\tok.n60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28480),
            .ce(),
            .sr(N__28236));
    defparam \tok.i2_4_lut_adj_139_LC_4_4_6 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_139_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_139_LC_4_4_6 .LUT_INIT=16'b1101101100100100;
    LogicCell40 \tok.i2_4_lut_adj_139_LC_4_4_6  (
            .in0(N__12327),
            .in1(N__12465),
            .in2(N__11854),
            .in3(N__11886),
            .lcout(\tok.depth_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_134_LC_4_4_7 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_134_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_134_LC_4_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \tok.i2_3_lut_adj_134_LC_4_4_7  (
            .in0(N__12464),
            .in1(N__11846),
            .in2(_gnd_net_),
            .in3(N__12326),
            .lcout(\tok.depth_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_48_LC_4_5_0 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_48_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_48_LC_4_5_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i3_4_lut_adj_48_LC_4_5_0  (
            .in0(N__12420),
            .in1(N__11903),
            .in2(N__11816),
            .in3(N__18306),
            .lcout(\tok.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_220_i9_2_lut_LC_4_5_1 .C_ON=1'b0;
    defparam \tok.T_7__I_0_220_i9_2_lut_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_220_i9_2_lut_LC_4_5_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \tok.T_7__I_0_220_i9_2_lut_LC_4_5_1  (
            .in0(N__18305),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20228),
            .lcout(\tok.n9_adj_766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i5605_4_lut_LC_4_5_2 .C_ON=1'b0;
    defparam \tok.uart.i5605_4_lut_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5605_4_lut_LC_4_5_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \tok.uart.i5605_4_lut_LC_4_5_2  (
            .in0(N__11894),
            .in1(N__18051),
            .in2(N__17812),
            .in3(N__18307),
            .lcout(n23),
            .ltout(n23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i5610_2_lut_3_lut_LC_4_5_3 .C_ON=1'b0;
    defparam \tok.uart.i5610_2_lut_3_lut_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5610_2_lut_3_lut_LC_4_5_3 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \tok.uart.i5610_2_lut_3_lut_LC_4_5_3  (
            .in0(N__11800),
            .in1(_gnd_net_),
            .in2(N__11804),
            .in3(N__17807),
            .lcout(\tok.uart.n1093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_119_i9_2_lut_LC_4_5_4 .C_ON=1'b0;
    defparam \tok.equal_119_i9_2_lut_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.equal_119_i9_2_lut_LC_4_5_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.equal_119_i9_2_lut_LC_4_5_4  (
            .in0(N__20227),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18304),
            .lcout(\tok.n9_adj_798 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_3_lut_LC_4_5_5 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_3_lut_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_3_lut_LC_4_5_5 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \tok.uart.i1_2_lut_3_lut_LC_4_5_5  (
            .in0(N__11801),
            .in1(N__17808),
            .in2(_gnd_net_),
            .in3(N__14332),
            .lcout(\tok.uart.n1023 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sentbits_147__i0_LC_4_5_6 .C_ON=1'b0;
    defparam \tok.uart.sentbits_147__i0_LC_4_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_147__i0_LC_4_5_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.uart.sentbits_147__i0_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12039),
            .lcout(\tok.uart.sentbits_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28486),
            .ce(N__11995),
            .sr(N__11980));
    defparam \tok.uart.sentbits_147__i1_LC_4_5_7 .C_ON=1'b0;
    defparam \tok.uart.sentbits_147__i1_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_147__i1_LC_4_5_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \tok.uart.sentbits_147__i1_LC_4_5_7  (
            .in0(N__12040),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12013),
            .lcout(\tok.uart.sentbits_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28486),
            .ce(N__11995),
            .sr(N__11980));
    defparam \tok.i2_4_lut_adj_64_LC_4_6_0 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_64_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_64_LC_4_6_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \tok.i2_4_lut_adj_64_LC_4_6_0  (
            .in0(N__11930),
            .in1(N__12422),
            .in2(N__11957),
            .in3(N__11942),
            .lcout(\tok.n5298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_119_LC_4_6_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_119_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_119_LC_4_6_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i1_2_lut_adj_119_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(N__22134),
            .in2(_gnd_net_),
            .in3(N__18026),
            .lcout(\tok.n5287 ),
            .ltout(\tok.n5287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_122_LC_4_6_2 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_122_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_122_LC_4_6_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \tok.i5_4_lut_adj_122_LC_4_6_2  (
            .in0(N__12233),
            .in1(N__12278),
            .in2(N__11924),
            .in3(N__16584),
            .lcout(\tok.n241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5149_2_lut_LC_4_6_3 .C_ON=1'b0;
    defparam \tok.i5149_2_lut_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5149_2_lut_LC_4_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i5149_2_lut_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__18835),
            .in2(_gnd_net_),
            .in3(N__18027),
            .lcout(),
            .ltout(\tok.n5312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_124_LC_4_6_4 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_124_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_124_LC_4_6_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \tok.i5_4_lut_adj_124_LC_4_6_4  (
            .in0(N__19060),
            .in1(N__11921),
            .in2(N__11909),
            .in3(N__14930),
            .lcout(\tok.n2515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_143_i15_2_lut_LC_4_6_5 .C_ON=1'b0;
    defparam \tok.equal_143_i15_2_lut_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.equal_143_i15_2_lut_LC_4_6_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \tok.equal_143_i15_2_lut_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__19059),
            .in2(_gnd_net_),
            .in3(N__18834),
            .lcout(),
            .ltout(\tok.n15_adj_817_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i3_4_lut_LC_4_6_6 .C_ON=1'b0;
    defparam \tok.uart.i3_4_lut_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i3_4_lut_LC_4_6_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.uart.i3_4_lut_LC_4_6_6  (
            .in0(N__19239),
            .in1(N__20232),
            .in2(N__11906),
            .in3(N__29984),
            .lcout(\tok.n898 ),
            .ltout(\tok.n898_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_LC_4_6_7 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_LC_4_6_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \tok.uart.i1_2_lut_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11897),
            .in3(N__22135),
            .lcout(\tok.uart.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5546_4_lut_LC_4_7_0 .C_ON=1'b0;
    defparam \tok.ram.i5546_4_lut_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5546_4_lut_LC_4_7_0 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \tok.ram.i5546_4_lut_LC_4_7_0  (
            .in0(N__15953),
            .in1(N__19895),
            .in2(N__12134),
            .in3(N__13013),
            .lcout(),
            .ltout(\tok.ram.n5608_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6_4_lut_adj_23_LC_4_7_1 .C_ON=1'b0;
    defparam \tok.ram.i6_4_lut_adj_23_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6_4_lut_adj_23_LC_4_7_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.ram.i6_4_lut_adj_23_LC_4_7_1  (
            .in0(N__15861),
            .in1(N__12132),
            .in2(N__12137),
            .in3(N__29985),
            .lcout(\tok.n3_adj_683 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_45_LC_4_7_2 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_45_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_45_LC_4_7_2 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_45_LC_4_7_2  (
            .in0(N__12133),
            .in1(N__18313),
            .in2(N__27106),
            .in3(N__20238),
            .lcout(),
            .ltout(\tok.n83_adj_678_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5458_2_lut_3_lut_LC_4_7_3 .C_ON=1'b0;
    defparam \tok.i5458_2_lut_3_lut_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5458_2_lut_3_lut_LC_4_7_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i5458_2_lut_3_lut_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(N__19038),
            .in2(N__12104),
            .in3(N__29986),
            .lcout(),
            .ltout(\tok.n5483_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i18_4_lut_LC_4_7_4 .C_ON=1'b0;
    defparam \tok.i18_4_lut_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i18_4_lut_LC_4_7_4 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \tok.i18_4_lut_LC_4_7_4  (
            .in0(N__12101),
            .in1(N__19240),
            .in2(N__12095),
            .in3(N__20239),
            .lcout(),
            .ltout(\tok.n5_adj_684_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_49_LC_4_7_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_49_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_49_LC_4_7_5 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \tok.i1_4_lut_adj_49_LC_4_7_5  (
            .in0(N__13014),
            .in1(N__16293),
            .in2(N__12092),
            .in3(N__16369),
            .lcout(n92_adj_868),
            .ltout(n92_adj_868_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_83_LC_4_7_6 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_83_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_83_LC_4_7_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \tok.i26_3_lut_adj_83_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(N__16171),
            .in2(N__12089),
            .in3(N__13041),
            .lcout(\tok.tc_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i5_LC_4_7_7 .C_ON=1'b0;
    defparam \tok.tc_i5_LC_4_7_7 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i5_LC_4_7_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.tc_i5_LC_4_7_7  (
            .in0(N__16172),
            .in1(_gnd_net_),
            .in2(N__13048),
            .in3(N__12071),
            .lcout(tc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28497),
            .ce(),
            .sr(N__28212));
    defparam \tok.i1546_3_lut_4_lut_LC_4_8_0 .C_ON=1'b0;
    defparam \tok.i1546_3_lut_4_lut_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1546_3_lut_4_lut_LC_4_8_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \tok.i1546_3_lut_4_lut_LC_4_8_0  (
            .in0(N__23793),
            .in1(N__16242),
            .in2(N__22541),
            .in3(N__15619),
            .lcout(\tok.table_wr_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2569_2_lut_3_lut_LC_4_8_1 .C_ON=1'b0;
    defparam \tok.i2569_2_lut_3_lut_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2569_2_lut_3_lut_LC_4_8_1 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \tok.i2569_2_lut_3_lut_LC_4_8_1  (
            .in0(N__15625),
            .in1(_gnd_net_),
            .in2(N__24782),
            .in3(N__22502),
            .lcout(\tok.table_wr_data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2570_2_lut_3_lut_LC_4_8_2 .C_ON=1'b0;
    defparam \tok.i2570_2_lut_3_lut_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2570_2_lut_3_lut_LC_4_8_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \tok.i2570_2_lut_3_lut_LC_4_8_2  (
            .in0(N__22501),
            .in1(N__28867),
            .in2(_gnd_net_),
            .in3(N__15626),
            .lcout(\tok.table_wr_data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1584_3_lut_4_lut_LC_4_8_3 .C_ON=1'b0;
    defparam \tok.i1584_3_lut_4_lut_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1584_3_lut_4_lut_LC_4_8_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \tok.i1584_3_lut_4_lut_LC_4_8_3  (
            .in0(N__15620),
            .in1(N__22492),
            .in2(N__25375),
            .in3(N__14967),
            .lcout(\tok.table_wr_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1622_3_lut_4_lut_LC_4_8_4 .C_ON=1'b0;
    defparam \tok.i1622_3_lut_4_lut_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1622_3_lut_4_lut_LC_4_8_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \tok.i1622_3_lut_4_lut_LC_4_8_4  (
            .in0(N__23932),
            .in1(N__12650),
            .in2(N__22540),
            .in3(N__15621),
            .lcout(\tok.table_wr_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1660_3_lut_4_lut_LC_4_8_5 .C_ON=1'b0;
    defparam \tok.i1660_3_lut_4_lut_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1660_3_lut_4_lut_LC_4_8_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \tok.i1660_3_lut_4_lut_LC_4_8_5  (
            .in0(N__15622),
            .in1(N__22496),
            .in2(N__24028),
            .in3(N__12710),
            .lcout(\tok.table_wr_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1812_3_lut_4_lut_LC_4_8_6 .C_ON=1'b0;
    defparam \tok.i1812_3_lut_4_lut_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1812_3_lut_4_lut_LC_4_8_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \tok.i1812_3_lut_4_lut_LC_4_8_6  (
            .in0(N__27213),
            .in1(N__13018),
            .in2(N__22542),
            .in3(N__15624),
            .lcout(\tok.table_wr_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1736_3_lut_4_lut_LC_4_8_7 .C_ON=1'b0;
    defparam \tok.i1736_3_lut_4_lut_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1736_3_lut_4_lut_LC_4_8_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \tok.i1736_3_lut_4_lut_LC_4_8_7  (
            .in0(N__15623),
            .in1(N__22497),
            .in2(N__23553),
            .in3(N__12948),
            .lcout(\tok.table_wr_data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2445_2_lut_3_lut_4_lut_LC_4_9_0 .C_ON=1'b0;
    defparam \tok.i2445_2_lut_3_lut_4_lut_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2445_2_lut_3_lut_4_lut_LC_4_9_0 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \tok.i2445_2_lut_3_lut_4_lut_LC_4_9_0  (
            .in0(N__22504),
            .in1(N__24351),
            .in2(N__15672),
            .in3(N__12923),
            .lcout(\tok.table_wr_data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2446_2_lut_3_lut_4_lut_LC_4_9_1 .C_ON=1'b0;
    defparam \tok.i2446_2_lut_3_lut_4_lut_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2446_2_lut_3_lut_4_lut_LC_4_9_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \tok.i2446_2_lut_3_lut_4_lut_LC_4_9_1  (
            .in0(N__12925),
            .in1(N__15663),
            .in2(N__24488),
            .in3(N__22507),
            .lcout(\tok.table_wr_data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2453_2_lut_3_lut_4_lut_LC_4_9_2 .C_ON=1'b0;
    defparam \tok.i2453_2_lut_3_lut_4_lut_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2453_2_lut_3_lut_4_lut_LC_4_9_2 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \tok.i2453_2_lut_3_lut_4_lut_LC_4_9_2  (
            .in0(N__22505),
            .in1(N__25060),
            .in2(N__15673),
            .in3(N__12924),
            .lcout(\tok.table_wr_data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2462_2_lut_3_lut_4_lut_LC_4_9_3 .C_ON=1'b0;
    defparam \tok.i2462_2_lut_3_lut_4_lut_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2462_2_lut_3_lut_4_lut_LC_4_9_3 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \tok.i2462_2_lut_3_lut_4_lut_LC_4_9_3  (
            .in0(N__12926),
            .in1(N__15667),
            .in2(N__27464),
            .in3(N__22508),
            .lcout(\tok.table_wr_data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2469_2_lut_3_lut_4_lut_LC_4_9_4 .C_ON=1'b0;
    defparam \tok.i2469_2_lut_3_lut_4_lut_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2469_2_lut_3_lut_4_lut_LC_4_9_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \tok.i2469_2_lut_3_lut_4_lut_LC_4_9_4  (
            .in0(N__22506),
            .in1(N__27538),
            .in2(N__15674),
            .in3(N__12928),
            .lcout(\tok.table_wr_data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2470_2_lut_3_lut_4_lut_LC_4_9_5 .C_ON=1'b0;
    defparam \tok.i2470_2_lut_3_lut_4_lut_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2470_2_lut_3_lut_4_lut_LC_4_9_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \tok.i2470_2_lut_3_lut_4_lut_LC_4_9_5  (
            .in0(N__12927),
            .in1(N__15671),
            .in2(N__28073),
            .in3(N__22509),
            .lcout(\tok.table_wr_data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1698_3_lut_4_lut_LC_4_9_6 .C_ON=1'b0;
    defparam \tok.i1698_3_lut_4_lut_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1698_3_lut_4_lut_LC_4_9_6 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \tok.i1698_3_lut_4_lut_LC_4_9_6  (
            .in0(N__22503),
            .in1(N__22853),
            .in2(N__12756),
            .in3(N__15594),
            .lcout(\tok.table_wr_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_121_LC_4_9_7 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_121_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_121_LC_4_9_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \tok.i2_3_lut_adj_121_LC_4_9_7  (
            .in0(N__18262),
            .in1(N__20231),
            .in2(_gnd_net_),
            .in3(N__29947),
            .lcout(\tok.n8_adj_790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_219_i11_2_lut_4_lut_LC_4_10_0 .C_ON=1'b0;
    defparam \tok.T_7__I_0_219_i11_2_lut_4_lut_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_219_i11_2_lut_4_lut_LC_4_10_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.T_7__I_0_219_i11_2_lut_4_lut_LC_4_10_0  (
            .in0(N__20166),
            .in1(N__17974),
            .in2(N__18315),
            .in3(N__29911),
            .lcout(\tok.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_118_i10_2_lut_LC_4_10_1 .C_ON=1'b0;
    defparam \tok.equal_118_i10_2_lut_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.equal_118_i10_2_lut_LC_4_10_1 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \tok.equal_118_i10_2_lut_LC_4_10_1  (
            .in0(N__29913),
            .in1(_gnd_net_),
            .in2(N__18023),
            .in3(_gnd_net_),
            .lcout(\tok.n10_adj_803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_2_lut_LC_4_10_2 .C_ON=1'b0;
    defparam \tok.i2_2_lut_2_lut_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_2_lut_LC_4_10_2 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \tok.i2_2_lut_2_lut_LC_4_10_2  (
            .in0(N__20162),
            .in1(_gnd_net_),
            .in2(N__18314),
            .in3(_gnd_net_),
            .lcout(\tok.n5318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_4_lut_LC_4_10_3 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_4_lut_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_4_lut_LC_4_10_3 .LUT_INIT=16'b1111101111111101;
    LogicCell40 \tok.i1_3_lut_4_lut_4_lut_LC_4_10_3  (
            .in0(N__29914),
            .in1(N__18258),
            .in2(N__18024),
            .in3(N__20167),
            .lcout(\tok.n5293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_135_i11_2_lut_4_lut_LC_4_10_4 .C_ON=1'b0;
    defparam \tok.equal_135_i11_2_lut_4_lut_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.equal_135_i11_2_lut_4_lut_LC_4_10_4 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \tok.equal_135_i11_2_lut_4_lut_LC_4_10_4  (
            .in0(N__20164),
            .in1(N__17975),
            .in2(N__18316),
            .in3(N__29912),
            .lcout(\tok.n11_adj_694 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_128_LC_4_10_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_128_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_128_LC_4_10_5 .LUT_INIT=16'b0110101111110111;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_128_LC_4_10_5  (
            .in0(N__29910),
            .in1(N__18250),
            .in2(N__18022),
            .in3(N__20165),
            .lcout(\tok.n10_adj_796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_233_i11_2_lut_4_lut_LC_4_10_6 .C_ON=1'b0;
    defparam \tok.T_7__I_0_233_i11_2_lut_4_lut_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_233_i11_2_lut_4_lut_LC_4_10_6 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \tok.T_7__I_0_233_i11_2_lut_4_lut_LC_4_10_6  (
            .in0(N__20168),
            .in1(N__17982),
            .in2(N__18317),
            .in3(N__29915),
            .lcout(\tok.n11_adj_681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_116_i9_2_lut_LC_4_10_7 .C_ON=1'b0;
    defparam \tok.equal_116_i9_2_lut_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.equal_116_i9_2_lut_LC_4_10_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \tok.equal_116_i9_2_lut_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(N__18251),
            .in2(_gnd_net_),
            .in3(N__20163),
            .lcout(\tok.n9_adj_802 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_213_i11_2_lut_4_lut_LC_4_11_0 .C_ON=1'b0;
    defparam \tok.T_7__I_0_213_i11_2_lut_4_lut_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_213_i11_2_lut_4_lut_LC_4_11_0 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \tok.T_7__I_0_213_i11_2_lut_4_lut_LC_4_11_0  (
            .in0(N__20122),
            .in1(N__17934),
            .in2(N__18280),
            .in3(N__29853),
            .lcout(\tok.n11_adj_788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_111_i11_2_lut_4_lut_LC_4_11_1 .C_ON=1'b0;
    defparam \tok.equal_111_i11_2_lut_4_lut_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.equal_111_i11_2_lut_4_lut_LC_4_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.equal_111_i11_2_lut_4_lut_LC_4_11_1  (
            .in0(N__29850),
            .in1(N__18194),
            .in2(N__17997),
            .in3(N__20120),
            .lcout(\tok.n11_adj_680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_122_i11_2_lut_4_lut_LC_4_11_2 .C_ON=1'b0;
    defparam \tok.equal_122_i11_2_lut_4_lut_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.equal_122_i11_2_lut_4_lut_LC_4_11_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.equal_122_i11_2_lut_4_lut_LC_4_11_2  (
            .in0(N__20121),
            .in1(N__17933),
            .in2(N__18279),
            .in3(N__29852),
            .lcout(\tok.n11_adj_706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_237_i11_2_lut_4_lut_LC_4_11_3 .C_ON=1'b0;
    defparam \tok.T_7__I_0_237_i11_2_lut_4_lut_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_237_i11_2_lut_4_lut_LC_4_11_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \tok.T_7__I_0_237_i11_2_lut_4_lut_LC_4_11_3  (
            .in0(N__20119),
            .in1(N__17926),
            .in2(N__29927),
            .in3(N__18193),
            .lcout(\tok.n11_adj_793 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_214_i14_2_lut_3_lut_4_lut_LC_4_11_4 .C_ON=1'b0;
    defparam \tok.T_7__I_0_214_i14_2_lut_3_lut_4_lut_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_214_i14_2_lut_3_lut_4_lut_LC_4_11_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \tok.T_7__I_0_214_i14_2_lut_3_lut_4_lut_LC_4_11_4  (
            .in0(N__18761),
            .in1(N__22063),
            .in2(N__18962),
            .in3(N__19153),
            .lcout(\tok.n14_adj_644 ),
            .ltout(\tok.n14_adj_644_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_154_i16_2_lut_LC_4_11_5 .C_ON=1'b0;
    defparam \tok.equal_154_i16_2_lut_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.equal_154_i16_2_lut_LC_4_11_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \tok.equal_154_i16_2_lut_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12269),
            .in3(N__13129),
            .lcout(\tok.n399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_4_lut_LC_4_11_6 .C_ON=1'b0;
    defparam \tok.i3_4_lut_4_lut_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_4_lut_LC_4_11_6 .LUT_INIT=16'b0111100100110000;
    LogicCell40 \tok.i3_4_lut_4_lut_LC_4_11_6  (
            .in0(N__18192),
            .in1(N__20118),
            .in2(N__17996),
            .in3(N__29851),
            .lcout(\tok.n8_adj_805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_4_lut_adj_142_LC_4_11_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_4_lut_adj_142_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_4_lut_adj_142_LC_4_11_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \tok.i1_2_lut_4_lut_adj_142_LC_4_11_7  (
            .in0(N__29854),
            .in1(N__18201),
            .in2(N__17998),
            .in3(N__20123),
            .lcout(\tok.n26_adj_750 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5256_4_lut_4_lut_LC_4_12_0 .C_ON=1'b0;
    defparam \tok.i5256_4_lut_4_lut_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5256_4_lut_4_lut_LC_4_12_0 .LUT_INIT=16'b1110111111000111;
    LogicCell40 \tok.i5256_4_lut_4_lut_LC_4_12_0  (
            .in0(N__17962),
            .in1(N__20124),
            .in2(N__18281),
            .in3(N__29855),
            .lcout(\tok.n5429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_67_LC_4_12_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_67_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_67_LC_4_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i1_2_lut_adj_67_LC_4_12_1  (
            .in0(N__18908),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18213),
            .lcout(\tok.n4_adj_712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_LC_4_12_2 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_LC_4_12_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.i1_2_lut_3_lut_LC_4_12_2  (
            .in0(N__19154),
            .in1(N__18765),
            .in2(_gnd_net_),
            .in3(N__18909),
            .lcout(\tok.n7_adj_785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_adj_153_LC_4_12_3 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_adj_153_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_adj_153_LC_4_12_3 .LUT_INIT=16'b1111111110000001;
    LogicCell40 \tok.i1_3_lut_4_lut_adj_153_LC_4_12_3  (
            .in0(N__29858),
            .in1(N__18208),
            .in2(N__20194),
            .in3(N__17965),
            .lcout(\tok.n4848 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i12_1_lut_2_lut_4_lut_LC_4_12_4 .C_ON=1'b0;
    defparam \tok.i12_1_lut_2_lut_4_lut_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i12_1_lut_2_lut_4_lut_LC_4_12_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \tok.i12_1_lut_2_lut_4_lut_LC_4_12_4  (
            .in0(N__17966),
            .in1(N__20132),
            .in2(N__18283),
            .in3(N__29860),
            .lcout(\tok.n20_adj_663 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i20_1_lut_2_lut_4_lut_LC_4_12_5 .C_ON=1'b0;
    defparam \tok.i20_1_lut_2_lut_4_lut_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i20_1_lut_2_lut_4_lut_LC_4_12_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \tok.i20_1_lut_2_lut_4_lut_LC_4_12_5  (
            .in0(N__29859),
            .in1(N__18209),
            .in2(N__20195),
            .in3(N__17967),
            .lcout(\tok.n8_adj_792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5220_2_lut_4_lut_4_lut_LC_4_12_6 .C_ON=1'b0;
    defparam \tok.i5220_2_lut_4_lut_4_lut_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5220_2_lut_4_lut_4_lut_LC_4_12_6 .LUT_INIT=16'b1110101111111111;
    LogicCell40 \tok.i5220_2_lut_4_lut_4_lut_LC_4_12_6  (
            .in0(N__17963),
            .in1(N__20125),
            .in2(N__18282),
            .in3(N__29856),
            .lcout(\tok.n5391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2547_2_lut_LC_4_12_7 .C_ON=1'b0;
    defparam \tok.i2547_2_lut_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2547_2_lut_LC_4_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i2547_2_lut_LC_4_12_7  (
            .in0(N__29857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17964),
            .lcout(\tok.n2607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i113_LC_5_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i113_LC_5_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i113_LC_5_2_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \tok.A_stk.tail_i0_i113_LC_5_2_3  (
            .in0(N__26502),
            .in1(N__12298),
            .in2(N__26056),
            .in3(N__12314),
            .lcout(tail_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28477),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i112_LC_5_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i112_LC_5_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i112_LC_5_2_6 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i112_LC_5_2_6  (
            .in0(N__14431),
            .in1(N__26012),
            .in2(N__14459),
            .in3(N__26501),
            .lcout(tail_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28477),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_151_LC_5_3_0 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_151_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_151_LC_5_3_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \tok.i50_4_lut_adj_151_LC_5_3_0  (
            .in0(N__16940),
            .in1(N__29607),
            .in2(N__16859),
            .in3(N__14735),
            .lcout(\tok.n27_adj_825 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_154_LC_5_3_1 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_154_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_154_LC_5_3_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \tok.i50_4_lut_adj_154_LC_5_3_1  (
            .in0(N__14657),
            .in1(N__16941),
            .in2(N__27353),
            .in3(N__16853),
            .lcout(),
            .ltout(\tok.n27_adj_828_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i5_LC_5_3_2 .C_ON=1'b0;
    defparam \tok.idx_i5_LC_5_3_2 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i5_LC_5_3_2 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \tok.idx_i5_LC_5_3_2  (
            .in0(N__16700),
            .in1(N__14697),
            .in2(N__12287),
            .in3(N__16734),
            .lcout(\tok.idx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28481),
            .ce(),
            .sr(N__28234));
    defparam \tok.i50_4_lut_adj_157_LC_5_3_3 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_157_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_157_LC_5_3_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \tok.i50_4_lut_adj_157_LC_5_3_3  (
            .in0(N__16942),
            .in1(N__16854),
            .in2(N__21894),
            .in3(N__14582),
            .lcout(),
            .ltout(\tok.n27_adj_831_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i6_LC_5_3_4 .C_ON=1'b0;
    defparam \tok.idx_i6_LC_5_3_4 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i6_LC_5_3_4 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \tok.idx_i6_LC_5_3_4  (
            .in0(N__16701),
            .in1(N__14622),
            .in2(N__12284),
            .in3(N__16735),
            .lcout(\tok.idx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28481),
            .ce(),
            .sr(N__28234));
    defparam \tok.i50_4_lut_adj_160_LC_5_3_5 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_160_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_160_LC_5_3_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \tok.i50_4_lut_adj_160_LC_5_3_5  (
            .in0(N__16943),
            .in1(N__16855),
            .in2(N__22321),
            .in3(N__14513),
            .lcout(),
            .ltout(\tok.n27_adj_833_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i7_LC_5_3_6 .C_ON=1'b0;
    defparam \tok.idx_i7_LC_5_3_6 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i7_LC_5_3_6 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \tok.idx_i7_LC_5_3_6  (
            .in0(N__16702),
            .in1(N__14545),
            .in2(N__12281),
            .in3(N__16736),
            .lcout(\tok.idx_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28481),
            .ce(),
            .sr(N__28234));
    defparam \tok.idx_i4_LC_5_3_7 .C_ON=1'b0;
    defparam \tok.idx_i4_LC_5_3_7 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i4_LC_5_3_7 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \tok.idx_i4_LC_5_3_7  (
            .in0(N__16733),
            .in1(N__16699),
            .in2(N__14778),
            .in3(N__12479),
            .lcout(\tok.idx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28481),
            .ce(),
            .sr(N__28234));
    defparam \tok.i1_2_lut_3_lut_4_lut_LC_5_4_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_LC_5_4_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_LC_5_4_0  (
            .in0(N__16923),
            .in1(N__12446),
            .in2(N__12421),
            .in3(N__22140),
            .lcout(\tok.n17_adj_777 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_136_LC_5_4_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_136_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_136_LC_5_4_1 .LUT_INIT=16'b0100000000000100;
    LogicCell40 \tok.i1_4_lut_adj_136_LC_5_4_1  (
            .in0(N__18351),
            .in1(N__18052),
            .in2(N__12380),
            .in3(N__20297),
            .lcout(),
            .ltout(\tok.n5285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_137_LC_5_4_2 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_137_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_137_LC_5_4_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \tok.i4_4_lut_adj_137_LC_5_4_2  (
            .in0(N__17416),
            .in1(N__12388),
            .in2(N__12473),
            .in3(N__30025),
            .lcout(\tok.n1_adj_715 ),
            .ltout(\tok.n1_adj_715_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2571_2_lut_LC_5_4_3 .C_ON=1'b0;
    defparam \tok.i2571_2_lut_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2571_2_lut_LC_5_4_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \tok.i2571_2_lut_LC_5_4_3  (
            .in0(N__12378),
            .in1(_gnd_net_),
            .in2(N__12470),
            .in3(_gnd_net_),
            .lcout(\tok.n190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_108_LC_5_4_4 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_108_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_108_LC_5_4_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \tok.i4_4_lut_adj_108_LC_5_4_4  (
            .in0(N__20298),
            .in1(N__18352),
            .in2(N__17420),
            .in3(N__18059),
            .lcout(),
            .ltout(\tok.n10_adj_763_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_4_lut_LC_5_4_5 .C_ON=1'b0;
    defparam \tok.i5_3_lut_4_lut_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_4_lut_LC_5_4_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \tok.i5_3_lut_4_lut_LC_5_4_5  (
            .in0(N__12389),
            .in1(N__12452),
            .in2(N__12425),
            .in3(N__12415),
            .lcout(\tok.n238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5175_2_lut_3_lut_LC_5_4_6 .C_ON=1'b0;
    defparam \tok.i5175_2_lut_3_lut_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5175_2_lut_3_lut_LC_5_4_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i5175_2_lut_3_lut_LC_5_4_6  (
            .in0(N__16922),
            .in1(N__22139),
            .in2(_gnd_net_),
            .in3(N__19246),
            .lcout(\tok.n5340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_162_LC_5_4_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_162_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_162_LC_5_4_7 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_162_LC_5_4_7  (
            .in0(N__12377),
            .in1(N__12357),
            .in2(N__16499),
            .in3(N__16432),
            .lcout(\tok.n4_adj_813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_54_LC_5_5_0 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_54_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_54_LC_5_5_0 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \tok.i27_4_lut_adj_54_LC_5_5_0  (
            .in0(N__20278),
            .in1(N__12503),
            .in2(N__12494),
            .in3(N__19256),
            .lcout(),
            .ltout(\tok.n13_adj_691_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_55_LC_5_5_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_55_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_55_LC_5_5_1 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \tok.i1_4_lut_adj_55_LC_5_5_1  (
            .in0(N__16353),
            .in1(N__16294),
            .in2(N__12530),
            .in3(N__15313),
            .lcout(n10_adj_871),
            .ltout(n10_adj_871_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_82_LC_5_5_2 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_82_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_82_LC_5_5_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \tok.i26_3_lut_adj_82_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__16134),
            .in2(N__12527),
            .in3(N__14105),
            .lcout(\tok.tc_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5541_4_lut_LC_5_5_3 .C_ON=1'b0;
    defparam \tok.ram.i5541_4_lut_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5541_4_lut_LC_5_5_3 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \tok.ram.i5541_4_lut_LC_5_5_3  (
            .in0(N__15964),
            .in1(N__19897),
            .in2(N__14084),
            .in3(N__15312),
            .lcout(),
            .ltout(\tok.ram.n5605_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6_4_lut_adj_24_LC_5_5_4 .C_ON=1'b0;
    defparam \tok.ram.i6_4_lut_adj_24_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6_4_lut_adj_24_LC_5_5_4 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.ram.i6_4_lut_adj_24_LC_5_5_4  (
            .in0(N__14083),
            .in1(N__15874),
            .in2(N__12506),
            .in3(N__30031),
            .lcout(\tok.n3_adj_690 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_51_LC_5_5_5 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_51_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_51_LC_5_5_5 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_51_LC_5_5_5  (
            .in0(N__14079),
            .in1(N__18350),
            .in2(N__17279),
            .in3(N__20277),
            .lcout(),
            .ltout(\tok.n83_adj_687_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5480_2_lut_3_lut_LC_5_5_6 .C_ON=1'b0;
    defparam \tok.i5480_2_lut_3_lut_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5480_2_lut_3_lut_LC_5_5_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i5480_2_lut_3_lut_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(N__19070),
            .in2(N__12497),
            .in3(N__30030),
            .lcout(\tok.n5505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i6_LC_5_5_7 .C_ON=1'b0;
    defparam \tok.tc_i6_LC_5_5_7 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i6_LC_5_5_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.tc_i6_LC_5_5_7  (
            .in0(N__16135),
            .in1(_gnd_net_),
            .in2(N__14113),
            .in3(N__12485),
            .lcout(tc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28492),
            .ce(),
            .sr(N__28213));
    defparam \tok.i125_4_lut_adj_198_LC_5_6_0 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_198_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_198_LC_5_6_0 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \tok.i125_4_lut_adj_198_LC_5_6_0  (
            .in0(N__18361),
            .in1(N__12612),
            .in2(N__17459),
            .in3(N__20311),
            .lcout(),
            .ltout(\tok.n83_adj_848_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5545_2_lut_3_lut_LC_5_6_1 .C_ON=1'b0;
    defparam \tok.i5545_2_lut_3_lut_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5545_2_lut_3_lut_LC_5_6_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i5545_2_lut_3_lut_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(N__19058),
            .in2(N__12620),
            .in3(N__30026),
            .lcout(\tok.n5610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5527_4_lut_LC_5_6_2 .C_ON=1'b0;
    defparam \tok.ram.i5527_4_lut_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5527_4_lut_LC_5_6_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.ram.i5527_4_lut_LC_5_6_2  (
            .in0(N__15960),
            .in1(N__12711),
            .in2(N__12617),
            .in3(N__19901),
            .lcout(),
            .ltout(\tok.ram.n5594_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6_4_lut_LC_5_6_3 .C_ON=1'b0;
    defparam \tok.ram.i6_4_lut_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6_4_lut_LC_5_6_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.ram.i6_4_lut_LC_5_6_3  (
            .in0(N__15860),
            .in1(N__12616),
            .in2(N__12590),
            .in3(N__30027),
            .lcout(),
            .ltout(\tok.n3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_LC_5_6_4 .C_ON=1'b0;
    defparam \tok.i27_4_lut_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_LC_5_6_4 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i27_4_lut_LC_5_6_4  (
            .in0(N__12587),
            .in1(N__19245),
            .in2(N__12581),
            .in3(N__20312),
            .lcout(),
            .ltout(\tok.n13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_LC_5_6_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_LC_5_6_5 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \tok.i1_4_lut_LC_5_6_5  (
            .in0(N__12712),
            .in1(N__16281),
            .in2(N__12578),
            .in3(N__16357),
            .lcout(n10_adj_866),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_4_lut_LC_5_6_6 .C_ON=1'b0;
    defparam \tok.uart.i1_4_lut_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_4_lut_LC_5_6_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \tok.uart.i1_4_lut_LC_5_6_6  (
            .in0(N__15995),
            .in1(N__17048),
            .in2(N__17330),
            .in3(N__12575),
            .lcout(rx_data_7__N_511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_65_LC_5_6_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_65_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_65_LC_5_6_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_65_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__19057),
            .in2(_gnd_net_),
            .in3(N__18360),
            .lcout(\tok.n101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i11_4_lut_adj_103_LC_5_7_0 .C_ON=1'b0;
    defparam \tok.i11_4_lut_adj_103_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i11_4_lut_adj_103_LC_5_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i11_4_lut_adj_103_LC_5_7_0  (
            .in0(N__12872),
            .in1(N__12560),
            .in2(N__12548),
            .in3(N__12887),
            .lcout(\tok.n27_adj_757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_81_LC_5_7_1 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_81_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_81_LC_5_7_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i5_4_lut_adj_81_LC_5_7_1  (
            .in0(N__12559),
            .in1(N__12544),
            .in2(N__21631),
            .in3(N__29266),
            .lcout(),
            .ltout(\tok.n21_adj_733_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i14_4_lut_adj_107_LC_5_7_2 .C_ON=1'b0;
    defparam \tok.i14_4_lut_adj_107_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i14_4_lut_adj_107_LC_5_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i14_4_lut_adj_107_LC_5_7_2  (
            .in0(N__12845),
            .in1(N__12857),
            .in2(N__12533),
            .in3(N__12851),
            .lcout(\tok.n30_adj_761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_71_LC_5_7_3 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_71_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_71_LC_5_7_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i6_4_lut_adj_71_LC_5_7_3  (
            .in0(N__12886),
            .in1(N__12871),
            .in2(N__22320),
            .in3(N__22757),
            .lcout(\tok.n22_adj_721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_79_LC_5_7_4 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_79_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_79_LC_5_7_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i7_4_lut_adj_79_LC_5_7_4  (
            .in0(N__12838),
            .in1(N__12796),
            .in2(N__25765),
            .in3(N__25158),
            .lcout(\tok.n23_adj_731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_4_lut_adj_33_LC_5_7_5 .C_ON=1'b0;
    defparam \tok.i8_4_lut_adj_33_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i8_4_lut_adj_33_LC_5_7_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i8_4_lut_adj_33_LC_5_7_5  (
            .in0(N__12826),
            .in1(N__12808),
            .in2(N__24862),
            .in3(N__29070),
            .lcout(\tok.n24_adj_651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i12_4_lut_adj_101_LC_5_7_6 .C_ON=1'b0;
    defparam \tok.i12_4_lut_adj_101_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i12_4_lut_adj_101_LC_5_7_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i12_4_lut_adj_101_LC_5_7_6  (
            .in0(N__12839),
            .in1(N__12827),
            .in2(N__12812),
            .in3(N__12797),
            .lcout(\tok.n28_adj_755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_LC_5_7_7 .C_ON=1'b0;
    defparam \tok.i5_4_lut_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_LC_5_7_7 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \tok.i5_4_lut_LC_5_7_7  (
            .in0(N__21619),
            .in1(N__24481),
            .in2(N__27460),
            .in3(N__29267),
            .lcout(\tok.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_2_lut_LC_5_8_0 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_2_lut_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_2_lut_LC_5_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_2_lut_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__12784),
            .in2(_gnd_net_),
            .in3(N__12719),
            .lcout(\tok.tc_plus_1_0 ),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\tok.n4754 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_3_lut_LC_5_8_1 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_3_lut_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_3_lut_LC_5_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_3_lut_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__15726),
            .in2(_gnd_net_),
            .in3(N__12686),
            .lcout(\tok.tc_plus_1_1 ),
            .ltout(),
            .carryin(\tok.n4754 ),
            .carryout(\tok.n4755 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_4_lut_LC_5_8_2 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_4_lut_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_4_lut_LC_5_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_4_lut_LC_5_8_2  (
            .in0(_gnd_net_),
            .in1(N__12683),
            .in2(_gnd_net_),
            .in3(N__12623),
            .lcout(\tok.tc_plus_1_2 ),
            .ltout(),
            .carryin(\tok.n4755 ),
            .carryout(\tok.n4756 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_5_lut_LC_5_8_3 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_5_lut_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_5_lut_LC_5_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_5_lut_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13090),
            .in3(N__13055),
            .lcout(\tok.tc_plus_1_3 ),
            .ltout(),
            .carryin(\tok.n4756 ),
            .carryout(\tok.n4757 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_6_lut_LC_5_8_4 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_6_lut_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_6_lut_LC_5_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_6_lut_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(N__16106),
            .in2(_gnd_net_),
            .in3(N__13052),
            .lcout(\tok.tc_plus_1_4 ),
            .ltout(),
            .carryin(\tok.n4757 ),
            .carryout(\tok.n4758 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_7_lut_LC_5_8_5 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_7_lut_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_7_lut_LC_5_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_7_lut_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(N__13040),
            .in2(_gnd_net_),
            .in3(N__12995),
            .lcout(\tok.tc_plus_1_5 ),
            .ltout(),
            .carryin(\tok.n4758 ),
            .carryout(\tok.n4759 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_8_lut_LC_5_8_6 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_8_lut_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_8_lut_LC_5_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_8_lut_LC_5_8_6  (
            .in0(_gnd_net_),
            .in1(N__14112),
            .in2(_gnd_net_),
            .in3(N__12992),
            .lcout(\tok.tc_plus_1_6 ),
            .ltout(),
            .carryin(\tok.n4759 ),
            .carryout(\tok.n4760 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_9_lut_LC_5_8_7 .C_ON=1'b0;
    defparam \tok.tc_7__I_0_9_lut_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_9_lut_LC_5_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_9_lut_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(N__12989),
            .in2(_gnd_net_),
            .in3(N__12962),
            .lcout(\tok.tc_plus_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5608_2_lut_3_lut_LC_5_9_0 .C_ON=1'b0;
    defparam \tok.i5608_2_lut_3_lut_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5608_2_lut_3_lut_LC_5_9_0 .LUT_INIT=16'b0000010000000100;
    LogicCell40 \tok.i5608_2_lut_3_lut_LC_5_9_0  (
            .in0(N__17611),
            .in1(N__18386),
            .in2(N__22510),
            .in3(_gnd_net_),
            .lcout(\tok.write_flag ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5234_4_lut_LC_5_9_1 .C_ON=1'b0;
    defparam \tok.i5234_4_lut_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5234_4_lut_LC_5_9_1 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \tok.i5234_4_lut_LC_5_9_1  (
            .in0(N__18385),
            .in1(N__17610),
            .in2(N__12932),
            .in3(N__15589),
            .lcout(\tok.n5406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_157_i15_2_lut_3_lut_LC_5_9_2 .C_ON=1'b0;
    defparam \tok.equal_157_i15_2_lut_3_lut_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.equal_157_i15_2_lut_3_lut_LC_5_9_2 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \tok.equal_157_i15_2_lut_3_lut_LC_5_9_2  (
            .in0(N__17528),
            .in1(N__15815),
            .in2(_gnd_net_),
            .in3(N__15423),
            .lcout(\tok.n15_adj_671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_LC_5_9_3 .C_ON=1'b0;
    defparam \tok.i5_3_lut_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_LC_5_9_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \tok.i5_3_lut_LC_5_9_3  (
            .in0(N__12893),
            .in1(_gnd_net_),
            .in2(N__23278),
            .in3(N__15590),
            .lcout(),
            .ltout(\tok.n14_adj_688_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2652_4_lut_LC_5_9_4 .C_ON=1'b0;
    defparam \tok.i2652_4_lut_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2652_4_lut_LC_5_9_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \tok.i2652_4_lut_LC_5_9_4  (
            .in0(N__13178),
            .in1(N__15814),
            .in2(N__13166),
            .in3(N__13097),
            .lcout(\tok.n2735 ),
            .ltout(\tok.n2735_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_4_i1_3_lut_LC_5_9_5 .C_ON=1'b0;
    defparam \tok.select_73_Select_4_i1_3_lut_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_4_i1_3_lut_LC_5_9_5 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \tok.select_73_Select_4_i1_3_lut_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(N__27756),
            .in2(N__13163),
            .in3(N__19042),
            .lcout(),
            .ltout(\tok.n1_adj_850_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_186_LC_5_9_6 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_186_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_186_LC_5_9_6 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \tok.i6_4_lut_adj_186_LC_5_9_6  (
            .in0(N__23212),
            .in1(N__13253),
            .in2(N__13160),
            .in3(N__21632),
            .lcout(\tok.n17_adj_853 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_155_i16_2_lut_3_lut_LC_5_9_7 .C_ON=1'b0;
    defparam \tok.equal_155_i16_2_lut_3_lut_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.equal_155_i16_2_lut_3_lut_LC_5_9_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \tok.equal_155_i16_2_lut_3_lut_LC_5_9_7  (
            .in0(N__15424),
            .in1(N__22450),
            .in2(_gnd_net_),
            .in3(N__17529),
            .lcout(\tok.n400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_98_LC_5_10_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_98_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_98_LC_5_10_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \tok.i1_4_lut_adj_98_LC_5_10_0  (
            .in0(N__13157),
            .in1(N__13151),
            .in2(N__16004),
            .in3(N__19681),
            .lcout(\tok.n5254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5210_4_lut_4_lut_LC_5_10_1 .C_ON=1'b0;
    defparam \tok.i5210_4_lut_4_lut_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5210_4_lut_4_lut_LC_5_10_1 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \tok.i5210_4_lut_4_lut_LC_5_10_1  (
            .in0(N__15419),
            .in1(N__23258),
            .in2(N__17531),
            .in3(N__15451),
            .lcout(\tok.n5380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_129_LC_5_10_2 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_129_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_129_LC_5_10_2 .LUT_INIT=16'b1111000111111111;
    LogicCell40 \tok.i4_4_lut_adj_129_LC_5_10_2  (
            .in0(N__17598),
            .in1(N__15417),
            .in2(N__13145),
            .in3(N__13128),
            .lcout(),
            .ltout(\tok.n5271_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_130_LC_5_10_3 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_130_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_130_LC_5_10_3 .LUT_INIT=16'b1111000111111111;
    LogicCell40 \tok.i2_4_lut_adj_130_LC_5_10_3  (
            .in0(N__15418),
            .in1(N__15450),
            .in2(N__13112),
            .in3(N__23377),
            .lcout(\tok.n5272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_56_LC_5_10_4 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_56_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_56_LC_5_10_4 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \tok.i6_4_lut_adj_56_LC_5_10_4  (
            .in0(N__13109),
            .in1(N__13103),
            .in2(N__17612),
            .in3(N__19680),
            .lcout(\tok.n15_adj_695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i4_LC_5_10_5 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i4_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i4_LC_5_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.rx_data_i0_i4_LC_5_10_5  (
            .in0(N__13262),
            .in1(N__23039),
            .in2(_gnd_net_),
            .in3(N__25679),
            .lcout(uart_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28523),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_4_i12_2_lut_3_lut_LC_5_10_6 .C_ON=1'b0;
    defparam \tok.select_73_Select_4_i12_2_lut_3_lut_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_4_i12_2_lut_3_lut_LC_5_10_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \tok.select_73_Select_4_i12_2_lut_3_lut_LC_5_10_6  (
            .in0(N__23259),
            .in1(N__13261),
            .in2(_gnd_net_),
            .in3(N__22411),
            .lcout(\tok.n12_adj_826 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_213_i15_2_lut_LC_5_10_7 .C_ON=1'b0;
    defparam \tok.T_7__I_0_213_i15_2_lut_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_213_i15_2_lut_LC_5_10_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.T_7__I_0_213_i15_2_lut_LC_5_10_7  (
            .in0(N__13237),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17487),
            .lcout(\tok.n15_adj_789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i3_LC_5_11_0 .C_ON=1'b0;
    defparam \tok.uart.sender_i3_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i3_LC_5_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i3_LC_5_11_0  (
            .in0(N__13208),
            .in1(N__14366),
            .in2(_gnd_net_),
            .in3(N__27755),
            .lcout(sender_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28527),
            .ce(N__14300),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i4_LC_5_11_1 .C_ON=1'b0;
    defparam \tok.uart.sender_i4_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i4_LC_5_11_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.sender_i4_LC_5_11_1  (
            .in0(N__14367),
            .in1(N__13202),
            .in2(_gnd_net_),
            .in3(N__21131),
            .lcout(\tok.uart.sender_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28527),
            .ce(N__14300),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i5_LC_5_11_2 .C_ON=1'b0;
    defparam \tok.uart.sender_i5_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i5_LC_5_11_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i5_LC_5_11_2  (
            .in0(N__13196),
            .in1(N__14368),
            .in2(_gnd_net_),
            .in3(N__22758),
            .lcout(\tok.uart.sender_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28527),
            .ce(N__14300),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i6_LC_5_11_3 .C_ON=1'b0;
    defparam \tok.uart.sender_i6_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i6_LC_5_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.sender_i6_LC_5_11_3  (
            .in0(N__14369),
            .in1(N__13190),
            .in2(_gnd_net_),
            .in3(N__29731),
            .lcout(\tok.uart.sender_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28527),
            .ce(N__14300),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i7_LC_5_11_4 .C_ON=1'b0;
    defparam \tok.uart.sender_i7_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i7_LC_5_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i7_LC_5_11_4  (
            .in0(N__13184),
            .in1(N__14370),
            .in2(_gnd_net_),
            .in3(N__29596),
            .lcout(\tok.uart.sender_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28527),
            .ce(N__14300),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i8_LC_5_11_5 .C_ON=1'b0;
    defparam \tok.uart.sender_i8_LC_5_11_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i8_LC_5_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.sender_i8_LC_5_11_5  (
            .in0(N__14371),
            .in1(N__14306),
            .in2(_gnd_net_),
            .in3(N__27347),
            .lcout(\tok.uart.sender_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28527),
            .ce(N__14300),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i9_LC_5_11_6 .C_ON=1'b0;
    defparam \tok.uart.sender_i9_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i9_LC_5_11_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i9_LC_5_11_6  (
            .in0(N__14408),
            .in1(N__14372),
            .in2(_gnd_net_),
            .in3(N__21893),
            .lcout(\tok.uart.sender_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28527),
            .ce(N__14300),
            .sr(_gnd_net_));
    defparam \tok.equal_114_i10_2_lut_LC_5_11_7 .C_ON=1'b0;
    defparam \tok.equal_114_i10_2_lut_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.equal_114_i10_2_lut_LC_5_11_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.equal_114_i10_2_lut_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__18002),
            .in2(_gnd_net_),
            .in3(N__29958),
            .lcout(\tok.n10_adj_643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i6_LC_5_12_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i6_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i6_LC_5_12_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.C_stk.tail_i0_i6_LC_5_12_0  (
            .in0(N__14024),
            .in1(N__14070),
            .in2(N__13721),
            .in3(N__13748),
            .lcout(\tok.C_stk.tail_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28530),
            .ce(N__13362),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i5265_3_lut_LC_5_12_1 .C_ON=1'b0;
    defparam \tok.C_stk.i5265_3_lut_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i5265_3_lut_LC_5_12_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i5265_3_lut_LC_5_12_1  (
            .in0(N__14053),
            .in1(N__14270),
            .in2(_gnd_net_),
            .in3(N__15314),
            .lcout(),
            .ltout(\tok.C_stk.n5438_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i6_LC_5_12_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i6_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i6_LC_5_12_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i6_LC_5_12_2  (
            .in0(N__14185),
            .in1(N__15517),
            .in2(N__14117),
            .in3(N__14114),
            .lcout(\tok.c_stk_r_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28530),
            .ce(N__13362),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i14_LC_5_12_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i14_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i14_LC_5_12_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.C_stk.tail_i0_i14_LC_5_12_3  (
            .in0(N__14054),
            .in1(N__13716),
            .in2(N__13396),
            .in3(N__14025),
            .lcout(\tok.tail_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28530),
            .ce(N__13362),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i22_LC_5_12_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i22_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i22_LC_5_12_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.C_stk.tail_i0_i22_LC_5_12_4  (
            .in0(N__14023),
            .in1(N__13747),
            .in2(N__13739),
            .in3(N__13720),
            .lcout(\tok.C_stk.tail_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28530),
            .ce(N__13362),
            .sr(_gnd_net_));
    defparam \tok.tc_i1_LC_5_13_0 .C_ON=1'b0;
    defparam \tok.tc_i1_LC_5_13_0 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i1_LC_5_13_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.tc_i1_LC_5_13_0  (
            .in0(N__15752),
            .in1(N__16204),
            .in2(_gnd_net_),
            .in3(N__15722),
            .lcout(tc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28535),
            .ce(),
            .sr(N__28128));
    defparam \tok.inv_106_i14_1_lut_LC_5_13_1 .C_ON=1'b0;
    defparam \tok.inv_106_i14_1_lut_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i14_1_lut_LC_5_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i14_1_lut_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23154),
            .lcout(\tok.n289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.reset_I_0_1_lut_LC_5_13_2 .C_ON=1'b0;
    defparam \tok.reset_I_0_1_lut_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.reset_I_0_1_lut_LC_5_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.reset_I_0_1_lut_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14507),
            .lcout(\tok.reset_N_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i16_LC_6_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i16_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i16_LC_6_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i16_LC_6_2_0  (
            .in0(N__14486),
            .in1(N__14417),
            .in2(_gnd_net_),
            .in3(N__26402),
            .lcout(\tok.A_stk.tail_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28482),
            .ce(N__26019),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i0_LC_6_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i0_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i0_LC_6_2_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i0_LC_6_2_1  (
            .in0(N__26401),
            .in1(_gnd_net_),
            .in2(N__14498),
            .in3(N__22840),
            .lcout(\tok.A_stk.tail_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28482),
            .ce(N__26019),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i32_LC_6_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i32_LC_6_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i32_LC_6_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i32_LC_6_2_2  (
            .in0(N__14477),
            .in1(N__14494),
            .in2(_gnd_net_),
            .in3(N__26403),
            .lcout(\tok.A_stk.tail_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28482),
            .ce(N__26019),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i48_LC_6_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i48_LC_6_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i48_LC_6_2_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i48_LC_6_2_3  (
            .in0(N__26404),
            .in1(N__14485),
            .in2(_gnd_net_),
            .in3(N__14468),
            .lcout(\tok.A_stk.tail_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28482),
            .ce(N__26019),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i64_LC_6_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i64_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i64_LC_6_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i64_LC_6_2_4  (
            .in0(N__14476),
            .in1(N__14441),
            .in2(_gnd_net_),
            .in3(N__26405),
            .lcout(\tok.A_stk.tail_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28482),
            .ce(N__26019),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i80_LC_6_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i80_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i80_LC_6_2_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i80_LC_6_2_5  (
            .in0(N__26406),
            .in1(_gnd_net_),
            .in2(N__14432),
            .in3(N__14467),
            .lcout(\tok.A_stk.tail_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28482),
            .ce(N__26019),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i96_LC_6_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i96_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i96_LC_6_2_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i96_LC_6_2_6  (
            .in0(N__14458),
            .in1(N__14440),
            .in2(_gnd_net_),
            .in3(N__26407),
            .lcout(tail_96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28482),
            .ce(N__26019),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i0_LC_6_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i0_LC_6_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i0_LC_6_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i0_LC_6_2_7  (
            .in0(N__14416),
            .in1(N__25466),
            .in2(_gnd_net_),
            .in3(N__27783),
            .lcout(\tok.S_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28482),
            .ce(N__26019),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_2_lut_LC_6_3_0 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_2_lut_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_2_lut_LC_6_3_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_2_lut_LC_6_3_0  (
            .in0(N__14849),
            .in1(N__14848),
            .in2(N__15229),
            .in3(N__14813),
            .lcout(\tok.n33 ),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\tok.n4747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_3_lut_LC_6_3_1 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_3_lut_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_3_lut_LC_6_3_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_3_lut_LC_6_3_1  (
            .in0(N__16631),
            .in1(N__16630),
            .in2(N__15233),
            .in3(N__14810),
            .lcout(\tok.n33_adj_814 ),
            .ltout(),
            .carryin(\tok.n4747 ),
            .carryout(\tok.n4748 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_4_lut_LC_6_3_2 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_4_lut_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_4_lut_LC_6_3_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_4_lut_LC_6_3_2  (
            .in0(N__16974),
            .in1(N__16973),
            .in2(N__15230),
            .in3(N__14807),
            .lcout(\tok.n33_adj_816 ),
            .ltout(),
            .carryin(\tok.n4748 ),
            .carryout(\tok.n4749 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_5_lut_LC_6_3_3 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_5_lut_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_5_lut_LC_6_3_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_5_lut_LC_6_3_3  (
            .in0(N__16769),
            .in1(N__16768),
            .in2(N__15234),
            .in3(N__14804),
            .lcout(\tok.n33_adj_821 ),
            .ltout(),
            .carryin(\tok.n4749 ),
            .carryout(\tok.n4750 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_6_lut_LC_6_3_4 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_6_lut_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_6_lut_LC_6_3_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_6_lut_LC_6_3_4  (
            .in0(N__14768),
            .in1(N__14767),
            .in2(N__15231),
            .in3(N__14729),
            .lcout(\tok.n33_adj_819 ),
            .ltout(),
            .carryin(\tok.n4750 ),
            .carryout(\tok.n4751 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_7_lut_LC_6_3_5 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_7_lut_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_7_lut_LC_6_3_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_7_lut_LC_6_3_5  (
            .in0(N__14696),
            .in1(N__14695),
            .in2(N__15235),
            .in3(N__14651),
            .lcout(\tok.n33_adj_811 ),
            .ltout(),
            .carryin(\tok.n4751 ),
            .carryout(\tok.n4752 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_8_lut_LC_6_3_6 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_8_lut_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_8_lut_LC_6_3_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_8_lut_LC_6_3_6  (
            .in0(N__14615),
            .in1(N__14614),
            .in2(N__15232),
            .in3(N__14576),
            .lcout(\tok.n33_adj_804 ),
            .ltout(),
            .carryin(\tok.n4752 ),
            .carryout(\tok.n4753 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_9_lut_LC_6_3_7 .C_ON=1'b0;
    defparam \tok.idx_7__I_0_9_lut_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_9_lut_LC_6_3_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_9_lut_LC_6_3_7  (
            .in0(N__14552),
            .in1(N__14553),
            .in2(N__15236),
            .in3(N__14516),
            .lcout(\tok.n33_adj_801 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_LC_6_4_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_LC_6_4_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.i1_2_lut_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(N__16837),
            .in2(_gnd_net_),
            .in3(N__15186),
            .lcout(\tok.n5 ),
            .ltout(\tok.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_72_LC_6_4_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_72_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_72_LC_6_4_1 .LUT_INIT=16'b1011101010111011;
    LogicCell40 \tok.i1_4_lut_adj_72_LC_6_4_1  (
            .in0(N__17768),
            .in1(N__15560),
            .in2(N__14897),
            .in3(N__16930),
            .lcout(stall_),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.stall_200_LC_6_4_2 .C_ON=1'b0;
    defparam \tok.stall_200_LC_6_4_2 .SEQ_MODE=4'b1010;
    defparam \tok.stall_200_LC_6_4_2 .LUT_INIT=16'b1100111111001101;
    LogicCell40 \tok.stall_200_LC_6_4_2  (
            .in0(N__16933),
            .in1(N__17771),
            .in2(N__15566),
            .in3(N__14894),
            .lcout(\tok.stall ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28493),
            .ce(),
            .sr(N__28237));
    defparam \tok.i1_4_lut_adj_132_LC_6_4_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_132_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_132_LC_6_4_3 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \tok.i1_4_lut_adj_132_LC_6_4_3  (
            .in0(N__17770),
            .in1(N__15562),
            .in2(N__16857),
            .in3(N__16931),
            .lcout(\tok.n5282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.search_clk_198_LC_6_4_4 .C_ON=1'b0;
    defparam \tok.search_clk_198_LC_6_4_4 .SEQ_MODE=4'b1010;
    defparam \tok.search_clk_198_LC_6_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.search_clk_198_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16844),
            .lcout(\tok.search_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28493),
            .ce(),
            .sr(N__28237));
    defparam \tok.i50_4_lut_LC_6_4_5 .C_ON=1'b0;
    defparam \tok.i50_4_lut_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_LC_6_4_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \tok.i50_4_lut_LC_6_4_5  (
            .in0(N__27770),
            .in1(N__14888),
            .in2(N__16856),
            .in3(N__16932),
            .lcout(),
            .ltout(\tok.n27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i0_LC_6_4_6 .C_ON=1'b0;
    defparam \tok.idx_i0_LC_6_4_6 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i0_LC_6_4_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \tok.idx_i0_LC_6_4_6  (
            .in0(N__14850),
            .in1(N__16693),
            .in2(N__14882),
            .in3(N__16729),
            .lcout(\tok.idx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28493),
            .ce(),
            .sr(N__28237));
    defparam \tok.i2622_2_lut_LC_6_4_7 .C_ON=1'b0;
    defparam \tok.i2622_2_lut_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2622_2_lut_LC_6_4_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i2622_2_lut_LC_6_4_7  (
            .in0(N__17769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15561),
            .lcout(\tok.n2699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_34_LC_6_5_0 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_34_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_34_LC_6_5_0 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \tok.i125_4_lut_adj_34_LC_6_5_0  (
            .in0(N__18367),
            .in1(N__15018),
            .in2(N__15395),
            .in3(N__20313),
            .lcout(),
            .ltout(\tok.n83_adj_652_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5442_2_lut_3_lut_LC_6_5_1 .C_ON=1'b0;
    defparam \tok.i5442_2_lut_3_lut_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5442_2_lut_3_lut_LC_6_5_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i5442_2_lut_3_lut_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__19071),
            .in2(N__14816),
            .in3(N__30028),
            .lcout(\tok.n5460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5518_4_lut_LC_6_5_2 .C_ON=1'b0;
    defparam \tok.ram.i5518_4_lut_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5518_4_lut_LC_6_5_2 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \tok.ram.i5518_4_lut_LC_6_5_2  (
            .in0(N__15965),
            .in1(N__14976),
            .in2(N__19904),
            .in3(N__15019),
            .lcout(),
            .ltout(\tok.ram.n5580_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6_4_lut_adj_21_LC_6_5_3 .C_ON=1'b0;
    defparam \tok.ram.i6_4_lut_adj_21_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6_4_lut_adj_21_LC_6_5_3 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.ram.i6_4_lut_adj_21_LC_6_5_3  (
            .in0(N__15020),
            .in1(N__15873),
            .in2(N__14993),
            .in3(N__30029),
            .lcout(),
            .ltout(\tok.n3_adj_659_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_37_LC_6_5_4 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_37_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_37_LC_6_5_4 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i27_4_lut_adj_37_LC_6_5_4  (
            .in0(N__14990),
            .in1(N__19258),
            .in2(N__14984),
            .in3(N__20315),
            .lcout(),
            .ltout(\tok.n13_adj_660_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_39_LC_6_5_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_39_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_39_LC_6_5_5 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \tok.i1_4_lut_adj_39_LC_6_5_5  (
            .in0(N__14977),
            .in1(N__16370),
            .in2(N__14948),
            .in3(N__16309),
            .lcout(n92_adj_867),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_LC_6_5_6 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_LC_6_5_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.i1_3_lut_4_lut_LC_6_5_6  (
            .in0(N__18368),
            .in1(N__19257),
            .in2(N__18836),
            .in3(N__20314),
            .lcout(),
            .ltout(\tok.n4_adj_778_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_115_LC_6_5_7 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_115_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_115_LC_6_5_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i2_4_lut_adj_115_LC_6_5_7  (
            .in0(N__18046),
            .in1(N__14923),
            .in2(N__14912),
            .in3(N__19072),
            .lcout(\tok.n797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_106_LC_6_6_0 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_106_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_106_LC_6_6_0 .LUT_INIT=16'b1111110111111110;
    LogicCell40 \tok.i10_4_lut_adj_106_LC_6_6_0  (
            .in0(N__29468),
            .in1(N__17018),
            .in2(N__15113),
            .in3(N__15274),
            .lcout(),
            .ltout(\tok.n26_adj_760_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5526_4_lut_LC_6_6_1 .C_ON=1'b0;
    defparam \tok.i5526_4_lut_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5526_4_lut_LC_6_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i5526_4_lut_LC_6_6_1  (
            .in0(N__15026),
            .in1(N__15104),
            .in2(N__14909),
            .in3(N__14906),
            .lcout(),
            .ltout(\tok.n5587_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_138_LC_6_6_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_138_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_138_LC_6_6_2 .LUT_INIT=16'b0000110001000100;
    LogicCell40 \tok.i1_4_lut_adj_138_LC_6_6_2  (
            .in0(N__15640),
            .in1(N__16949),
            .in2(N__14900),
            .in3(N__15242),
            .lcout(\tok.found_slot ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_102_LC_6_6_3 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_102_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_102_LC_6_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i10_4_lut_adj_102_LC_6_6_3  (
            .in0(N__15128),
            .in1(N__17036),
            .in2(N__15275),
            .in3(N__15143),
            .lcout(),
            .ltout(\tok.n26_adj_756_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i15_4_lut_adj_126_LC_6_6_4 .C_ON=1'b0;
    defparam \tok.i15_4_lut_adj_126_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i15_4_lut_adj_126_LC_6_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i15_4_lut_adj_126_LC_6_6_4  (
            .in0(N__15257),
            .in1(N__15062),
            .in2(N__15251),
            .in3(N__15248),
            .lcout(\tok.found_slot_N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_adj_145_LC_6_6_5 .C_ON=1'b0;
    defparam \tok.i2_2_lut_adj_145_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_adj_145_LC_6_6_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i2_2_lut_adj_145_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__15641),
            .in2(_gnd_net_),
            .in3(N__15185),
            .lcout(\tok.write_slot ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_LC_6_6_6 .C_ON=1'b0;
    defparam \tok.i4_4_lut_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_LC_6_6_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i4_4_lut_LC_6_6_6  (
            .in0(N__15142),
            .in1(N__15127),
            .in2(N__27351),
            .in3(N__29724),
            .lcout(\tok.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_105_LC_6_7_0 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_105_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_105_LC_6_7_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i2_4_lut_adj_105_LC_6_7_0  (
            .in0(N__21109),
            .in1(N__15076),
            .in2(N__15098),
            .in3(N__29597),
            .lcout(\tok.n18_adj_759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_104_LC_6_7_1 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_104_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_104_LC_6_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_104_LC_6_7_1  (
            .in0(N__15040),
            .in1(N__15094),
            .in2(N__15080),
            .in3(N__15055),
            .lcout(\tok.n25_adj_758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5505_4_lut_LC_6_7_2 .C_ON=1'b0;
    defparam \tok.i5505_4_lut_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5505_4_lut_LC_6_7_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i5505_4_lut_LC_6_7_2  (
            .in0(N__15056),
            .in1(N__21886),
            .in2(N__27782),
            .in3(N__15041),
            .lcout(\tok.n5590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_175_LC_6_7_3 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_175_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_175_LC_6_7_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i2_3_lut_adj_175_LC_6_7_3  (
            .in0(N__25159),
            .in1(N__20657),
            .in2(_gnd_net_),
            .in3(N__23402),
            .lcout(\tok.n6_adj_843 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i6_LC_6_7_4 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i6_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i6_LC_6_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i6_LC_6_7_4  (
            .in0(N__22916),
            .in1(N__25660),
            .in2(_gnd_net_),
            .in3(N__15356),
            .lcout(uart_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28510),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_6_i12_2_lut_3_lut_LC_6_7_7 .C_ON=1'b0;
    defparam \tok.select_73_Select_6_i12_2_lut_3_lut_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_6_i12_2_lut_3_lut_LC_6_7_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \tok.select_73_Select_6_i12_2_lut_3_lut_LC_6_7_7  (
            .in0(N__15355),
            .in1(N__22511),
            .in2(_gnd_net_),
            .in3(N__23314),
            .lcout(\tok.n12_adj_824 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_176_LC_6_8_0 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_176_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_176_LC_6_8_0 .LUT_INIT=16'b1110111111101110;
    LogicCell40 \tok.i3_4_lut_adj_176_LC_6_8_0  (
            .in0(N__15347),
            .in1(N__23813),
            .in2(N__23335),
            .in3(N__15337),
            .lcout(),
            .ltout(\tok.n31_adj_844_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_177_LC_6_8_1 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_177_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_177_LC_6_8_1 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i3_4_lut_adj_177_LC_6_8_1  (
            .in0(N__22539),
            .in1(N__18047),
            .in2(N__15341),
            .in3(N__19511),
            .lcout(\tok.n10_adj_845 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i3_LC_6_8_3 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i3_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i3_LC_6_8_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.uart.rx_data_i0_i3_LC_6_8_3  (
            .in0(N__15338),
            .in1(_gnd_net_),
            .in2(N__15329),
            .in3(N__25680),
            .lcout(uart_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28517),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_4_lut_adj_188_LC_6_8_4 .C_ON=1'b0;
    defparam \tok.i3_4_lut_4_lut_adj_188_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_4_lut_adj_188_LC_6_8_4 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \tok.i3_4_lut_4_lut_adj_188_LC_6_8_4  (
            .in0(N__28730),
            .in1(N__23665),
            .in2(N__18509),
            .in3(N__29167),
            .lcout(\tok.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i2_LC_6_8_5 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i2_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i2_LC_6_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.uart.capture_i0_i2_LC_6_8_5  (
            .in0(N__21183),
            .in1(N__17344),
            .in2(_gnd_net_),
            .in3(N__22975),
            .lcout(capture_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28517),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i4_LC_6_8_6 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i4_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i4_LC_6_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.capture_i0_i4_LC_6_8_6  (
            .in0(N__22977),
            .in1(N__23035),
            .in2(_gnd_net_),
            .in3(N__15324),
            .lcout(capture_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28517),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i3_LC_6_8_7 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i3_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i3_LC_6_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i3_LC_6_8_7  (
            .in0(N__15325),
            .in1(N__17343),
            .in2(_gnd_net_),
            .in3(N__22976),
            .lcout(capture_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28517),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1774_3_lut_4_lut_LC_6_9_0 .C_ON=1'b0;
    defparam \tok.i1774_3_lut_4_lut_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1774_3_lut_4_lut_LC_6_9_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \tok.i1774_3_lut_4_lut_LC_6_9_0  (
            .in0(N__23667),
            .in1(N__15311),
            .in2(N__22547),
            .in3(N__15629),
            .lcout(\tok.table_wr_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_219_i10_2_lut_LC_6_9_1 .C_ON=1'b0;
    defparam \tok.T_7__I_0_219_i10_2_lut_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_219_i10_2_lut_LC_6_9_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \tok.T_7__I_0_219_i10_2_lut_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__18034),
            .in2(_gnd_net_),
            .in3(N__30013),
            .lcout(\tok.n10_adj_747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2573_3_lut_4_lut_LC_6_9_2 .C_ON=1'b0;
    defparam \tok.i2573_3_lut_4_lut_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2573_3_lut_4_lut_LC_6_9_2 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \tok.i2573_3_lut_4_lut_LC_6_9_2  (
            .in0(N__15432),
            .in1(N__15627),
            .in2(N__22545),
            .in3(N__17613),
            .lcout(\tok.n2635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2620_3_lut_4_lut_LC_6_9_3 .C_ON=1'b0;
    defparam \tok.i2620_3_lut_4_lut_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2620_3_lut_4_lut_LC_6_9_3 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \tok.i2620_3_lut_4_lut_LC_6_9_3  (
            .in0(N__15628),
            .in1(N__15464),
            .in2(N__26979),
            .in3(N__22523),
            .lcout(\tok.n2697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2460_3_lut_4_lut_LC_6_9_4 .C_ON=1'b0;
    defparam \tok.i2460_3_lut_4_lut_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2460_3_lut_4_lut_LC_6_9_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \tok.i2460_3_lut_4_lut_LC_6_9_4  (
            .in0(N__15433),
            .in1(N__15508),
            .in2(N__22546),
            .in3(N__17614),
            .lcout(\tok.n2520 ),
            .ltout(\tok.n2520_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2587_4_lut_LC_6_9_5 .C_ON=1'b0;
    defparam \tok.i2587_4_lut_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2587_4_lut_LC_6_9_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \tok.i2587_4_lut_LC_6_9_5  (
            .in0(N__22527),
            .in1(N__15458),
            .in2(N__15437),
            .in3(N__15434),
            .lcout(\tok.n2661 ),
            .ltout(\tok.n2661_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_179_LC_6_9_6 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_179_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_179_LC_6_9_6 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \tok.i2_4_lut_adj_179_LC_6_9_6  (
            .in0(N__15391),
            .in1(N__25369),
            .in2(N__15368),
            .in3(N__26958),
            .lcout(),
            .ltout(\tok.n9_adj_847_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5562_4_lut_LC_6_9_7 .C_ON=1'b0;
    defparam \tok.i5562_4_lut_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i5562_4_lut_LC_6_9_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i5562_4_lut_LC_6_9_7  (
            .in0(N__15365),
            .in1(N__18398),
            .in2(N__15359),
            .in3(N__19754),
            .lcout(\tok.n5566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_LC_6_10_0 .C_ON=1'b0;
    defparam \tok.i2_3_lut_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_LC_6_10_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \tok.i2_3_lut_LC_6_10_0  (
            .in0(N__15971),
            .in1(N__18420),
            .in2(_gnd_net_),
            .in3(N__18983),
            .lcout(\tok.n880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_116_i14_2_lut_3_lut_4_lut_LC_6_10_1 .C_ON=1'b0;
    defparam \tok.equal_116_i14_2_lut_3_lut_4_lut_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.equal_116_i14_2_lut_3_lut_4_lut_LC_6_10_1 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \tok.equal_116_i14_2_lut_3_lut_4_lut_LC_6_10_1  (
            .in0(N__22109),
            .in1(N__18791),
            .in2(N__19043),
            .in3(N__19217),
            .lcout(\tok.n14_adj_701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_6_10_2 .C_ON=1'b0;
    defparam \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_6_10_2 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_6_10_2  (
            .in0(N__19216),
            .in1(N__18979),
            .in2(N__18815),
            .in3(N__22108),
            .lcout(\tok.n14_adj_807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5260_4_lut_LC_6_10_3 .C_ON=1'b0;
    defparam \tok.i5260_4_lut_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5260_4_lut_LC_6_10_3 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \tok.i5260_4_lut_LC_6_10_3  (
            .in0(N__15806),
            .in1(N__17483),
            .in2(N__16013),
            .in3(N__15794),
            .lcout(),
            .ltout(\tok.n5433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_133_LC_6_10_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_133_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_133_LC_6_10_4 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \tok.i1_4_lut_adj_133_LC_6_10_4  (
            .in0(N__15767),
            .in1(N__15758),
            .in2(N__15788),
            .in3(N__15785),
            .lcout(\tok.n2743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_131_LC_6_10_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_131_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_131_LC_6_10_5 .LUT_INIT=16'b1110111011100000;
    LogicCell40 \tok.i1_4_lut_adj_131_LC_6_10_5  (
            .in0(N__15680),
            .in1(N__17482),
            .in2(N__15779),
            .in3(N__15766),
            .lcout(\tok.n5175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_88_LC_6_10_6 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_88_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_88_LC_6_10_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.i26_3_lut_adj_88_LC_6_10_6  (
            .in0(N__15748),
            .in1(N__16162),
            .in2(_gnd_net_),
            .in3(N__15727),
            .lcout(\tok.tc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i8_LC_6_10_7 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i8_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i8_LC_6_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.uart.capture_i0_i8_LC_6_10_7  (
            .in0(N__22993),
            .in1(N__15991),
            .in2(_gnd_net_),
            .in3(N__22978),
            .lcout(capture_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28528),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_213_i14_2_lut_3_lut_4_lut_LC_6_11_0 .C_ON=1'b0;
    defparam \tok.T_7__I_0_213_i14_2_lut_3_lut_4_lut_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_213_i14_2_lut_3_lut_4_lut_LC_6_11_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \tok.T_7__I_0_213_i14_2_lut_3_lut_4_lut_LC_6_11_0  (
            .in0(N__18777),
            .in1(N__19167),
            .in2(N__22107),
            .in3(N__19044),
            .lcout(\tok.n14_adj_765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_174_LC_6_11_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_174_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_174_LC_6_11_1 .LUT_INIT=16'b1111111111101011;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_174_LC_6_11_1  (
            .in0(N__18016),
            .in1(N__20240),
            .in2(N__30014),
            .in3(N__18354),
            .lcout(\tok.n2_adj_808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5250_3_lut_4_lut_LC_6_11_2 .C_ON=1'b0;
    defparam \tok.i5250_3_lut_4_lut_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5250_3_lut_4_lut_LC_6_11_2 .LUT_INIT=16'b1111111100111111;
    LogicCell40 \tok.i5250_3_lut_4_lut_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__29962),
            .in2(N__20279),
            .in3(N__18017),
            .lcout(\tok.n5423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_143_LC_6_11_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_143_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_143_LC_6_11_3 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_143_LC_6_11_3  (
            .in0(N__18019),
            .in1(N__20245),
            .in2(N__30016),
            .in3(N__18356),
            .lcout(\tok.n42_adj_751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i9_LC_6_11_4 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i9_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i9_LC_6_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i9_LC_6_11_4  (
            .in0(N__17151),
            .in1(N__15990),
            .in2(_gnd_net_),
            .in3(N__22982),
            .lcout(capture_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28531),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_173_LC_6_11_5 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_173_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_173_LC_6_11_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_173_LC_6_11_5  (
            .in0(N__19168),
            .in1(N__22077),
            .in2(_gnd_net_),
            .in3(N__18778),
            .lcout(\tok.n878 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5588_4_lut_4_lut_LC_6_11_6 .C_ON=1'b0;
    defparam \tok.i5588_4_lut_4_lut_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5588_4_lut_4_lut_LC_6_11_6 .LUT_INIT=16'b0011000101110101;
    LogicCell40 \tok.i5588_4_lut_4_lut_LC_6_11_6  (
            .in0(N__18357),
            .in1(N__29969),
            .in2(N__20280),
            .in3(N__18020),
            .lcout(\tok.n5470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2549_2_lut_4_lut_LC_6_11_7 .C_ON=1'b0;
    defparam \tok.i2549_2_lut_4_lut_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2549_2_lut_4_lut_LC_6_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \tok.i2549_2_lut_4_lut_LC_6_11_7  (
            .in0(N__18018),
            .in1(N__20244),
            .in2(N__30015),
            .in3(N__18355),
            .lcout(\tok.n2609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5514_4_lut_LC_6_12_1 .C_ON=1'b0;
    defparam \tok.ram.i5514_4_lut_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5514_4_lut_LC_6_12_1 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.ram.i5514_4_lut_LC_6_12_1  (
            .in0(N__15946),
            .in1(N__16251),
            .in2(N__16072),
            .in3(N__19888),
            .lcout(),
            .ltout(\tok.ram.n5577_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6_4_lut_adj_22_LC_6_12_2 .C_ON=1'b0;
    defparam \tok.ram.i6_4_lut_adj_22_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6_4_lut_adj_22_LC_6_12_2 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \tok.ram.i6_4_lut_adj_22_LC_6_12_2  (
            .in0(N__30020),
            .in1(N__16067),
            .in2(N__15893),
            .in3(N__15882),
            .lcout(\tok.n3_adj_672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_42_LC_6_12_4 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_42_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_42_LC_6_12_4 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \tok.i27_4_lut_adj_42_LC_6_12_4  (
            .in0(N__15821),
            .in1(N__19215),
            .in2(N__16034),
            .in3(N__20276),
            .lcout(),
            .ltout(\tok.n13_adj_673_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_44_LC_6_12_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_44_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_44_LC_6_12_5 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \tok.i1_4_lut_adj_44_LC_6_12_5  (
            .in0(N__16394),
            .in1(N__16316),
            .in2(N__16256),
            .in3(N__16252),
            .lcout(n10_adj_870),
            .ltout(n10_adj_870_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_85_LC_6_12_6 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_85_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_85_LC_6_12_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \tok.i26_3_lut_adj_85_LC_6_12_6  (
            .in0(_gnd_net_),
            .in1(N__16094),
            .in2(N__16223),
            .in3(N__16163),
            .lcout(\tok.tc_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i4_LC_6_12_7 .C_ON=1'b0;
    defparam \tok.tc_i4_LC_6_12_7 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i4_LC_6_12_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.tc_i4_LC_6_12_7  (
            .in0(N__16164),
            .in1(_gnd_net_),
            .in2(N__16104),
            .in3(N__16112),
            .lcout(tc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28536),
            .ce(),
            .sr(N__28174));
    defparam \tok.i5568_3_lut_LC_6_13_1 .C_ON=1'b0;
    defparam \tok.i5568_3_lut_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5568_3_lut_LC_6_13_1 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \tok.i5568_3_lut_LC_6_13_1  (
            .in0(N__28751),
            .in1(N__18083),
            .in2(_gnd_net_),
            .in3(N__23931),
            .lcout(\tok.n5571 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_40_LC_6_13_5 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_40_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_40_LC_6_13_5 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_40_LC_6_13_5  (
            .in0(N__16073),
            .in1(N__18334),
            .in2(N__17402),
            .in3(N__20230),
            .lcout(),
            .ltout(\tok.n83_adj_665_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5463_2_lut_3_lut_LC_6_13_6 .C_ON=1'b0;
    defparam \tok.i5463_2_lut_3_lut_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5463_2_lut_3_lut_LC_6_13_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i5463_2_lut_3_lut_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__19053),
            .in2(N__16037),
            .in3(N__30021),
            .lcout(\tok.n5487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i110_LC_7_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i110_LC_7_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i110_LC_7_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i110_LC_7_2_0  (
            .in0(N__17201),
            .in1(N__16024),
            .in2(_gnd_net_),
            .in3(N__26393),
            .lcout(tail_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28487),
            .ce(N__26047),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i94_LC_7_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i94_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i94_LC_7_2_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i94_LC_7_2_1  (
            .in0(N__26400),
            .in1(N__17215),
            .in2(_gnd_net_),
            .in3(N__16561),
            .lcout(\tok.A_stk.tail_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28487),
            .ce(N__26047),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i78_LC_7_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i78_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i78_LC_7_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i78_LC_7_2_2  (
            .in0(N__16025),
            .in1(N__16552),
            .in2(_gnd_net_),
            .in3(N__26399),
            .lcout(\tok.A_stk.tail_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28487),
            .ce(N__26047),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i62_LC_7_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i62_LC_7_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i62_LC_7_2_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i62_LC_7_2_3  (
            .in0(N__26398),
            .in1(N__16543),
            .in2(_gnd_net_),
            .in3(N__16562),
            .lcout(\tok.A_stk.tail_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28487),
            .ce(N__26047),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i46_LC_7_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i46_LC_7_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i46_LC_7_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i46_LC_7_2_4  (
            .in0(N__16534),
            .in1(N__16553),
            .in2(_gnd_net_),
            .in3(N__26397),
            .lcout(\tok.A_stk.tail_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28487),
            .ce(N__26047),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i30_LC_7_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i30_LC_7_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i30_LC_7_2_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i30_LC_7_2_5  (
            .in0(N__26396),
            .in1(N__25072),
            .in2(_gnd_net_),
            .in3(N__16544),
            .lcout(\tok.A_stk.tail_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28487),
            .ce(N__26047),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i14_LC_7_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i14_LC_7_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i14_LC_7_2_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i14_LC_7_2_6  (
            .in0(N__16535),
            .in1(N__26395),
            .in2(_gnd_net_),
            .in3(N__28868),
            .lcout(\tok.A_stk.tail_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28487),
            .ce(N__26047),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i111_LC_7_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i111_LC_7_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i111_LC_7_2_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i111_LC_7_2_7  (
            .in0(N__26394),
            .in1(N__16526),
            .in2(_gnd_net_),
            .in3(N__24667),
            .lcout(tail_111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28487),
            .ce(N__26047),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_140_LC_7_3_0 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_140_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_140_LC_7_3_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \tok.i50_4_lut_adj_140_LC_7_3_0  (
            .in0(N__16939),
            .in1(N__16505),
            .in2(N__16858),
            .in3(N__21143),
            .lcout(\tok.n27_adj_815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_69_LC_7_3_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_69_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_69_LC_7_3_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.i1_2_lut_adj_69_LC_7_3_1  (
            .in0(_gnd_net_),
            .in1(N__16498),
            .in2(_gnd_net_),
            .in3(N__16442),
            .lcout(),
            .ltout(\tok.depth_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_96_LC_7_3_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_96_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_96_LC_7_3_2 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \tok.i1_4_lut_adj_96_LC_7_3_2  (
            .in0(N__28582),
            .in1(N__16934),
            .in2(N__16412),
            .in3(N__16409),
            .lcout(\tok.n995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_144_LC_7_3_3 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_144_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_144_LC_7_3_3 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \tok.i50_4_lut_adj_144_LC_7_3_3  (
            .in0(N__22761),
            .in1(N__16848),
            .in2(N__16948),
            .in3(N__16400),
            .lcout(),
            .ltout(\tok.n27_adj_818_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i2_LC_7_3_4 .C_ON=1'b0;
    defparam \tok.idx_i2_LC_7_3_4 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i2_LC_7_3_4 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \tok.idx_i2_LC_7_3_4  (
            .in0(N__16975),
            .in1(N__16697),
            .in2(N__17009),
            .in3(N__16731),
            .lcout(\tok.idx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28494),
            .ce(),
            .sr(N__28232));
    defparam \tok.i50_4_lut_adj_148_LC_7_3_5 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_148_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_148_LC_7_3_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \tok.i50_4_lut_adj_148_LC_7_3_5  (
            .in0(N__16935),
            .in1(N__16865),
            .in2(N__29738),
            .in3(N__16849),
            .lcout(),
            .ltout(\tok.n27_adj_822_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i3_LC_7_3_6 .C_ON=1'b0;
    defparam \tok.idx_i3_LC_7_3_6 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i3_LC_7_3_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \tok.idx_i3_LC_7_3_6  (
            .in0(N__16770),
            .in1(N__16698),
            .in2(N__16805),
            .in3(N__16732),
            .lcout(\tok.idx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28494),
            .ce(),
            .sr(N__28232));
    defparam \tok.idx_i1_LC_7_3_7 .C_ON=1'b0;
    defparam \tok.idx_i1_LC_7_3_7 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i1_LC_7_3_7 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \tok.idx_i1_LC_7_3_7  (
            .in0(N__16730),
            .in1(N__16632),
            .in2(N__16703),
            .in3(N__16667),
            .lcout(\tok.idx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28494),
            .ce(),
            .sr(N__28232));
    defparam \tok.i567_2_lut_4_lut_LC_7_4_0 .C_ON=1'b0;
    defparam \tok.i567_2_lut_4_lut_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i567_2_lut_4_lut_LC_7_4_0 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \tok.i567_2_lut_4_lut_LC_7_4_0  (
            .in0(N__16586),
            .in1(N__17677),
            .in2(N__16598),
            .in3(N__19324),
            .lcout(rd_15__N_301),
            .ltout(rd_15__N_301_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i120_LC_7_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i120_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i120_LC_7_4_1 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \tok.A_stk.tail_i0_i120_LC_7_4_1  (
            .in0(N__26194),
            .in1(N__18616),
            .in2(N__16601),
            .in3(N__18596),
            .lcout(tail_120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28498),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i119_LC_7_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i119_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i119_LC_7_4_2 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i119_LC_7_4_2  (
            .in0(N__18653),
            .in1(N__25870),
            .in2(N__18682),
            .in3(N__26193),
            .lcout(tail_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28498),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2563_2_lut_4_lut_LC_7_4_3 .C_ON=1'b0;
    defparam \tok.i2563_2_lut_4_lut_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2563_2_lut_4_lut_LC_7_4_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \tok.i2563_2_lut_4_lut_LC_7_4_3  (
            .in0(N__19323),
            .in1(N__16594),
            .in2(N__17678),
            .in3(N__16585),
            .lcout(A_stk_delta_1),
            .ltout(A_stk_delta_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i117_LC_7_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i117_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i117_LC_7_4_4 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \tok.A_stk.tail_i0_i117_LC_7_4_4  (
            .in0(N__24914),
            .in1(N__24925),
            .in2(N__16565),
            .in3(N__25869),
            .lcout(tail_117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28498),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i121_LC_7_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i121_LC_7_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i121_LC_7_4_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \tok.A_stk.tail_i0_i121_LC_7_4_5  (
            .in0(N__26195),
            .in1(N__18481),
            .in2(N__25926),
            .in3(N__18470),
            .lcout(tail_121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28498),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i115_LC_7_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i115_LC_7_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i115_LC_7_4_6 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i115_LC_7_4_6  (
            .in0(N__18536),
            .in1(N__25868),
            .in2(N__18551),
            .in3(N__26192),
            .lcout(tail_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28498),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i126_LC_7_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i126_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i126_LC_7_4_7 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \tok.A_stk.tail_i0_i126_LC_7_4_7  (
            .in0(N__26196),
            .in1(N__17219),
            .in2(N__25927),
            .in3(N__17197),
            .lcout(tail_126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28498),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i95_LC_7_5_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i95_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i95_LC_7_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i95_LC_7_5_0  (
            .in0(N__17176),
            .in1(N__24641),
            .in2(_gnd_net_),
            .in3(N__26246),
            .lcout(\tok.A_stk.tail_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28505),
            .ce(N__26020),
            .sr(_gnd_net_));
    defparam \tok.or_99_i9_2_lut_3_lut_LC_7_5_2 .C_ON=1'b0;
    defparam \tok.or_99_i9_2_lut_3_lut_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i9_2_lut_3_lut_LC_7_5_2 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \tok.or_99_i9_2_lut_3_lut_LC_7_5_2  (
            .in0(N__22170),
            .in1(N__29586),
            .in2(_gnd_net_),
            .in3(N__22144),
            .lcout(\tok.n181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i2_3_lut_adj_28_LC_7_5_6 .C_ON=1'b0;
    defparam \tok.uart.i2_3_lut_adj_28_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_3_lut_adj_28_LC_7_5_6 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \tok.uart.i2_3_lut_adj_28_LC_7_5_6  (
            .in0(N__17077),
            .in1(_gnd_net_),
            .in2(N__17111),
            .in3(N__17158),
            .lcout(\tok.uart.n5235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i5204_2_lut_LC_7_5_7 .C_ON=1'b0;
    defparam \tok.uart.i5204_2_lut_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5204_2_lut_LC_7_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.uart.i5204_2_lut_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(N__17107),
            .in2(_gnd_net_),
            .in3(N__17076),
            .lcout(\tok.uart.n5374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.key_rd_15__I_0_241_i14_2_lut_LC_7_6_0 .C_ON=1'b0;
    defparam \tok.key_rd_15__I_0_241_i14_2_lut_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.key_rd_15__I_0_241_i14_2_lut_LC_7_6_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.key_rd_15__I_0_241_i14_2_lut_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__17035),
            .in2(_gnd_net_),
            .in3(N__23157),
            .lcout(\tok.n14_adj_647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i0_LC_7_6_1 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i0_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i0_LC_7_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.uart.rx_data_i0_i0_LC_7_6_1  (
            .in0(N__25661),
            .in1(N__17306),
            .in2(_gnd_net_),
            .in3(N__17293),
            .lcout(uart_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28511),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i0_LC_7_6_4 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i0_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i0_LC_7_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i0_LC_7_6_4  (
            .in0(N__17305),
            .in1(N__17320),
            .in2(_gnd_net_),
            .in3(N__22973),
            .lcout(capture_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28511),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i1_LC_7_6_5 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i1_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i1_LC_7_6_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.uart.capture_i0_i1_LC_7_6_5  (
            .in0(N__22974),
            .in1(N__17304),
            .in2(_gnd_net_),
            .in3(N__21184),
            .lcout(capture_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28511),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_125_LC_7_6_6 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_125_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_125_LC_7_6_6 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \tok.i2_4_lut_adj_125_LC_7_6_6  (
            .in0(N__23410),
            .in1(N__29469),
            .in2(N__17294),
            .in3(N__23334),
            .lcout(),
            .ltout(\tok.n6_adj_794_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_159_LC_7_6_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_159_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_159_LC_7_6_7 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \tok.i1_4_lut_adj_159_LC_7_6_7  (
            .in0(N__22781),
            .in1(N__20477),
            .in2(N__17282),
            .in3(N__22550),
            .lcout(\tok.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_5_i3_3_lut_LC_7_7_0 .C_ON=1'b0;
    defparam \tok.select_73_Select_5_i3_3_lut_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_5_i3_3_lut_LC_7_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \tok.select_73_Select_5_i3_3_lut_LC_7_7_0  (
            .in0(N__28949),
            .in1(N__27754),
            .in2(_gnd_net_),
            .in3(N__18818),
            .lcout(\tok.n3_adj_859 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5577_4_lut_LC_7_7_1 .C_ON=1'b0;
    defparam \tok.i5577_4_lut_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5577_4_lut_LC_7_7_1 .LUT_INIT=16'b1111000011110110;
    LogicCell40 \tok.i5577_4_lut_LC_7_7_1  (
            .in0(N__21111),
            .in1(N__19259),
            .in2(N__19430),
            .in3(N__28950),
            .lcout(),
            .ltout(\tok.n5553_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5576_4_lut_LC_7_7_2 .C_ON=1'b0;
    defparam \tok.i5576_4_lut_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5576_4_lut_LC_7_7_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i5576_4_lut_LC_7_7_2  (
            .in0(N__17275),
            .in1(N__23573),
            .in2(N__17249),
            .in3(N__26973),
            .lcout(\tok.n5552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_adj_111_LC_7_7_3 .C_ON=1'b0;
    defparam \tok.i3_3_lut_adj_111_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_adj_111_LC_7_7_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \tok.i3_3_lut_adj_111_LC_7_7_3  (
            .in0(N__26974),
            .in1(N__17246),
            .in2(_gnd_net_),
            .in3(N__19613),
            .lcout(\tok.n15_adj_770 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_adj_84_LC_7_7_4 .C_ON=1'b0;
    defparam \tok.i3_3_lut_adj_84_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_adj_84_LC_7_7_4 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \tok.i3_3_lut_adj_84_LC_7_7_4  (
            .in0(N__17234),
            .in1(N__26972),
            .in2(_gnd_net_),
            .in3(N__19625),
            .lcout(),
            .ltout(\tok.n14_adj_735_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_91_LC_7_7_5 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_91_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_91_LC_7_7_5 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \tok.i7_4_lut_adj_91_LC_7_7_5  (
            .in0(N__27940),
            .in1(N__20798),
            .in2(N__17423),
            .in3(N__29598),
            .lcout(\tok.n18_adj_739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_99_i6_3_lut_LC_7_7_6 .C_ON=1'b0;
    defparam \tok.or_99_i6_3_lut_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i6_3_lut_LC_7_7_6 .LUT_INIT=16'b1111111101100110;
    LogicCell40 \tok.or_99_i6_3_lut_LC_7_7_6  (
            .in0(N__19049),
            .in1(N__18817),
            .in2(_gnd_net_),
            .in3(N__21110),
            .lcout(\tok.n184 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_100_LC_7_7_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_100_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_100_LC_7_7_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \tok.i1_2_lut_adj_100_LC_7_7_7  (
            .in0(N__18816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19048),
            .lcout(\tok.n6_adj_754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_185_LC_7_8_0 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_185_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_185_LC_7_8_0 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \tok.i2_4_lut_adj_185_LC_7_8_0  (
            .in0(N__27850),
            .in1(N__20642),
            .in2(N__29608),
            .in3(N__27633),
            .lcout(\tok.n13_adj_852 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_adj_184_LC_7_8_1 .C_ON=1'b0;
    defparam \tok.i5_3_lut_adj_184_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_adj_184_LC_7_8_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i5_3_lut_adj_184_LC_7_8_1  (
            .in0(N__17401),
            .in1(N__23696),
            .in2(_gnd_net_),
            .in3(N__26954),
            .lcout(),
            .ltout(\tok.n16_adj_851_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5507_4_lut_LC_7_8_2 .C_ON=1'b0;
    defparam \tok.i5507_4_lut_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5507_4_lut_LC_7_8_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i5507_4_lut_LC_7_8_2  (
            .in0(N__19037),
            .in1(N__19442),
            .in2(N__17375),
            .in3(N__28971),
            .lcout(),
            .ltout(\tok.n5562_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5569_4_lut_LC_7_8_3 .C_ON=1'b0;
    defparam \tok.i5569_4_lut_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5569_4_lut_LC_7_8_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i5569_4_lut_LC_7_8_3  (
            .in0(N__17372),
            .in1(N__17351),
            .in2(N__17360),
            .in3(N__17357),
            .lcout(\tok.n5561 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_4_lut_adj_187_LC_7_8_4 .C_ON=1'b0;
    defparam \tok.i3_4_lut_4_lut_adj_187_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_4_lut_adj_187_LC_7_8_4 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \tok.i3_4_lut_4_lut_adj_187_LC_7_8_4  (
            .in0(N__23776),
            .in1(N__17825),
            .in2(N__28762),
            .in3(N__29149),
            .lcout(\tok.n14_adj_854 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i2_LC_7_8_7 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i2_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i2_LC_7_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.uart.rx_data_i0_i2_LC_7_8_7  (
            .in0(N__17345),
            .in1(N__23365),
            .in2(_gnd_net_),
            .in3(N__25681),
            .lcout(uart_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28524),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5570_4_lut_LC_7_9_0 .C_ON=1'b0;
    defparam \tok.i5570_4_lut_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5570_4_lut_LC_7_9_0 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \tok.i5570_4_lut_LC_7_9_0  (
            .in0(N__19349),
            .in1(N__26960),
            .in2(N__17570),
            .in3(N__20012),
            .lcout(),
            .ltout(\tok.n5463_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5555_4_lut_LC_7_9_1 .C_ON=1'b0;
    defparam \tok.i5555_4_lut_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5555_4_lut_LC_7_9_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i5555_4_lut_LC_7_9_1  (
            .in0(N__19913),
            .in1(N__17543),
            .in2(N__17534),
            .in3(N__27563),
            .lcout(\tok.n5462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_109_LC_7_9_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_109_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_109_LC_7_9_2 .LUT_INIT=16'b0101010101011101;
    LogicCell40 \tok.i1_4_lut_adj_109_LC_7_9_2  (
            .in0(N__29148),
            .in1(N__17530),
            .in2(N__17638),
            .in3(N__17491),
            .lcout(\tok.n8_adj_767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_215_i15_2_lut_3_lut_LC_7_9_3 .C_ON=1'b0;
    defparam \tok.T_7__I_0_215_i15_2_lut_3_lut_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_215_i15_2_lut_3_lut_LC_7_9_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.T_7__I_0_215_i15_2_lut_3_lut_LC_7_9_3  (
            .in0(N__18421),
            .in1(N__19693),
            .in2(_gnd_net_),
            .in3(N__19050),
            .lcout(\tok.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5170_2_lut_LC_7_9_4 .C_ON=1'b0;
    defparam \tok.i5170_2_lut_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5170_2_lut_LC_7_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i5170_2_lut_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__26710),
            .in2(_gnd_net_),
            .in3(N__28904),
            .lcout(\tok.n5334 ),
            .ltout(\tok.n5334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_166_LC_7_9_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_166_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_166_LC_7_9_5 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \tok.i1_4_lut_adj_166_LC_7_9_5  (
            .in0(N__26959),
            .in1(N__17458),
            .in2(N__17426),
            .in3(N__18335),
            .lcout(\tok.n8_adj_837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_181_LC_7_9_6 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_181_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_181_LC_7_9_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i1_2_lut_adj_181_LC_7_9_6  (
            .in0(N__19051),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18422),
            .lcout(\tok.n14_adj_679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i2_1_lut_LC_7_9_7 .C_ON=1'b0;
    defparam \tok.inv_106_i2_1_lut_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i2_1_lut_LC_7_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i2_1_lut_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21103),
            .lcout(\tok.n301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i11_LC_7_10_0 .C_ON=1'b0;
    defparam \tok.A_i11_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \tok.A_i11_LC_7_10_0 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \tok.A_i11_LC_7_10_0  (
            .in0(N__27452),
            .in1(N__26858),
            .in2(N__28636),
            .in3(N__19919),
            .lcout(\tok.A_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28532),
            .ce(N__28285),
            .sr(N__28192));
    defparam \tok.A_i12_LC_7_10_1 .C_ON=1'b0;
    defparam \tok.A_i12_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \tok.A_i12_LC_7_10_1 .LUT_INIT=16'b1111011111000100;
    LogicCell40 \tok.A_i12_LC_7_10_1  (
            .in0(N__26859),
            .in1(N__28618),
            .in2(N__20942),
            .in3(N__25061),
            .lcout(\tok.A_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28532),
            .ce(N__28285),
            .sr(N__28192));
    defparam \tok.A_i1_LC_7_10_2 .C_ON=1'b0;
    defparam \tok.A_i1_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \tok.A_i1_LC_7_10_2 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \tok.A_i1_LC_7_10_2  (
            .in0(N__28619),
            .in1(N__26860),
            .in2(N__17663),
            .in3(N__22886),
            .lcout(\tok.A_low_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28532),
            .ce(N__28285),
            .sr(N__28192));
    defparam \tok.A_i2_LC_7_10_3 .C_ON=1'b0;
    defparam \tok.A_i2_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \tok.A_i2_LC_7_10_3 .LUT_INIT=16'b1100111110101010;
    LogicCell40 \tok.A_i2_LC_7_10_3  (
            .in0(N__24031),
            .in1(N__19517),
            .in2(N__26869),
            .in3(N__28620),
            .lcout(\tok.A_low_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28532),
            .ce(N__28285),
            .sr(N__28192));
    defparam \tok.A_i3_LC_7_10_4 .C_ON=1'b0;
    defparam \tok.A_i3_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \tok.A_i3_LC_7_10_4 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \tok.A_i3_LC_7_10_4  (
            .in0(N__23924),
            .in1(N__26864),
            .in2(N__28637),
            .in3(N__19760),
            .lcout(\tok.A_low_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28532),
            .ce(N__28285),
            .sr(N__28192));
    defparam \tok.A_i4_LC_7_10_5 .C_ON=1'b0;
    defparam \tok.A_i4_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \tok.A_i4_LC_7_10_5 .LUT_INIT=16'b1110111000101110;
    LogicCell40 \tok.A_i4_LC_7_10_5  (
            .in0(N__25374),
            .in1(N__28624),
            .in2(N__26870),
            .in3(N__17654),
            .lcout(\tok.A_low_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28532),
            .ce(N__28285),
            .sr(N__28192));
    defparam \tok.A_i5_LC_7_10_6 .C_ON=1'b0;
    defparam \tok.A_i5_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \tok.A_i5_LC_7_10_6 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \tok.A_i5_LC_7_10_6  (
            .in0(N__28625),
            .in1(N__26868),
            .in2(N__23794),
            .in3(N__17648),
            .lcout(\tok.A_low_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28532),
            .ce(N__28285),
            .sr(N__28192));
    defparam \tok.i2_4_lut_LC_7_10_7 .C_ON=1'b0;
    defparam \tok.i2_4_lut_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_LC_7_10_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i2_4_lut_LC_7_10_7  (
            .in0(N__24030),
            .in1(N__29545),
            .in2(N__23792),
            .in3(N__21084),
            .lcout(\tok.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i7_1_lut_LC_7_11_0 .C_ON=1'b0;
    defparam \tok.inv_106_i7_1_lut_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i7_1_lut_LC_7_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i7_1_lut_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21867),
            .lcout(\tok.n296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_110_LC_7_11_1 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_110_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_110_LC_7_11_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i2_3_lut_adj_110_LC_7_11_1  (
            .in0(N__21868),
            .in1(N__20783),
            .in2(_gnd_net_),
            .in3(N__27914),
            .lcout(\tok.n14_adj_769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_220_i15_2_lut_3_lut_LC_7_11_2 .C_ON=1'b0;
    defparam \tok.T_7__I_0_220_i15_2_lut_3_lut_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_220_i15_2_lut_3_lut_LC_7_11_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.T_7__I_0_220_i15_2_lut_3_lut_LC_7_11_2  (
            .in0(N__17639),
            .in1(N__22480),
            .in2(_gnd_net_),
            .in3(N__17615),
            .lcout(\tok.n15_adj_655 ),
            .ltout(\tok.n15_adj_655_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_135_LC_7_11_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_135_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_135_LC_7_11_3 .LUT_INIT=16'b0000110001011101;
    LogicCell40 \tok.i1_4_lut_adj_135_LC_7_11_3  (
            .in0(N__17745),
            .in1(N__17813),
            .in2(N__17774),
            .in3(N__27913),
            .lcout(\tok.uart_stall ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.valid_54_LC_7_11_4 .C_ON=1'b0;
    defparam \tok.uart.valid_54_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.valid_54_LC_7_11_4 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \tok.uart.valid_54_LC_7_11_4  (
            .in0(N__17749),
            .in1(N__22481),
            .in2(_gnd_net_),
            .in3(N__23308),
            .lcout(\tok.uart_rx_valid ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28537),
            .ce(N__17732),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_3_lut_4_lut_LC_7_11_5 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_3_lut_4_lut_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_3_lut_4_lut_LC_7_11_5 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \tok.uart.i1_2_lut_3_lut_4_lut_LC_7_11_5  (
            .in0(N__23307),
            .in1(N__25688),
            .in2(N__17750),
            .in3(N__22485),
            .lcout(\tok.uart.n953 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_233_i15_2_lut_LC_7_11_6 .C_ON=1'b0;
    defparam \tok.T_7__I_0_233_i15_2_lut_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_233_i15_2_lut_LC_7_11_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.T_7__I_0_233_i15_2_lut_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__22479),
            .in2(_gnd_net_),
            .in3(N__23306),
            .lcout(\tok.n15_adj_667 ),
            .ltout(\tok.n15_adj_667_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_117_LC_7_11_7 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_117_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_117_LC_7_11_7 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \tok.i2_4_lut_adj_117_LC_7_11_7  (
            .in0(N__22303),
            .in1(N__24861),
            .in2(N__17723),
            .in3(N__27649),
            .lcout(\tok.n13_adj_780 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_171_LC_7_12_0 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_171_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_171_LC_7_12_0 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \tok.i3_4_lut_adj_171_LC_7_12_0  (
            .in0(N__30019),
            .in1(N__26975),
            .in2(N__17720),
            .in3(N__26762),
            .lcout(\tok.n11_adj_840 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_LC_7_12_1 .C_ON=1'b0;
    defparam \tok.i2_2_lut_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_LC_7_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i2_2_lut_LC_7_12_1  (
            .in0(N__18358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30018),
            .lcout(),
            .ltout(\tok.n28_adj_771_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5446_4_lut_LC_7_12_2 .C_ON=1'b0;
    defparam \tok.i5446_4_lut_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5446_4_lut_LC_7_12_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \tok.i5446_4_lut_LC_7_12_2  (
            .in0(N__20270),
            .in1(N__19046),
            .in2(N__17690),
            .in3(N__18021),
            .lcout(),
            .ltout(\tok.n5467_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i49_4_lut_LC_7_12_3 .C_ON=1'b0;
    defparam \tok.i49_4_lut_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i49_4_lut_LC_7_12_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.i49_4_lut_LC_7_12_3  (
            .in0(N__19047),
            .in1(N__17687),
            .in2(N__17681),
            .in3(N__19244),
            .lcout(\tok.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2626_1_lut_LC_7_12_4 .C_ON=1'b0;
    defparam \tok.i2626_1_lut_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2626_1_lut_LC_7_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.i2626_1_lut_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29119),
            .lcout(\tok.n82 ),
            .ltout(\tok.n82_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_2_lut_LC_7_12_5 .C_ON=1'b0;
    defparam \tok.sub_100_add_2_2_lut_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_2_lut_LC_7_12_5 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \tok.sub_100_add_2_2_lut_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__24190),
            .in2(N__18425),
            .in3(N__20271),
            .lcout(\tok.n14_adj_764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2625_2_lut_3_lut_LC_7_12_6 .C_ON=1'b0;
    defparam \tok.i2625_2_lut_3_lut_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2625_2_lut_3_lut_LC_7_12_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i2625_2_lut_3_lut_LC_7_12_6  (
            .in0(N__19738),
            .in1(N__18414),
            .in2(_gnd_net_),
            .in3(N__19045),
            .lcout(\tok.n2703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_178_LC_7_12_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_178_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_178_LC_7_12_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i1_2_lut_adj_178_LC_7_12_7  (
            .in0(N__19457),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17837),
            .lcout(\tok.n8_adj_846 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_80_LC_7_13_0 .C_ON=1'b1;
    defparam \tok.i1_2_lut_adj_80_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_80_LC_7_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i1_2_lut_adj_80_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__20229),
            .in2(_gnd_net_),
            .in3(N__18318),
            .lcout(\tok.n41 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\tok.n4761 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_3_lut_LC_7_13_1 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_3_lut_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_3_lut_LC_7_13_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_100_add_2_3_lut_LC_7_13_1  (
            .in0(N__18072),
            .in1(_gnd_net_),
            .in2(N__18353),
            .in3(N__18086),
            .lcout(\tok.n23_adj_718 ),
            .ltout(),
            .carryin(\tok.n4761 ),
            .carryout(\tok.n4762 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_4_lut_LC_7_13_2 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_4_lut_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_4_lut_LC_7_13_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_100_add_2_4_lut_LC_7_13_2  (
            .in0(N__18074),
            .in1(N__30017),
            .in2(_gnd_net_),
            .in3(N__18077),
            .lcout(\tok.n15_adj_664 ),
            .ltout(),
            .carryin(\tok.n4762 ),
            .carryout(\tok.n4763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_5_lut_LC_7_13_3 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_5_lut_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_5_lut_LC_7_13_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_100_add_2_5_lut_LC_7_13_3  (
            .in0(N__18073),
            .in1(N__18025),
            .in2(N__24219),
            .in3(N__17828),
            .lcout(\tok.n11_adj_830 ),
            .ltout(),
            .carryin(\tok.n4763 ),
            .carryout(\tok.n4764 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_6_lut_LC_7_13_4 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_6_lut_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_6_lut_LC_7_13_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_100_add_2_6_lut_LC_7_13_4  (
            .in0(N__27725),
            .in1(N__19052),
            .in2(_gnd_net_),
            .in3(N__17816),
            .lcout(\tok.n212 ),
            .ltout(),
            .carryin(\tok.n4764 ),
            .carryout(\tok.n4765 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_7_lut_LC_7_13_5 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_7_lut_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_7_lut_LC_7_13_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_100_add_2_7_lut_LC_7_13_5  (
            .in0(N__21115),
            .in1(N__18804),
            .in2(_gnd_net_),
            .in3(N__18512),
            .lcout(\tok.n211 ),
            .ltout(),
            .carryin(\tok.n4765 ),
            .carryout(\tok.n4766 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_8_lut_LC_7_13_6 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_8_lut_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_8_lut_LC_7_13_6 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_100_add_2_8_lut_LC_7_13_6  (
            .in0(N__22750),
            .in1(N__19214),
            .in2(N__24209),
            .in3(N__18494),
            .lcout(\tok.n210 ),
            .ltout(),
            .carryin(\tok.n4766 ),
            .carryout(\tok.n4767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_9_lut_LC_7_13_7 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_9_lut_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_9_lut_LC_7_13_7 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_100_add_2_9_lut_LC_7_13_7  (
            .in0(N__29702),
            .in1(N__22110),
            .in2(N__24220),
            .in3(N__18491),
            .lcout(\tok.n209 ),
            .ltout(),
            .carryin(\tok.n4767 ),
            .carryout(\tok.n4768 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_10_lut_LC_7_14_0 .C_ON=1'b0;
    defparam \tok.sub_100_add_2_10_lut_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_10_lut_LC_7_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_100_add_2_10_lut_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__24189),
            .in2(_gnd_net_),
            .in3(N__18488),
            .lcout(\tok.n191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i105_LC_8_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i105_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i105_LC_8_2_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i105_LC_8_2_0  (
            .in0(N__26408),
            .in1(N__18485),
            .in2(_gnd_net_),
            .in3(N__18451),
            .lcout(tail_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28495),
            .ce(N__26048),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i89_LC_8_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i89_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i89_LC_8_2_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i89_LC_8_2_1  (
            .in0(N__18463),
            .in1(N__18442),
            .in2(_gnd_net_),
            .in3(N__26413),
            .lcout(\tok.A_stk.tail_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28495),
            .ce(N__26048),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i73_LC_8_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i73_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i73_LC_8_2_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i73_LC_8_2_2  (
            .in0(N__26412),
            .in1(N__18452),
            .in2(_gnd_net_),
            .in3(N__18433),
            .lcout(\tok.A_stk.tail_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28495),
            .ce(N__26048),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i57_LC_8_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i57_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i57_LC_8_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i57_LC_8_2_3  (
            .in0(N__18580),
            .in1(N__18443),
            .in2(_gnd_net_),
            .in3(N__26411),
            .lcout(\tok.A_stk.tail_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28495),
            .ce(N__26048),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i41_LC_8_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i41_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i41_LC_8_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i41_LC_8_2_4  (
            .in0(N__26410),
            .in1(N__18571),
            .in2(_gnd_net_),
            .in3(N__18434),
            .lcout(\tok.A_stk.tail_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28495),
            .ce(N__26048),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i25_LC_8_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i25_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i25_LC_8_2_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \tok.A_stk.tail_i0_i25_LC_8_2_5  (
            .in0(N__18581),
            .in1(_gnd_net_),
            .in2(N__18563),
            .in3(N__26409),
            .lcout(\tok.A_stk.tail_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28495),
            .ce(N__26048),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i9_LC_8_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i9_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i9_LC_8_2_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i9_LC_8_2_6  (
            .in0(N__26414),
            .in1(N__18572),
            .in2(_gnd_net_),
            .in3(N__27513),
            .lcout(\tok.A_stk.tail_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28495),
            .ce(N__26048),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i9_LC_8_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i9_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i9_LC_8_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i9_LC_8_2_7  (
            .in0(N__18559),
            .in1(N__25473),
            .in2(_gnd_net_),
            .in3(N__29081),
            .lcout(\tok.S_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28495),
            .ce(N__26048),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i99_LC_8_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i99_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i99_LC_8_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i99_LC_8_3_0  (
            .in0(N__26286),
            .in1(N__18550),
            .in2(_gnd_net_),
            .in3(N__20560),
            .lcout(tail_99),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28499),
            .ce(N__26061),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i83_LC_8_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i83_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i83_LC_8_3_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i83_LC_8_3_1  (
            .in0(N__26623),
            .in1(N__18535),
            .in2(_gnd_net_),
            .in3(N__26284),
            .lcout(\tok.A_stk.tail_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28499),
            .ce(N__26061),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i20_LC_8_3_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i20_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i20_LC_8_3_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i20_LC_8_3_2  (
            .in0(N__26280),
            .in1(N__18692),
            .in2(_gnd_net_),
            .in3(N__20548),
            .lcout(\tok.A_stk.tail_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28499),
            .ce(N__26061),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i100_LC_8_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i100_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i100_LC_8_3_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i100_LC_8_3_3  (
            .in0(N__20453),
            .in1(N__18523),
            .in2(_gnd_net_),
            .in3(N__26279),
            .lcout(tail_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28499),
            .ce(N__26061),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i84_LC_8_3_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i84_LC_8_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i84_LC_8_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i84_LC_8_3_4  (
            .in0(N__26285),
            .in1(N__20464),
            .in2(_gnd_net_),
            .in3(N__18709),
            .lcout(\tok.A_stk.tail_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28499),
            .ce(N__26061),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i68_LC_8_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i68_LC_8_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i68_LC_8_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i68_LC_8_3_5  (
            .in0(N__18524),
            .in1(N__18700),
            .in2(_gnd_net_),
            .in3(N__26283),
            .lcout(\tok.A_stk.tail_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28499),
            .ce(N__26061),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i52_LC_8_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i52_LC_8_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i52_LC_8_3_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i52_LC_8_3_6  (
            .in0(N__26282),
            .in1(N__18691),
            .in2(_gnd_net_),
            .in3(N__18710),
            .lcout(\tok.A_stk.tail_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28499),
            .ce(N__26061),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i36_LC_8_3_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i36_LC_8_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i36_LC_8_3_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i36_LC_8_3_7  (
            .in0(N__18664),
            .in1(N__18701),
            .in2(_gnd_net_),
            .in3(N__26281),
            .lcout(\tok.A_stk.tail_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28499),
            .ce(N__26061),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i103_LC_8_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i103_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i103_LC_8_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i103_LC_8_4_0  (
            .in0(N__18683),
            .in1(N__18628),
            .in2(_gnd_net_),
            .in3(N__26238),
            .lcout(tail_103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28506),
            .ce(N__25968),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i55_LC_8_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i55_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i55_LC_8_4_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i55_LC_8_4_1  (
            .in0(N__26241),
            .in1(_gnd_net_),
            .in2(N__18641),
            .in3(N__20575),
            .lcout(\tok.A_stk.tail_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28506),
            .ce(N__25968),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i71_LC_8_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i71_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i71_LC_8_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i71_LC_8_4_2  (
            .in0(N__18629),
            .in1(N__20587),
            .in2(_gnd_net_),
            .in3(N__26242),
            .lcout(\tok.A_stk.tail_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28506),
            .ce(N__25968),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i88_LC_8_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i88_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i88_LC_8_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i88_LC_8_4_3  (
            .in0(N__26245),
            .in1(N__18592),
            .in2(_gnd_net_),
            .in3(N__20392),
            .lcout(\tok.A_stk.tail_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28506),
            .ce(N__25968),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i4_LC_8_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i4_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i4_LC_8_4_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i4_LC_8_4_4  (
            .in0(N__18665),
            .in1(N__26240),
            .in2(_gnd_net_),
            .in3(N__23742),
            .lcout(\tok.A_stk.tail_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28506),
            .ce(N__25968),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i72_LC_8_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i72_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i72_LC_8_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i72_LC_8_4_5  (
            .in0(N__26243),
            .in1(N__18605),
            .in2(_gnd_net_),
            .in3(N__21988),
            .lcout(\tok.A_stk.tail_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28506),
            .ce(N__25968),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i87_LC_8_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i87_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i87_LC_8_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i87_LC_8_4_6  (
            .in0(N__18652),
            .in1(N__18637),
            .in2(_gnd_net_),
            .in3(N__26244),
            .lcout(\tok.A_stk.tail_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28506),
            .ce(N__25968),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i104_LC_8_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i104_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i104_LC_8_4_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i104_LC_8_4_7  (
            .in0(N__26239),
            .in1(N__18617),
            .in2(_gnd_net_),
            .in3(N__18604),
            .lcout(tail_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28506),
            .ce(N__25968),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_123_LC_8_5_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_123_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_123_LC_8_5_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.i1_2_lut_adj_123_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__18830),
            .in2(_gnd_net_),
            .in3(N__22141),
            .lcout(\tok.n9_adj_786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5447_4_lut_LC_8_5_1 .C_ON=1'b0;
    defparam \tok.i5447_4_lut_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5447_4_lut_LC_8_5_1 .LUT_INIT=16'b1111000011110110;
    LogicCell40 \tok.i5447_4_lut_LC_8_5_1  (
            .in0(N__22143),
            .in1(N__22760),
            .in2(N__19418),
            .in3(N__28978),
            .lcout(),
            .ltout(\tok.n5548_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5445_4_lut_LC_8_5_2 .C_ON=1'b0;
    defparam \tok.i5445_4_lut_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5445_4_lut_LC_8_5_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i5445_4_lut_LC_8_5_2  (
            .in0(N__19307),
            .in1(N__23432),
            .in2(N__19283),
            .in3(N__26994),
            .lcout(\tok.n5547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i227_2_lut_LC_8_5_3 .C_ON=1'b0;
    defparam \tok.i227_2_lut_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i227_2_lut_LC_8_5_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \tok.i227_2_lut_LC_8_5_3  (
            .in0(N__18832),
            .in1(_gnd_net_),
            .in2(N__19073),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\tok.n285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_6_i1_4_lut_LC_8_5_4 .C_ON=1'b0;
    defparam \tok.select_73_Select_6_i1_4_lut_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_6_i1_4_lut_LC_8_5_4 .LUT_INIT=16'b0000000011101101;
    LogicCell40 \tok.select_73_Select_6_i1_4_lut_LC_8_5_4  (
            .in0(N__19238),
            .in1(N__22759),
            .in2(N__19280),
            .in3(N__26763),
            .lcout(),
            .ltout(\tok.n1_adj_862_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_199_LC_8_5_5 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_199_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_199_LC_8_5_5 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \tok.i6_4_lut_adj_199_LC_8_5_5  (
            .in0(N__19277),
            .in1(N__23213),
            .in2(N__19262),
            .in3(N__25771),
            .lcout(\tok.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i237_2_lut_3_lut_LC_8_5_6 .C_ON=1'b0;
    defparam \tok.i237_2_lut_3_lut_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i237_2_lut_3_lut_LC_8_5_6 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \tok.i237_2_lut_3_lut_LC_8_5_6  (
            .in0(N__19237),
            .in1(N__19066),
            .in2(_gnd_net_),
            .in3(N__18831),
            .lcout(\tok.n6_adj_650 ),
            .ltout(\tok.n6_adj_650_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i245_2_lut_LC_8_5_7 .C_ON=1'b0;
    defparam \tok.i245_2_lut_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i245_2_lut_LC_8_5_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \tok.i245_2_lut_LC_8_5_7  (
            .in0(N__22142),
            .in1(_gnd_net_),
            .in2(N__18713),
            .in3(_gnd_net_),
            .lcout(\tok.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_35_LC_8_6_1 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_35_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_35_LC_8_6_1 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \tok.i2_4_lut_adj_35_LC_8_6_1  (
            .in0(N__27652),
            .in1(N__20615),
            .in2(N__22313),
            .in3(N__27882),
            .lcout(),
            .ltout(\tok.n13_adj_654_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5578_4_lut_LC_8_6_2 .C_ON=1'b0;
    defparam \tok.i5578_4_lut_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5578_4_lut_LC_8_6_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i5578_4_lut_LC_8_6_2  (
            .in0(N__20351),
            .in1(N__20927),
            .in2(N__19391),
            .in3(N__19388),
            .lcout(),
            .ltout(\tok.n5546_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i8_LC_8_6_3 .C_ON=1'b0;
    defparam \tok.A_i8_LC_8_6_3 .SEQ_MODE=4'b1010;
    defparam \tok.A_i8_LC_8_6_3 .LUT_INIT=16'b1111011111000100;
    LogicCell40 \tok.A_i8_LC_8_6_3  (
            .in0(N__26828),
            .in1(N__28589),
            .in2(N__19382),
            .in3(N__23543),
            .lcout(A_low_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28518),
            .ce(N__28300),
            .sr(N__28205));
    defparam \tok.i2_4_lut_adj_195_LC_8_6_4 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_195_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_195_LC_8_6_4 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \tok.i2_4_lut_adj_195_LC_8_6_4  (
            .in0(N__21834),
            .in1(N__20624),
            .in2(N__27887),
            .in3(N__27651),
            .lcout(),
            .ltout(\tok.n13_adj_641_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5582_4_lut_LC_8_6_5 .C_ON=1'b0;
    defparam \tok.i5582_4_lut_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i5582_4_lut_LC_8_6_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i5582_4_lut_LC_8_6_5  (
            .in0(N__19379),
            .in1(N__19367),
            .in2(N__19361),
            .in3(N__19358),
            .lcout(),
            .ltout(\tok.n5551_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i7_LC_8_6_6 .C_ON=1'b0;
    defparam \tok.A_i7_LC_8_6_6 .SEQ_MODE=4'b1010;
    defparam \tok.A_i7_LC_8_6_6 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \tok.A_i7_LC_8_6_6  (
            .in0(N__28588),
            .in1(N__26827),
            .in2(N__19352),
            .in3(N__23633),
            .lcout(\tok.A_low_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28518),
            .ce(N__28300),
            .sr(N__28205));
    defparam \tok.add_104_2_lut_LC_8_7_0 .C_ON=1'b1;
    defparam \tok.add_104_2_lut_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_2_lut_LC_8_7_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \tok.add_104_2_lut_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__27738),
            .in2(N__22880),
            .in3(N__19598),
            .lcout(\tok.n5465 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\tok.n4784 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_3_lut_LC_8_7_1 .C_ON=1'b1;
    defparam \tok.add_104_3_lut_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_3_lut_LC_8_7_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_3_lut_LC_8_7_1  (
            .in0(N__19595),
            .in1(N__21107),
            .in2(N__24035),
            .in3(N__19340),
            .lcout(\tok.n17_adj_812 ),
            .ltout(),
            .carryin(\tok.n4784 ),
            .carryout(\tok.n4785 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_4_lut_LC_8_7_2 .C_ON=1'b1;
    defparam \tok.add_104_4_lut_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_4_lut_LC_8_7_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_4_lut_LC_8_7_2  (
            .in0(N__19591),
            .in1(N__22732),
            .in2(N__23920),
            .in3(N__19337),
            .lcout(\tok.n16_adj_810 ),
            .ltout(),
            .carryin(\tok.n4785 ),
            .carryout(\tok.n4786 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_5_lut_LC_8_7_3 .C_ON=1'b1;
    defparam \tok.add_104_5_lut_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_5_lut_LC_8_7_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_5_lut_LC_8_7_3  (
            .in0(N__19594),
            .in1(N__29700),
            .in2(N__25373),
            .in3(N__19445),
            .lcout(\tok.n4_adj_806 ),
            .ltout(),
            .carryin(\tok.n4786 ),
            .carryout(\tok.n4787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_6_lut_LC_8_7_4 .C_ON=1'b1;
    defparam \tok.add_104_6_lut_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_6_lut_LC_8_7_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_6_lut_LC_8_7_4  (
            .in0(N__19593),
            .in1(N__29585),
            .in2(N__23762),
            .in3(N__19436),
            .lcout(\tok.n5564 ),
            .ltout(),
            .carryin(\tok.n4787 ),
            .carryout(\tok.n4788 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_7_lut_LC_8_7_5 .C_ON=1'b1;
    defparam \tok.add_104_7_lut_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_7_lut_LC_8_7_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_7_lut_LC_8_7_5  (
            .in0(N__19597),
            .in1(N__27303),
            .in2(N__27209),
            .in3(N__19433),
            .lcout(\tok.n5_adj_800 ),
            .ltout(),
            .carryin(\tok.n4788 ),
            .carryout(\tok.n4789 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_8_lut_LC_8_7_6 .C_ON=1'b1;
    defparam \tok.add_104_8_lut_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_8_lut_LC_8_7_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_8_lut_LC_8_7_6  (
            .in0(N__19592),
            .in1(N__21830),
            .in2(N__23666),
            .in3(N__19421),
            .lcout(\tok.n5554 ),
            .ltout(),
            .carryin(\tok.n4789 ),
            .carryout(\tok.n4790 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_9_lut_LC_8_7_7 .C_ON=1'b1;
    defparam \tok.add_104_9_lut_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_9_lut_LC_8_7_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_9_lut_LC_8_7_7  (
            .in0(N__19596),
            .in1(N__22258),
            .in2(N__23533),
            .in3(N__19406),
            .lcout(\tok.n5549 ),
            .ltout(),
            .carryin(\tok.n4790 ),
            .carryout(\tok.n4791 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_10_lut_LC_8_8_0 .C_ON=1'b1;
    defparam \tok.add_104_10_lut_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_10_lut_LC_8_8_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_10_lut_LC_8_8_0  (
            .in0(N__19590),
            .in1(N__29447),
            .in2(N__28066),
            .in3(N__19403),
            .lcout(\tok.n5_adj_669 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\tok.n4792 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_11_lut_LC_8_8_1 .C_ON=1'b1;
    defparam \tok.add_104_11_lut_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_11_lut_LC_8_8_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_11_lut_LC_8_8_1  (
            .in0(N__19601),
            .in1(N__29061),
            .in2(N__27531),
            .in3(N__19400),
            .lcout(\tok.n25 ),
            .ltout(),
            .carryin(\tok.n4792 ),
            .carryout(\tok.n4793 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_12_lut_LC_8_8_2 .C_ON=1'b1;
    defparam \tok.add_104_12_lut_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_12_lut_LC_8_8_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_12_lut_LC_8_8_2  (
            .in0(N__19587),
            .in1(N__29249),
            .in2(N__27459),
            .in3(N__19397),
            .lcout(\tok.n24_adj_703 ),
            .ltout(),
            .carryin(\tok.n4793 ),
            .carryout(\tok.n4794 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_13_lut_LC_8_8_3 .C_ON=1'b1;
    defparam \tok.add_104_13_lut_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_13_lut_LC_8_8_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_13_lut_LC_8_8_3  (
            .in0(N__19599),
            .in1(N__25146),
            .in2(N__25059),
            .in3(N__19394),
            .lcout(\tok.n5_adj_726 ),
            .ltout(),
            .carryin(\tok.n4794 ),
            .carryout(\tok.n4795 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_14_lut_LC_8_8_4 .C_ON=1'b1;
    defparam \tok.add_104_14_lut_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_14_lut_LC_8_8_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_14_lut_LC_8_8_4  (
            .in0(N__19586),
            .in1(N__21611),
            .in2(N__24477),
            .in3(N__19619),
            .lcout(\tok.n5_adj_734 ),
            .ltout(),
            .carryin(\tok.n4795 ),
            .carryout(\tok.n4796 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_15_lut_LC_8_8_5 .C_ON=1'b1;
    defparam \tok.add_104_15_lut_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_15_lut_LC_8_8_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_15_lut_LC_8_8_5  (
            .in0(N__19600),
            .in1(N__23150),
            .in2(N__24369),
            .in3(N__19616),
            .lcout(\tok.n5_adj_732 ),
            .ltout(),
            .carryin(\tok.n4796 ),
            .carryout(\tok.n4797 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_16_lut_LC_8_8_6 .C_ON=1'b1;
    defparam \tok.add_104_16_lut_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_16_lut_LC_8_8_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_16_lut_LC_8_8_6  (
            .in0(N__19589),
            .in1(N__28859),
            .in2(N__25772),
            .in3(N__19604),
            .lcout(\tok.n5_adj_716 ),
            .ltout(),
            .carryin(\tok.n4797 ),
            .carryout(\tok.n4798 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_17_lut_LC_8_8_7 .C_ON=1'b0;
    defparam \tok.add_104_17_lut_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_17_lut_LC_8_8_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \tok.add_104_17_lut_LC_8_8_7  (
            .in0(N__24860),
            .in1(N__19588),
            .in2(N__24778),
            .in3(N__19526),
            .lcout(\tok.n5_adj_713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5561_4_lut_LC_8_9_0 .C_ON=1'b0;
    defparam \tok.i5561_4_lut_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5561_4_lut_LC_8_9_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i5561_4_lut_LC_8_9_0  (
            .in0(N__22340),
            .in1(N__19523),
            .in2(N__20882),
            .in3(N__21011),
            .lcout(\tok.n5574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5242_4_lut_LC_8_9_1 .C_ON=1'b0;
    defparam \tok.i5242_4_lut_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5242_4_lut_LC_8_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \tok.i5242_4_lut_LC_8_9_1  (
            .in0(N__26940),
            .in1(N__21910),
            .in2(N__27878),
            .in3(N__19510),
            .lcout(),
            .ltout(\tok.n5414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_149_LC_8_9_2 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_149_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_149_LC_8_9_2 .LUT_INIT=16'b1111111101001111;
    LogicCell40 \tok.i6_4_lut_adj_149_LC_8_9_2  (
            .in0(N__22528),
            .in1(N__19499),
            .in2(N__19487),
            .in3(N__19484),
            .lcout(\tok.n904 ),
            .ltout(\tok.n904_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i47_3_lut_LC_8_9_3 .C_ON=1'b0;
    defparam \tok.i47_3_lut_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i47_3_lut_LC_8_9_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.i47_3_lut_LC_8_9_3  (
            .in0(N__27855),
            .in1(_gnd_net_),
            .in2(N__19478),
            .in3(N__22710),
            .lcout(),
            .ltout(\tok.n5346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_172_LC_8_9_4 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_172_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_172_LC_8_9_4 .LUT_INIT=16'b1101111111001111;
    LogicCell40 \tok.i6_4_lut_adj_172_LC_8_9_4  (
            .in0(N__22529),
            .in1(N__19475),
            .in2(N__19460),
            .in3(N__23225),
            .lcout(),
            .ltout(\tok.n14_adj_841_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5557_4_lut_LC_8_9_5 .C_ON=1'b0;
    defparam \tok.i5557_4_lut_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i5557_4_lut_LC_8_9_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.i5557_4_lut_LC_8_9_5  (
            .in0(N__19790),
            .in1(N__29750),
            .in2(N__19775),
            .in3(N__19772),
            .lcout(\tok.n5569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i49_3_lut_LC_8_9_6 .C_ON=1'b0;
    defparam \tok.i49_3_lut_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i49_3_lut_LC_8_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.i49_3_lut_LC_8_9_6  (
            .in0(N__29687),
            .in1(N__27854),
            .in2(_gnd_net_),
            .in3(N__27629),
            .lcout(\tok.n45_adj_849 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i3_1_lut_LC_8_9_7 .C_ON=1'b0;
    defparam \tok.inv_106_i3_1_lut_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i3_1_lut_LC_8_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i3_1_lut_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22709),
            .lcout(\tok.n300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_57_LC_8_10_0 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_57_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_57_LC_8_10_0 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \tok.i1_3_lut_adj_57_LC_8_10_0  (
            .in0(N__29345),
            .in1(N__21875),
            .in2(_gnd_net_),
            .in3(N__19745),
            .lcout(\tok.n45_adj_696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_50_LC_8_10_1 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_50_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_50_LC_8_10_1 .LUT_INIT=16'b1100110011101111;
    LogicCell40 \tok.i3_4_lut_adj_50_LC_8_10_1  (
            .in0(N__27325),
            .in1(N__19706),
            .in2(N__21314),
            .in3(N__26751),
            .lcout(\tok.n10_adj_686 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_LC_8_10_2 .C_ON=1'b0;
    defparam \tok.i1_3_lut_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_LC_8_10_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \tok.i1_3_lut_LC_8_10_2  (
            .in0(N__29344),
            .in1(N__27324),
            .in2(_gnd_net_),
            .in3(N__19744),
            .lcout(),
            .ltout(\tok.n45_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_46_LC_8_10_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_46_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_46_LC_8_10_3 .LUT_INIT=16'b0011000000110010;
    LogicCell40 \tok.i1_4_lut_adj_46_LC_8_10_3  (
            .in0(N__19724),
            .in1(N__19642),
            .in2(N__19709),
            .in3(N__19699),
            .lcout(\tok.n39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_58_LC_8_10_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_58_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_58_LC_8_10_4 .LUT_INIT=16'b0000111100000100;
    LogicCell40 \tok.i1_4_lut_adj_58_LC_8_10_4  (
            .in0(N__19700),
            .in1(N__19667),
            .in2(N__19646),
            .in3(N__19634),
            .lcout(),
            .ltout(\tok.n39_adj_697_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_60_LC_8_10_5 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_60_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_60_LC_8_10_5 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \tok.i3_4_lut_adj_60_LC_8_10_5  (
            .in0(N__21876),
            .in1(N__21311),
            .in2(N__19628),
            .in3(N__26752),
            .lcout(),
            .ltout(\tok.n10_adj_700_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5441_4_lut_LC_8_10_6 .C_ON=1'b0;
    defparam \tok.i5441_4_lut_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5441_4_lut_LC_8_10_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i5441_4_lut_LC_8_10_6  (
            .in0(N__27371),
            .in1(N__22616),
            .in2(N__19922),
            .in3(N__20852),
            .lcout(\tok.n5536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_180_LC_8_10_7 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_180_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_180_LC_8_10_7 .LUT_INIT=16'b0000101000111011;
    LogicCell40 \tok.i3_4_lut_adj_180_LC_8_10_7  (
            .in0(N__22882),
            .in1(N__20296),
            .in2(N__28789),
            .in3(N__28939),
            .lcout(\tok.n11_adj_730 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_66_LC_8_11_0 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_66_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_66_LC_8_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i10_4_lut_adj_66_LC_8_11_0  (
            .in0(N__27327),
            .in1(N__23111),
            .in2(N__29470),
            .in3(N__29701),
            .lcout(),
            .ltout(\tok.n26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i15_4_lut_LC_8_11_1 .C_ON=1'b0;
    defparam \tok.i15_4_lut_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i15_4_lut_LC_8_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i15_4_lut_LC_8_11_1  (
            .in0(N__19805),
            .in1(N__19796),
            .in2(N__19907),
            .in3(N__19811),
            .lcout(\tok.tc__7__N_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_LC_8_11_2 .C_ON=1'b0;
    defparam \tok.i9_4_lut_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_LC_8_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_LC_8_11_2  (
            .in0(N__27690),
            .in1(N__29552),
            .in2(N__21108),
            .in3(N__21865),
            .lcout(\tok.n25_adj_710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i12_4_lut_LC_8_11_3 .C_ON=1'b0;
    defparam \tok.i12_4_lut_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i12_4_lut_LC_8_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i12_4_lut_LC_8_11_3  (
            .in0(N__29038),
            .in1(N__25767),
            .in2(N__24844),
            .in3(N__25116),
            .lcout(\tok.n28_adj_708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i11_4_lut_LC_8_11_4 .C_ON=1'b0;
    defparam \tok.i11_4_lut_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i11_4_lut_LC_8_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i11_4_lut_LC_8_11_4  (
            .in0(N__22268),
            .in1(N__29215),
            .in2(N__22731),
            .in3(N__21595),
            .lcout(\tok.n27_adj_709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_94_LC_8_11_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_94_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_94_LC_8_11_5 .LUT_INIT=16'b0000110001011101;
    LogicCell40 \tok.i1_4_lut_adj_94_LC_8_11_5  (
            .in0(N__23112),
            .in1(N__29464),
            .in2(N__28979),
            .in3(N__27876),
            .lcout(\tok.n12_adj_745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_74_LC_8_11_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_74_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_74_LC_8_11_6 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \tok.i1_4_lut_adj_74_LC_8_11_6  (
            .in0(N__27874),
            .in1(N__28972),
            .in2(N__25145),
            .in3(N__21866),
            .lcout(\tok.n12_adj_723 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_116_LC_8_11_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_116_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_116_LC_8_11_7 .LUT_INIT=16'b0100010001001111;
    LogicCell40 \tok.i1_4_lut_adj_116_LC_8_11_7  (
            .in0(N__28973),
            .in1(N__29240),
            .in2(N__24845),
            .in3(N__27875),
            .lcout(\tok.n12_adj_779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_191_LC_8_12_0 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_191_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_191_LC_8_12_0 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \tok.i2_3_lut_adj_191_LC_8_12_0  (
            .in0(N__26747),
            .in1(N__20321),
            .in2(_gnd_net_),
            .in3(N__20272),
            .lcout(\tok.n10_adj_858 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_adj_97_LC_8_12_1 .C_ON=1'b0;
    defparam \tok.i5_3_lut_adj_97_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_adj_97_LC_8_12_1 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \tok.i5_3_lut_adj_97_LC_8_12_1  (
            .in0(N__26984),
            .in1(N__20003),
            .in2(_gnd_net_),
            .in3(N__19988),
            .lcout(\tok.n16_adj_749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_114_LC_8_12_2 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_114_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_114_LC_8_12_2 .LUT_INIT=16'b1101110111001101;
    LogicCell40 \tok.i3_4_lut_adj_114_LC_8_12_2  (
            .in0(N__26748),
            .in1(N__20342),
            .in2(N__21313),
            .in3(N__25167),
            .lcout(),
            .ltout(\tok.n14_adj_776_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_120_LC_8_12_3 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_120_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_120_LC_8_12_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_120_LC_8_12_3  (
            .in0(N__24071),
            .in1(N__19979),
            .in2(N__19973),
            .in3(N__19970),
            .lcout(),
            .ltout(\tok.n20_adj_784_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5572_4_lut_LC_8_12_4 .C_ON=1'b0;
    defparam \tok.i5572_4_lut_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5572_4_lut_LC_8_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i5572_4_lut_LC_8_12_4  (
            .in0(N__20699),
            .in1(N__19928),
            .in2(N__19964),
            .in3(N__19961),
            .lcout(\tok.n5513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_15_i9_2_lut_LC_8_12_5 .C_ON=1'b0;
    defparam \tok.select_73_Select_15_i9_2_lut_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_15_i9_2_lut_LC_8_12_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.select_73_Select_15_i9_2_lut_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__24767),
            .in2(_gnd_net_),
            .in3(N__28777),
            .lcout(\tok.n9_adj_781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_adj_118_LC_8_12_6 .C_ON=1'b0;
    defparam \tok.i5_3_lut_adj_118_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_adj_118_LC_8_12_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \tok.i5_3_lut_adj_118_LC_8_12_6  (
            .in0(N__19955),
            .in1(N__19946),
            .in2(_gnd_net_),
            .in3(N__26983),
            .lcout(\tok.n16_adj_782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_8_13_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_8_13_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_8_13_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_8_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_4_lut_adj_182_LC_8_13_2 .C_ON=1'b0;
    defparam \tok.i3_4_lut_4_lut_adj_182_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_4_lut_adj_182_LC_8_13_2 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i3_4_lut_4_lut_adj_182_LC_8_13_2  (
            .in0(N__28781),
            .in1(N__20357),
            .in2(N__23554),
            .in3(N__29139),
            .lcout(\tok.n14_adj_658 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_11_i2_3_lut_3_lut_LC_8_13_4 .C_ON=1'b0;
    defparam \tok.select_73_Select_11_i2_3_lut_3_lut_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_11_i2_3_lut_3_lut_LC_8_13_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \tok.select_73_Select_11_i2_3_lut_3_lut_LC_8_13_4  (
            .in0(N__29310),
            .in1(N__29138),
            .in2(_gnd_net_),
            .in3(N__22269),
            .lcout(\tok.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_15_i2_3_lut_3_lut_LC_8_14_6 .C_ON=1'b0;
    defparam \tok.select_73_Select_15_i2_3_lut_3_lut_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_15_i2_3_lut_3_lut_LC_8_14_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \tok.select_73_Select_15_i2_3_lut_3_lut_LC_8_14_6  (
            .in0(N__29319),
            .in1(N__29160),
            .in2(_gnd_net_),
            .in3(N__25166),
            .lcout(\tok.n2_adj_775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i102_LC_9_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i102_LC_9_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i102_LC_9_2_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i102_LC_9_2_3  (
            .in0(N__20333),
            .in1(N__20603),
            .in2(_gnd_net_),
            .in3(N__26526),
            .lcout(tail_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28500),
            .ce(N__26049),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i125_LC_9_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i125_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i125_LC_9_3_0 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i125_LC_9_3_0  (
            .in0(N__21443),
            .in1(N__26011),
            .in2(N__21460),
            .in3(N__26455),
            .lcout(tail_125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28507),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i123_LC_9_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i123_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i123_LC_9_3_1 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \tok.A_stk.tail_i0_i123_LC_9_3_1  (
            .in0(N__26453),
            .in1(N__21557),
            .in2(N__26055),
            .in3(N__21361),
            .lcout(tail_123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28507),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i124_LC_9_3_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i124_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i124_LC_9_3_2 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i124_LC_9_3_2  (
            .in0(N__21509),
            .in1(N__26010),
            .in2(N__21530),
            .in3(N__26454),
            .lcout(tail_124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28507),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i118_LC_9_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i118_LC_9_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i118_LC_9_3_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \tok.A_stk.tail_i0_i118_LC_9_3_3  (
            .in0(N__26451),
            .in1(N__20332),
            .in2(N__26054),
            .in3(N__20380),
            .lcout(tail_118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28507),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i122_LC_9_3_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i122_LC_9_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i122_LC_9_3_4 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i122_LC_9_3_4  (
            .in0(N__25211),
            .in1(N__26006),
            .in2(N__25228),
            .in3(N__26452),
            .lcout(tail_122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28507),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i116_LC_9_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i116_LC_9_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i116_LC_9_3_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \tok.A_stk.tail_i0_i116_LC_9_3_5  (
            .in0(N__26450),
            .in1(N__20468),
            .in2(N__26053),
            .in3(N__20449),
            .lcout(tail_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28507),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i114_LC_9_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i114_LC_9_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i114_LC_9_3_6 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i114_LC_9_3_6  (
            .in0(N__20419),
            .in1(N__25999),
            .in2(N__20437),
            .in3(N__26449),
            .lcout(tail_114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28507),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i23_LC_9_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i23_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i23_LC_9_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i23_LC_9_4_0  (
            .in0(N__20576),
            .in1(N__21745),
            .in2(_gnd_net_),
            .in3(N__26343),
            .lcout(\tok.A_stk.tail_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28512),
            .ce(N__26031),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i70_LC_9_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i70_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i70_LC_9_4_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i70_LC_9_4_1  (
            .in0(N__26347),
            .in1(N__20602),
            .in2(_gnd_net_),
            .in3(N__20524),
            .lcout(\tok.A_stk.tail_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28512),
            .ce(N__26031),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i98_LC_9_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i98_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i98_LC_9_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i98_LC_9_4_2  (
            .in0(N__20438),
            .in1(N__20401),
            .in2(_gnd_net_),
            .in3(N__26350),
            .lcout(tail_98),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28512),
            .ce(N__26031),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i66_LC_9_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i66_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i66_LC_9_4_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i66_LC_9_4_3  (
            .in0(N__26346),
            .in1(_gnd_net_),
            .in2(N__20405),
            .in3(N__21692),
            .lcout(\tok.A_stk.tail_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28512),
            .ce(N__26031),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i82_LC_9_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i82_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i82_LC_9_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i82_LC_9_4_4  (
            .in0(N__20420),
            .in1(N__21703),
            .in2(_gnd_net_),
            .in3(N__26348),
            .lcout(\tok.A_stk.tail_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28512),
            .ce(N__26031),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i56_LC_9_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i56_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i56_LC_9_4_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i56_LC_9_4_5  (
            .in0(N__26345),
            .in1(N__21977),
            .in2(_gnd_net_),
            .in3(N__20393),
            .lcout(\tok.A_stk.tail_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28512),
            .ce(N__26031),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i54_LC_9_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i54_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i54_LC_9_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i54_LC_9_4_6  (
            .in0(N__20366),
            .in1(N__20500),
            .in2(_gnd_net_),
            .in3(N__26344),
            .lcout(\tok.A_stk.tail_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28512),
            .ce(N__26031),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i86_LC_9_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i86_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i86_LC_9_4_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i86_LC_9_4_7  (
            .in0(N__26349),
            .in1(N__20381),
            .in2(_gnd_net_),
            .in3(N__20365),
            .lcout(\tok.A_stk.tail_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28512),
            .ce(N__26031),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i39_LC_9_5_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i39_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i39_LC_9_5_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i39_LC_9_5_0  (
            .in0(N__26508),
            .in1(N__20488),
            .in2(_gnd_net_),
            .in3(N__20588),
            .lcout(\tok.A_stk.tail_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28519),
            .ce(N__26021),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i67_LC_9_5_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i67_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i67_LC_9_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i67_LC_9_5_1  (
            .in0(N__26096),
            .in1(N__20564),
            .in2(_gnd_net_),
            .in3(N__26509),
            .lcout(\tok.A_stk.tail_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28519),
            .ce(N__26021),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i4_LC_9_5_2 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i4_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i4_LC_9_5_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i4_LC_9_5_2  (
            .in0(N__20549),
            .in1(N__25498),
            .in2(_gnd_net_),
            .in3(N__29599),
            .lcout(\tok.S_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28519),
            .ce(N__26021),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i6_LC_9_5_3 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i6_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i6_LC_9_5_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.head_i0_i6_LC_9_5_3  (
            .in0(N__25499),
            .in1(N__20536),
            .in2(_gnd_net_),
            .in3(N__21835),
            .lcout(\tok.S_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28519),
            .ce(N__26021),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i6_LC_9_5_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i6_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i6_LC_9_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i6_LC_9_5_4  (
            .in0(N__26510),
            .in1(N__20513),
            .in2(_gnd_net_),
            .in3(N__23648),
            .lcout(\tok.A_stk.tail_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28519),
            .ce(N__26021),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i22_LC_9_5_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i22_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i22_LC_9_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i22_LC_9_5_5  (
            .in0(N__20504),
            .in1(N__20537),
            .in2(_gnd_net_),
            .in3(N__26506),
            .lcout(\tok.A_stk.tail_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28519),
            .ce(N__26021),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i38_LC_9_5_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i38_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i38_LC_9_5_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i38_LC_9_5_6  (
            .in0(N__26507),
            .in1(_gnd_net_),
            .in2(N__20528),
            .in3(N__20512),
            .lcout(\tok.A_stk.tail_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28519),
            .ce(N__26021),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i7_LC_9_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i7_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i7_LC_9_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i7_LC_9_5_7  (
            .in0(N__23523),
            .in1(N__20489),
            .in2(_gnd_net_),
            .in3(N__26511),
            .lcout(\tok.A_stk.tail_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28519),
            .ce(N__26021),
            .sr(_gnd_net_));
    defparam \tok.add_109_2_lut_LC_9_6_0 .C_ON=1'b1;
    defparam \tok.add_109_2_lut_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_2_lut_LC_9_6_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_2_lut_LC_9_6_0  (
            .in0(N__20843),
            .in1(N__22881),
            .in2(_gnd_net_),
            .in3(N__20666),
            .lcout(\tok.n3_adj_692 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\tok.n4799 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_3_lut_LC_9_6_1 .C_ON=1'b1;
    defparam \tok.add_109_3_lut_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_3_lut_LC_9_6_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_3_lut_LC_9_6_1  (
            .in0(N__20839),
            .in1(N__24029),
            .in2(_gnd_net_),
            .in3(N__20663),
            .lcout(\tok.n14_adj_662 ),
            .ltout(),
            .carryin(\tok.n4799 ),
            .carryout(\tok.n4800 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_4_lut_LC_9_6_2 .C_ON=1'b1;
    defparam \tok.add_109_4_lut_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_4_lut_LC_9_6_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_4_lut_LC_9_6_2  (
            .in0(N__20842),
            .in1(N__23913),
            .in2(_gnd_net_),
            .in3(N__20660),
            .lcout(\tok.n12_adj_832 ),
            .ltout(),
            .carryin(\tok.n4800 ),
            .carryout(\tok.n4801 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_5_lut_LC_9_6_3 .C_ON=1'b1;
    defparam \tok.add_109_5_lut_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_5_lut_LC_9_6_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_5_lut_LC_9_6_3  (
            .in0(N__20838),
            .in1(N__25335),
            .in2(_gnd_net_),
            .in3(N__20645),
            .lcout(\tok.n22_adj_829 ),
            .ltout(),
            .carryin(\tok.n4801 ),
            .carryout(\tok.n4802 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_6_lut_LC_9_6_4 .C_ON=1'b1;
    defparam \tok.add_109_6_lut_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_6_lut_LC_9_6_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_6_lut_LC_9_6_4  (
            .in0(N__20765),
            .in1(N__23732),
            .in2(_gnd_net_),
            .in3(N__20630),
            .lcout(\tok.n10_adj_827 ),
            .ltout(),
            .carryin(\tok.n4802 ),
            .carryout(\tok.n4803 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_7_lut_LC_9_6_5 .C_ON=1'b1;
    defparam \tok.add_109_7_lut_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_7_lut_LC_9_6_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_7_lut_LC_9_6_5  (
            .in0(N__20767),
            .in1(N__27188),
            .in2(_gnd_net_),
            .in3(N__20627),
            .lcout(\tok.n10_adj_823 ),
            .ltout(),
            .carryin(\tok.n4803 ),
            .carryout(\tok.n4804 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_8_lut_LC_9_6_6 .C_ON=1'b1;
    defparam \tok.add_109_8_lut_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_8_lut_LC_9_6_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_8_lut_LC_9_6_6  (
            .in0(N__20766),
            .in1(N__23629),
            .in2(_gnd_net_),
            .in3(N__20618),
            .lcout(\tok.n10_adj_820 ),
            .ltout(),
            .carryin(\tok.n4804 ),
            .carryout(\tok.n4805 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_9_lut_LC_9_6_7 .C_ON=1'b1;
    defparam \tok.add_109_9_lut_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_9_lut_LC_9_6_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_9_lut_LC_9_6_7  (
            .in0(N__20768),
            .in1(N__23519),
            .in2(_gnd_net_),
            .in3(N__20609),
            .lcout(\tok.n10_adj_653 ),
            .ltout(),
            .carryin(\tok.n4805 ),
            .carryout(\tok.n4806 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_10_lut_LC_9_7_0 .C_ON=1'b1;
    defparam \tok.add_109_10_lut_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_10_lut_LC_9_7_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_10_lut_LC_9_7_0  (
            .in0(N__20750),
            .in1(N__28057),
            .in2(_gnd_net_),
            .in3(N__20606),
            .lcout(\tok.n10_adj_666 ),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\tok.n4807 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_11_lut_LC_9_7_1 .C_ON=1'b1;
    defparam \tok.add_109_11_lut_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_11_lut_LC_9_7_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_11_lut_LC_9_7_1  (
            .in0(N__20841),
            .in1(N__27539),
            .in2(_gnd_net_),
            .in3(N__20846),
            .lcout(\tok.n23_adj_682 ),
            .ltout(),
            .carryin(\tok.n4807 ),
            .carryout(\tok.n4808 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_12_lut_LC_9_7_2 .C_ON=1'b1;
    defparam \tok.add_109_12_lut_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_12_lut_LC_9_7_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_12_lut_LC_9_7_2  (
            .in0(N__20840),
            .in1(N__27441),
            .in2(_gnd_net_),
            .in3(N__20804),
            .lcout(\tok.n22_adj_698 ),
            .ltout(),
            .carryin(\tok.n4808 ),
            .carryout(\tok.n4809 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_13_lut_LC_9_7_3 .C_ON=1'b1;
    defparam \tok.add_109_13_lut_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_13_lut_LC_9_7_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_13_lut_LC_9_7_3  (
            .in0(N__20762),
            .in1(N__25054),
            .in2(_gnd_net_),
            .in3(N__20801),
            .lcout(\tok.n5534 ),
            .ltout(),
            .carryin(\tok.n4809 ),
            .carryout(\tok.n4810 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_14_lut_LC_9_7_4 .C_ON=1'b1;
    defparam \tok.add_109_14_lut_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_14_lut_LC_9_7_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_14_lut_LC_9_7_4  (
            .in0(N__20748),
            .in1(N__24464),
            .in2(_gnd_net_),
            .in3(N__20789),
            .lcout(\tok.n10_adj_738 ),
            .ltout(),
            .carryin(\tok.n4810 ),
            .carryout(\tok.n4811 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_15_lut_LC_9_7_5 .C_ON=1'b1;
    defparam \tok.add_109_15_lut_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_15_lut_LC_9_7_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_15_lut_LC_9_7_5  (
            .in0(N__20763),
            .in1(N__24365),
            .in2(_gnd_net_),
            .in3(N__20786),
            .lcout(\tok.n5525 ),
            .ltout(),
            .carryin(\tok.n4811 ),
            .carryout(\tok.n4812 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_16_lut_LC_9_7_6 .C_ON=1'b1;
    defparam \tok.add_109_16_lut_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_16_lut_LC_9_7_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_16_lut_LC_9_7_6  (
            .in0(N__20749),
            .in1(N__28866),
            .in2(_gnd_net_),
            .in3(N__20771),
            .lcout(\tok.n10_adj_768 ),
            .ltout(),
            .carryin(\tok.n4812 ),
            .carryout(\tok.n4813 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_17_lut_LC_9_7_7 .C_ON=1'b0;
    defparam \tok.add_109_17_lut_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_17_lut_LC_9_7_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \tok.add_109_17_lut_LC_9_7_7  (
            .in0(N__24777),
            .in1(N__20751),
            .in2(_gnd_net_),
            .in3(N__20702),
            .lcout(\tok.n5516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_90_LC_9_8_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_90_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_90_LC_9_8_0 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \tok.i1_4_lut_adj_90_LC_9_8_0  (
            .in0(N__21612),
            .in1(N__26760),
            .in2(N__20900),
            .in3(N__27624),
            .lcout(),
            .ltout(\tok.n12_adj_737_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_92_LC_9_8_1 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_92_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_92_LC_9_8_1 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \tok.i9_4_lut_adj_92_LC_9_8_1  (
            .in0(N__20684),
            .in1(N__22322),
            .in2(N__20669),
            .in3(N__28970),
            .lcout(\tok.n20_adj_740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_7_i1_4_lut_LC_9_8_3 .C_ON=1'b0;
    defparam \tok.select_73_Select_7_i1_4_lut_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_7_i1_4_lut_LC_9_8_3 .LUT_INIT=16'b0101010001000101;
    LogicCell40 \tok.select_73_Select_7_i1_4_lut_LC_9_8_3  (
            .in0(N__26761),
            .in1(N__29728),
            .in2(N__22187),
            .in3(N__22146),
            .lcout(),
            .ltout(\tok.n1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_36_LC_9_8_4 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_36_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_36_LC_9_8_4 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \tok.i6_4_lut_adj_36_LC_9_8_4  (
            .in0(N__23208),
            .in1(N__20915),
            .in2(N__20930),
            .in3(N__24843),
            .lcout(\tok.n17_adj_656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_7_i12_2_lut_3_lut_LC_9_8_5 .C_ON=1'b0;
    defparam \tok.select_73_Select_7_i12_2_lut_3_lut_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_7_i12_2_lut_3_lut_LC_9_8_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \tok.select_73_Select_7_i12_2_lut_3_lut_LC_9_8_5  (
            .in0(N__20908),
            .in1(N__22548),
            .in2(_gnd_net_),
            .in3(N__23332),
            .lcout(\tok.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i7_LC_9_8_6 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i7_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i7_LC_9_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i7_LC_9_8_6  (
            .in0(N__23008),
            .in1(N__25692),
            .in2(_gnd_net_),
            .in3(N__20909),
            .lcout(uart_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28533),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_99_i13_2_lut_3_lut_LC_9_8_7 .C_ON=1'b0;
    defparam \tok.or_99_i13_2_lut_3_lut_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i13_2_lut_3_lut_LC_9_8_7 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \tok.or_99_i13_2_lut_3_lut_LC_9_8_7  (
            .in0(N__22182),
            .in1(N__29448),
            .in2(_gnd_net_),
            .in3(N__22145),
            .lcout(\tok.n177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_168_LC_9_9_0 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_168_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_168_LC_9_9_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \tok.i2_3_lut_adj_168_LC_9_9_0  (
            .in0(N__20891),
            .in1(N__28758),
            .in2(_gnd_net_),
            .in3(N__24039),
            .lcout(\tok.n9_adj_838 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_47_LC_9_9_1 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_47_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_47_LC_9_9_1 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \tok.i1_3_lut_adj_47_LC_9_9_1  (
            .in0(N__20873),
            .in1(N__21135),
            .in2(_gnd_net_),
            .in3(N__23336),
            .lcout(),
            .ltout(\tok.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_53_LC_9_9_2 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_53_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_53_LC_9_9_2 .LUT_INIT=16'b1010101011111110;
    LogicCell40 \tok.i2_4_lut_adj_53_LC_9_9_2  (
            .in0(N__20861),
            .in1(N__24608),
            .in2(N__20855),
            .in3(N__22549),
            .lcout(\tok.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i59_3_lut_adj_63_LC_9_9_3 .C_ON=1'b0;
    defparam \tok.i59_3_lut_adj_63_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i59_3_lut_adj_63_LC_9_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.i59_3_lut_adj_63_LC_9_9_3  (
            .in0(N__29270),
            .in1(N__27857),
            .in2(_gnd_net_),
            .in3(N__27631),
            .lcout(\tok.n5350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i1_LC_9_9_4 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i1_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i1_LC_9_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i1_LC_9_9_4  (
            .in0(N__21188),
            .in1(N__25694),
            .in2(_gnd_net_),
            .in3(N__22600),
            .lcout(uart_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28538),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i59_3_lut_LC_9_9_5 .C_ON=1'b0;
    defparam \tok.i59_3_lut_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i59_3_lut_LC_9_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.i59_3_lut_LC_9_9_5  (
            .in0(N__29079),
            .in1(N__27858),
            .in2(_gnd_net_),
            .in3(N__27632),
            .lcout(),
            .ltout(\tok.n5342_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5560_4_lut_LC_9_9_6 .C_ON=1'b0;
    defparam \tok.i5560_4_lut_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5560_4_lut_LC_9_9_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.i5560_4_lut_LC_9_9_6  (
            .in0(N__27476),
            .in1(N__21158),
            .in2(N__21152),
            .in3(N__21149),
            .lcout(\tok.n5539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i44_3_lut_LC_9_9_7 .C_ON=1'b0;
    defparam \tok.i44_3_lut_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i44_3_lut_LC_9_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.i44_3_lut_LC_9_9_7  (
            .in0(N__21136),
            .in1(N__27856),
            .in2(_gnd_net_),
            .in3(N__27630),
            .lcout(\tok.n5336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_11_i9_2_lut_LC_9_10_0 .C_ON=1'b0;
    defparam \tok.select_73_Select_11_i9_2_lut_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_11_i9_2_lut_LC_9_10_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \tok.select_73_Select_11_i9_2_lut_LC_9_10_0  (
            .in0(N__28782),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25055),
            .lcout(\tok.n9_adj_725 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_adj_76_LC_9_10_1 .C_ON=1'b0;
    defparam \tok.i5_3_lut_adj_76_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_adj_76_LC_9_10_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i5_3_lut_adj_76_LC_9_10_1  (
            .in0(N__21005),
            .in1(N__20987),
            .in2(_gnd_net_),
            .in3(N__26993),
            .lcout(\tok.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_75_LC_9_10_2 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_75_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_75_LC_9_10_2 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \tok.i2_4_lut_adj_75_LC_9_10_2  (
            .in0(N__25157),
            .in1(N__29704),
            .in2(N__27953),
            .in3(N__27625),
            .lcout(),
            .ltout(\tok.n13_adj_724_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_78_LC_9_10_3 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_78_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_78_LC_9_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_78_LC_9_10_3  (
            .in0(N__24509),
            .in1(N__21230),
            .in2(N__20975),
            .in3(N__20972),
            .lcout(),
            .ltout(\tok.n20_adj_729_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5567_4_lut_LC_9_10_4 .C_ON=1'b0;
    defparam \tok.i5567_4_lut_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5567_4_lut_LC_9_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i5567_4_lut_LC_9_10_4  (
            .in0(N__20966),
            .in1(N__20957),
            .in2(N__20951),
            .in3(N__20948),
            .lcout(\tok.n5531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_73_LC_9_10_5 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_73_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_73_LC_9_10_5 .LUT_INIT=16'b1010101011101111;
    LogicCell40 \tok.i3_4_lut_adj_73_LC_9_10_5  (
            .in0(N__21239),
            .in1(N__22299),
            .in2(N__21312),
            .in3(N__26749),
            .lcout(\tok.n14_adj_722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i11_1_lut_LC_9_10_6 .C_ON=1'b0;
    defparam \tok.inv_106_i11_1_lut_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i11_1_lut_LC_9_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i11_1_lut_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29253),
            .lcout(\tok.n292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i12_1_lut_LC_9_10_7 .C_ON=1'b0;
    defparam \tok.inv_106_i12_1_lut_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i12_1_lut_LC_9_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i12_1_lut_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25156),
            .lcout(\tok.n291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5583_4_lut_LC_9_11_0 .C_ON=1'b0;
    defparam \tok.i5583_4_lut_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5583_4_lut_LC_9_11_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.i5583_4_lut_LC_9_11_0  (
            .in0(N__24404),
            .in1(N__21248),
            .in2(N__21197),
            .in3(N__21224),
            .lcout(),
            .ltout(\tok.n5527_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i13_LC_9_11_1 .C_ON=1'b0;
    defparam \tok.A_i13_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \tok.A_i13_LC_9_11_1 .LUT_INIT=16'b1110010011101110;
    LogicCell40 \tok.A_i13_LC_9_11_1  (
            .in0(N__28652),
            .in1(N__24480),
            .in2(N__21215),
            .in3(N__26855),
            .lcout(\tok.A_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28542),
            .ce(N__28296),
            .sr(N__28230));
    defparam \tok.A_i14_LC_9_11_2 .C_ON=1'b0;
    defparam \tok.A_i14_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \tok.A_i14_LC_9_11_2 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \tok.A_i14_LC_9_11_2  (
            .in0(N__26856),
            .in1(N__28653),
            .in2(N__24374),
            .in3(N__21320),
            .lcout(\tok.A_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28542),
            .ce(N__28296),
            .sr(N__28230));
    defparam \tok.A_i16_LC_9_11_3 .C_ON=1'b0;
    defparam \tok.A_i16_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \tok.A_i16_LC_9_11_3 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \tok.A_i16_LC_9_11_3  (
            .in0(N__24746),
            .in1(N__26857),
            .in2(N__28658),
            .in3(N__21212),
            .lcout(\tok.A_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28542),
            .ce(N__28296),
            .sr(N__28230));
    defparam \tok.A_i10_LC_9_11_5 .C_ON=1'b0;
    defparam \tok.A_i10_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \tok.A_i10_LC_9_11_5 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \tok.A_i10_LC_9_11_5  (
            .in0(N__27550),
            .in1(N__26854),
            .in2(N__28657),
            .in3(N__21206),
            .lcout(\tok.A_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28542),
            .ce(N__28296),
            .sr(N__28230));
    defparam \tok.i5181_2_lut_LC_9_11_6 .C_ON=1'b0;
    defparam \tok.i5181_2_lut_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5181_2_lut_LC_9_11_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i5181_2_lut_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__27877),
            .in2(_gnd_net_),
            .in3(N__21599),
            .lcout(\tok.n5348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_4_lut_LC_9_11_7 .C_ON=1'b0;
    defparam \tok.i8_4_lut_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i8_4_lut_LC_9_11_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i8_4_lut_LC_9_11_7  (
            .in0(N__27549),
            .in1(N__24825),
            .in2(N__24760),
            .in3(N__29039),
            .lcout(\tok.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_95_LC_9_12_0 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_95_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_95_LC_9_12_0 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \tok.i2_4_lut_adj_95_LC_9_12_0  (
            .in0(N__27343),
            .in1(N__23116),
            .in2(N__27959),
            .in3(N__27650),
            .lcout(),
            .ltout(\tok.n13_adj_746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_99_LC_9_12_1 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_99_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_99_LC_9_12_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_99_LC_9_12_1  (
            .in0(N__24278),
            .in1(N__21269),
            .in2(N__21350),
            .in3(N__21347),
            .lcout(),
            .ltout(\tok.n20_adj_753_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5581_4_lut_LC_9_12_2 .C_ON=1'b0;
    defparam \tok.i5581_4_lut_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5581_4_lut_LC_9_12_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i5581_4_lut_LC_9_12_2  (
            .in0(N__21341),
            .in1(N__21329),
            .in2(N__21323),
            .in3(N__21263),
            .lcout(\tok.n5522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_93_LC_9_12_3 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_93_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_93_LC_9_12_3 .LUT_INIT=16'b1010101011111011;
    LogicCell40 \tok.i3_4_lut_adj_93_LC_9_12_3  (
            .in0(N__21257),
            .in1(N__21304),
            .in2(N__29065),
            .in3(N__26750),
            .lcout(\tok.n14_adj_744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_13_i9_2_lut_LC_9_12_5 .C_ON=1'b0;
    defparam \tok.select_73_Select_13_i9_2_lut_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_13_i9_2_lut_LC_9_12_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.select_73_Select_13_i9_2_lut_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__24370),
            .in2(_gnd_net_),
            .in3(N__28783),
            .lcout(\tok.n9_adj_748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_13_i2_3_lut_3_lut_LC_9_12_7 .C_ON=1'b0;
    defparam \tok.select_73_Select_13_i2_3_lut_3_lut_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_13_i2_3_lut_3_lut_LC_9_12_7 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \tok.select_73_Select_13_i2_3_lut_3_lut_LC_9_12_7  (
            .in0(N__29343),
            .in1(N__29153),
            .in2(_gnd_net_),
            .in3(N__29040),
            .lcout(\tok.n2_adj_743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_101_i13_2_lut_LC_9_13_3 .C_ON=1'b0;
    defparam \tok.or_101_i13_2_lut_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.or_101_i13_2_lut_LC_9_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.or_101_i13_2_lut_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__29349),
            .in2(_gnd_net_),
            .in3(N__29460),
            .lcout(),
            .ltout(\tok.n204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_4_lut_LC_9_13_4 .C_ON=1'b0;
    defparam \tok.i5_4_lut_4_lut_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_4_lut_LC_9_13_4 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i5_4_lut_4_lut_LC_9_13_4  (
            .in0(N__29171),
            .in1(N__24479),
            .in2(N__21251),
            .in3(N__28790),
            .lcout(\tok.n16_adj_741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i109_LC_11_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i109_LC_11_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i109_LC_11_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i109_LC_11_2_0  (
            .in0(N__21467),
            .in1(N__21424),
            .in2(_gnd_net_),
            .in3(N__26574),
            .lcout(tail_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28508),
            .ce(N__26073),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i93_LC_11_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i93_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i93_LC_11_2_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i93_LC_11_2_1  (
            .in0(N__26580),
            .in1(N__21436),
            .in2(_gnd_net_),
            .in3(N__21412),
            .lcout(\tok.A_stk.tail_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28508),
            .ce(N__26073),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i77_LC_11_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i77_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i77_LC_11_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i77_LC_11_2_2  (
            .in0(N__21425),
            .in1(N__21403),
            .in2(_gnd_net_),
            .in3(N__26579),
            .lcout(\tok.A_stk.tail_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28508),
            .ce(N__26073),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i61_LC_11_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i61_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i61_LC_11_2_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i61_LC_11_2_3  (
            .in0(N__26578),
            .in1(N__21394),
            .in2(_gnd_net_),
            .in3(N__21413),
            .lcout(\tok.A_stk.tail_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28508),
            .ce(N__26073),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i45_LC_11_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i45_LC_11_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i45_LC_11_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i45_LC_11_2_4  (
            .in0(N__21385),
            .in1(N__21404),
            .in2(_gnd_net_),
            .in3(N__26577),
            .lcout(\tok.A_stk.tail_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28508),
            .ce(N__26073),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i29_LC_11_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i29_LC_11_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i29_LC_11_2_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.A_stk.tail_i0_i29_LC_11_2_5  (
            .in0(N__26576),
            .in1(_gnd_net_),
            .in2(N__21377),
            .in3(N__21395),
            .lcout(\tok.A_stk.tail_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28508),
            .ce(N__26073),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i13_LC_11_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i13_LC_11_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i13_LC_11_2_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i13_LC_11_2_6  (
            .in0(N__21386),
            .in1(N__26575),
            .in2(_gnd_net_),
            .in3(N__24319),
            .lcout(\tok.A_stk.tail_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28508),
            .ce(N__26073),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i13_LC_11_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i13_LC_11_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i13_LC_11_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i13_LC_11_2_7  (
            .in0(N__21373),
            .in1(N__25512),
            .in2(_gnd_net_),
            .in3(N__23162),
            .lcout(\tok.S_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28508),
            .ce(N__26073),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i107_LC_11_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i107_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i107_LC_11_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i107_LC_11_3_0  (
            .in0(N__21365),
            .in1(N__21541),
            .in2(_gnd_net_),
            .in3(N__26560),
            .lcout(tail_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28513),
            .ce(N__26058),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i91_LC_11_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i91_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i91_LC_11_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i91_LC_11_3_1  (
            .in0(N__26566),
            .in1(N__21553),
            .in2(_gnd_net_),
            .in3(N__25564),
            .lcout(\tok.A_stk.tail_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28513),
            .ce(N__26058),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i75_LC_11_3_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i75_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i75_LC_11_3_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i75_LC_11_3_2  (
            .in0(N__21542),
            .in1(N__25553),
            .in2(_gnd_net_),
            .in3(N__26564),
            .lcout(\tok.A_stk.tail_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28513),
            .ce(N__26058),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i108_LC_11_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i108_LC_11_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i108_LC_11_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i108_LC_11_3_3  (
            .in0(N__26561),
            .in1(N__21529),
            .in2(_gnd_net_),
            .in3(N__21493),
            .lcout(tail_108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28513),
            .ce(N__26058),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i92_LC_11_3_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i92_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i92_LC_11_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i92_LC_11_3_4  (
            .in0(N__21505),
            .in1(N__21484),
            .in2(_gnd_net_),
            .in3(N__26567),
            .lcout(\tok.A_stk.tail_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28513),
            .ce(N__26058),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i76_LC_11_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i76_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i76_LC_11_3_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i76_LC_11_3_5  (
            .in0(N__26565),
            .in1(N__21494),
            .in2(_gnd_net_),
            .in3(N__21475),
            .lcout(\tok.A_stk.tail_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28513),
            .ce(N__26058),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i60_LC_11_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i60_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i60_LC_11_3_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i60_LC_11_3_6  (
            .in0(N__21673),
            .in1(N__21485),
            .in2(_gnd_net_),
            .in3(N__26563),
            .lcout(\tok.A_stk.tail_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28513),
            .ce(N__26058),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i44_LC_11_3_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i44_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i44_LC_11_3_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i44_LC_11_3_7  (
            .in0(N__26562),
            .in1(N__21662),
            .in2(_gnd_net_),
            .in3(N__21476),
            .lcout(\tok.A_stk.tail_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28513),
            .ce(N__26058),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_LC_11_4_0 .C_ON=1'b0;
    defparam \tok.i6_4_lut_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_LC_11_4_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i6_4_lut_LC_11_4_0  (
            .in0(N__23880),
            .in1(N__22311),
            .in2(N__23507),
            .in3(N__22762),
            .lcout(\tok.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i2_LC_11_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i2_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i2_LC_11_4_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i2_LC_11_4_2  (
            .in0(N__21733),
            .in1(N__25450),
            .in2(_gnd_net_),
            .in3(N__22763),
            .lcout(\tok.S_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28520),
            .ce(N__26035),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i7_LC_11_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i7_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i7_LC_11_4_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.head_i0_i7_LC_11_4_3  (
            .in0(N__22312),
            .in1(N__21752),
            .in2(_gnd_net_),
            .in3(N__25451),
            .lcout(\tok.S_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28520),
            .ce(N__26035),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i2_LC_11_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i2_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i2_LC_11_4_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \tok.A_stk.tail_i0_i2_LC_11_4_4  (
            .in0(N__23881),
            .in1(_gnd_net_),
            .in2(N__26582),
            .in3(N__21725),
            .lcout(\tok.A_stk.tail_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28520),
            .ce(N__26035),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i18_LC_11_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i18_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i18_LC_11_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i18_LC_11_4_5  (
            .in0(N__21716),
            .in1(N__21734),
            .in2(_gnd_net_),
            .in3(N__26512),
            .lcout(\tok.A_stk.tail_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28520),
            .ce(N__26035),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i34_LC_11_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i34_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i34_LC_11_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i34_LC_11_4_6  (
            .in0(N__26516),
            .in1(N__21724),
            .in2(_gnd_net_),
            .in3(N__21691),
            .lcout(\tok.A_stk.tail_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28520),
            .ce(N__26035),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i50_LC_11_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i50_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i50_LC_11_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i50_LC_11_4_7  (
            .in0(N__21715),
            .in1(N__21707),
            .in2(_gnd_net_),
            .in3(N__26517),
            .lcout(\tok.A_stk.tail_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28520),
            .ce(N__26035),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i12_LC_11_5_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i12_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i12_LC_11_5_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i12_LC_11_5_0  (
            .in0(N__21661),
            .in1(N__26527),
            .in2(_gnd_net_),
            .in3(N__24457),
            .lcout(\tok.A_stk.tail_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28525),
            .ce(N__26059),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i28_LC_11_5_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i28_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i28_LC_11_5_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.A_stk.tail_i0_i28_LC_11_5_1  (
            .in0(N__26529),
            .in1(_gnd_net_),
            .in2(N__21647),
            .in3(N__21677),
            .lcout(\tok.A_stk.tail_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28525),
            .ce(N__26059),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i12_LC_11_5_2 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i12_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i12_LC_11_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.head_i0_i12_LC_11_5_2  (
            .in0(N__21635),
            .in1(N__21643),
            .in2(_gnd_net_),
            .in3(N__25500),
            .lcout(\tok.S_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28525),
            .ce(N__26059),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i13_1_lut_LC_11_5_3 .C_ON=1'b0;
    defparam \tok.inv_106_i13_1_lut_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i13_1_lut_LC_11_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i13_1_lut_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21634),
            .lcout(\tok.n290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i8_LC_11_5_4 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i8_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i8_LC_11_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.head_i0_i8_LC_11_5_4  (
            .in0(N__29452),
            .in1(N__22018),
            .in2(_gnd_net_),
            .in3(N__25501),
            .lcout(\tok.S_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28525),
            .ce(N__26059),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i8_LC_11_5_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i8_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i8_LC_11_5_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i8_LC_11_5_5  (
            .in0(N__26531),
            .in1(_gnd_net_),
            .in2(N__22010),
            .in3(N__28035),
            .lcout(\tok.A_stk.tail_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28525),
            .ce(N__26059),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i24_LC_11_5_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i24_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i24_LC_11_5_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i24_LC_11_5_6  (
            .in0(N__21973),
            .in1(N__22019),
            .in2(_gnd_net_),
            .in3(N__26528),
            .lcout(\tok.A_stk.tail_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28525),
            .ce(N__26059),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i40_LC_11_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i40_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i40_LC_11_5_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.A_stk.tail_i0_i40_LC_11_5_7  (
            .in0(N__26530),
            .in1(_gnd_net_),
            .in2(N__22009),
            .in3(N__21995),
            .lcout(\tok.A_stk.tail_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28525),
            .ce(N__26059),
            .sr(_gnd_net_));
    defparam \tok.i14_4_lut_LC_11_6_0 .C_ON=1'b0;
    defparam \tok.i14_4_lut_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i14_4_lut_LC_11_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i14_4_lut_LC_11_6_0  (
            .in0(N__21959),
            .in1(N__25190),
            .in2(N__21950),
            .in3(N__21932),
            .lcout(),
            .ltout(\tok.n30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5151_3_lut_LC_11_6_1 .C_ON=1'b0;
    defparam \tok.i5151_3_lut_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5151_3_lut_LC_11_6_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \tok.i5151_3_lut_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__21758),
            .in2(N__21917),
            .in3(N__21914),
            .lcout(\tok.n4908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_LC_11_6_2 .C_ON=1'b0;
    defparam \tok.i3_4_lut_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_LC_11_6_2 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \tok.i3_4_lut_LC_11_6_2  (
            .in0(N__28028),
            .in1(N__29459),
            .in2(N__24341),
            .in3(N__23158),
            .lcout(\tok.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_38_LC_11_6_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_38_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_38_LC_11_6_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i1_4_lut_adj_38_LC_11_6_3  (
            .in0(N__22872),
            .in1(N__21864),
            .in2(N__23677),
            .in3(N__27774),
            .lcout(),
            .ltout(\tok.n17_adj_661_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i13_4_lut_LC_11_6_4 .C_ON=1'b0;
    defparam \tok.i13_4_lut_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i13_4_lut_LC_11_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i13_4_lut_LC_11_6_4  (
            .in0(N__25535),
            .in1(N__21782),
            .in2(N__21767),
            .in3(N__21764),
            .lcout(\tok.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_163_LC_11_7_0 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_163_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_163_LC_11_7_0 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \tok.i2_3_lut_adj_163_LC_11_7_0  (
            .in0(N__23951),
            .in1(N__29075),
            .in2(_gnd_net_),
            .in3(N__23406),
            .lcout(\tok.n6_adj_834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_59_LC_11_7_1 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_59_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_59_LC_11_7_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i1_3_lut_adj_59_LC_11_7_1  (
            .in0(N__22764),
            .in1(N__22646),
            .in2(_gnd_net_),
            .in3(N__23331),
            .lcout(),
            .ltout(\tok.n4_adj_699_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_62_LC_11_7_2 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_62_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_62_LC_11_7_2 .LUT_INIT=16'b1100110011111110;
    LogicCell40 \tok.i2_4_lut_adj_62_LC_11_7_2  (
            .in0(N__24536),
            .in1(N__22634),
            .in2(N__22619),
            .in3(N__22544),
            .lcout(\tok.n9_adj_705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_164_LC_11_7_3 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_164_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_164_LC_11_7_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i1_3_lut_adj_164_LC_11_7_3  (
            .in0(N__22604),
            .in1(N__22586),
            .in2(_gnd_net_),
            .in3(N__23330),
            .lcout(),
            .ltout(\tok.n5_adj_835_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_165_LC_11_7_4 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_165_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_165_LC_11_7_4 .LUT_INIT=16'b1100110011111110;
    LogicCell40 \tok.i3_4_lut_adj_165_LC_11_7_4  (
            .in0(N__22574),
            .in1(N__22568),
            .in2(N__22553),
            .in3(N__22543),
            .lcout(\tok.n10_adj_836 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i8_1_lut_LC_11_7_5 .C_ON=1'b0;
    defparam \tok.inv_106_i8_1_lut_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i8_1_lut_LC_11_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i8_1_lut_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22310),
            .lcout(\tok.n295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i10_1_lut_LC_11_7_6 .C_ON=1'b0;
    defparam \tok.inv_106_i10_1_lut_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i10_1_lut_LC_11_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i10_1_lut_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29074),
            .lcout(\tok.n293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_99_i15_2_lut_3_lut_LC_11_7_7 .C_ON=1'b0;
    defparam \tok.or_99_i15_2_lut_3_lut_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i15_2_lut_3_lut_LC_11_7_7 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \tok.or_99_i15_2_lut_3_lut_LC_11_7_7  (
            .in0(N__29269),
            .in1(N__22186),
            .in2(_gnd_net_),
            .in3(N__22151),
            .lcout(\tok.n175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_inv_0_i1_1_lut_LC_11_8_0 .C_ON=1'b0;
    defparam \tok.sub_105_inv_0_i1_1_lut_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_inv_0_i1_1_lut_LC_11_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.sub_105_inv_0_i1_1_lut_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27766),
            .lcout(\tok.n17_adj_711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_169_LC_11_8_1 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_169_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_169_LC_11_8_1 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \tok.i2_3_lut_adj_169_LC_11_8_1  (
            .in0(N__23825),
            .in1(N__29271),
            .in2(_gnd_net_),
            .in3(N__23411),
            .lcout(),
            .ltout(\tok.n6_adj_839_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_170_LC_11_8_2 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_170_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_170_LC_11_8_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i3_4_lut_adj_170_LC_11_8_2  (
            .in0(N__23366),
            .in1(N__23351),
            .in2(N__23339),
            .in3(N__23333),
            .lcout(\tok.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5550_2_lut_LC_11_8_3 .C_ON=1'b0;
    defparam \tok.i5550_2_lut_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5550_2_lut_LC_11_8_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \tok.i5550_2_lut_LC_11_8_3  (
            .in0(N__23204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23155),
            .lcout(\tok.n5559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_4_lut_LC_11_8_4 .C_ON=1'b0;
    defparam \tok.i4_4_lut_4_lut_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_4_lut_LC_11_8_4 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \tok.i4_4_lut_4_lut_LC_11_8_4  (
            .in0(N__23069),
            .in1(N__29178),
            .in2(N__23054),
            .in3(N__26765),
            .lcout(\tok.n16_adj_855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i6_LC_11_8_5 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i6_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i6_LC_11_8_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.uart.capture_i0_i6_LC_11_8_5  (
            .in0(N__22906),
            .in1(_gnd_net_),
            .in2(N__25615),
            .in3(N__22971),
            .lcout(capture_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28539),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i5_LC_11_8_6 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i5_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i5_LC_11_8_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.uart.capture_i0_i5_LC_11_8_6  (
            .in0(N__22970),
            .in1(N__23023),
            .in2(_gnd_net_),
            .in3(N__25611),
            .lcout(capture_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28539),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i7_LC_11_8_7 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i7_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i7_LC_11_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.uart.capture_i0_i7_LC_11_8_7  (
            .in0(N__22905),
            .in1(N__23012),
            .in2(_gnd_net_),
            .in3(N__22972),
            .lcout(capture_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28539),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_2_lut_LC_11_9_0 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_2_lut_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_2_lut_LC_11_9_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_2_lut_LC_11_9_0  (
            .in0(N__24592),
            .in1(N__22892),
            .in2(N__22871),
            .in3(N__22769),
            .lcout(\tok.n11_adj_809 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\tok.n4769 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_3_lut_LC_11_9_1 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_3_lut_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_3_lut_LC_11_9_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_3_lut_LC_11_9_1  (
            .in0(N__24588),
            .in1(N__24059),
            .in2(N__24043),
            .in3(N__23942),
            .lcout(\tok.n20_adj_799 ),
            .ltout(),
            .carryin(\tok.n4769 ),
            .carryout(\tok.n4770 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_4_lut_LC_11_9_2 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_4_lut_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_4_lut_LC_11_9_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_4_lut_LC_11_9_2  (
            .in0(N__24591),
            .in1(N__23906),
            .in2(N__23840),
            .in3(N__23816),
            .lcout(\tok.n22_adj_797 ),
            .ltout(),
            .carryin(\tok.n4770 ),
            .carryout(\tok.n4771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_5_lut_LC_11_9_3 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_5_lut_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_5_lut_LC_11_9_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_5_lut_LC_11_9_3  (
            .in0(N__24589),
            .in1(N__25339),
            .in2(N__25529),
            .in3(N__23798),
            .lcout(\tok.n10_adj_791 ),
            .ltout(),
            .carryin(\tok.n4771 ),
            .carryout(\tok.n4772 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_6_lut_LC_11_9_4 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_6_lut_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_6_lut_LC_11_9_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_6_lut_LC_11_9_4  (
            .in0(N__24141),
            .in1(N__23775),
            .in2(N__27362),
            .in3(N__23684),
            .lcout(\tok.n6_adj_762 ),
            .ltout(),
            .carryin(\tok.n4772 ),
            .carryout(\tok.n4773 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_7_lut_LC_11_9_5 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_7_lut_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_7_lut_LC_11_9_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_7_lut_LC_11_9_5  (
            .in0(N__24135),
            .in1(N__27227),
            .in2(N__27214),
            .in3(N__23681),
            .lcout(\tok.n6_adj_717 ),
            .ltout(),
            .carryin(\tok.n4773 ),
            .carryout(\tok.n4774 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_8_lut_LC_11_9_6 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_8_lut_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_8_lut_LC_11_9_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_8_lut_LC_11_9_6  (
            .in0(N__24142),
            .in1(N__23664),
            .in2(N__23588),
            .in3(N__23561),
            .lcout(\tok.n6 ),
            .ltout(),
            .carryin(\tok.n4774 ),
            .carryout(\tok.n4775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_9_lut_LC_11_9_7 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_9_lut_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_9_lut_LC_11_9_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_9_lut_LC_11_9_7  (
            .in0(N__24134),
            .in1(N__23506),
            .in2(N__23444),
            .in3(N__23417),
            .lcout(\tok.n6_adj_657 ),
            .ltout(),
            .carryin(\tok.n4775 ),
            .carryout(\tok.n4776 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_10_lut_LC_11_10_0 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_10_lut_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_10_lut_LC_11_10_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_10_lut_LC_11_10_0  (
            .in0(N__24139),
            .in1(N__29360),
            .in2(N__28067),
            .in3(N__23414),
            .lcout(\tok.n5544 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\tok.n4777 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_11_lut_LC_11_10_1 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_11_lut_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_11_lut_LC_11_10_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_11_lut_LC_11_10_1  (
            .in0(N__24590),
            .in1(N__27545),
            .in2(N__24620),
            .in3(N__24596),
            .lcout(\tok.n28 ),
            .ltout(),
            .carryin(\tok.n4777 ),
            .carryout(\tok.n4778 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_12_lut_LC_11_10_2 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_12_lut_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_12_lut_LC_11_10_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_12_lut_LC_11_10_2  (
            .in0(N__24593),
            .in1(N__27440),
            .in2(N__24548),
            .in3(N__24527),
            .lcout(\tok.n27_adj_704 ),
            .ltout(),
            .carryin(\tok.n4778 ),
            .carryout(\tok.n4779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_13_lut_LC_11_10_3 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_13_lut_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_13_lut_LC_11_10_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_13_lut_LC_11_10_3  (
            .in0(N__24136),
            .in1(N__25041),
            .in2(N__24524),
            .in3(N__24500),
            .lcout(\tok.n6_adj_728 ),
            .ltout(),
            .carryin(\tok.n4779 ),
            .carryout(\tok.n4780 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_14_lut_LC_11_10_4 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_14_lut_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_14_lut_LC_11_10_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_14_lut_LC_11_10_4  (
            .in0(N__24140),
            .in1(N__24497),
            .in2(N__24478),
            .in3(N__24392),
            .lcout(\tok.n6_adj_742 ),
            .ltout(),
            .carryin(\tok.n4780 ),
            .carryout(\tok.n4781 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_15_lut_LC_11_10_5 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_15_lut_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_15_lut_LC_11_10_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_15_lut_LC_11_10_5  (
            .in0(N__24137),
            .in1(N__24389),
            .in2(N__24364),
            .in3(N__24266),
            .lcout(\tok.n6_adj_752 ),
            .ltout(),
            .carryin(\tok.n4781 ),
            .carryout(\tok.n4782 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_16_lut_LC_11_10_6 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_16_lut_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_16_lut_LC_11_10_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_16_lut_LC_11_10_6  (
            .in0(N__24138),
            .in1(N__28857),
            .in2(N__25184),
            .in3(N__24263),
            .lcout(\tok.n5520 ),
            .ltout(),
            .carryin(\tok.n4782 ),
            .carryout(\tok.n4783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_16_THRU_CRY_0_LC_11_10_7 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_16_THRU_CRY_0_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_16_THRU_CRY_0_LC_11_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \tok.sub_105_add_2_16_THRU_CRY_0_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__24226),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\tok.n4783 ),
            .carryout(\tok.n4783_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_17_lut_LC_11_11_0 .C_ON=1'b0;
    defparam \tok.sub_105_add_2_17_lut_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_17_lut_LC_11_11_0 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \tok.sub_105_add_2_17_lut_LC_11_11_0  (
            .in0(N__24758),
            .in1(N__24143),
            .in2(N__24872),
            .in3(N__24074),
            .lcout(\tok.n6_adj_783 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i16_1_lut_LC_11_11_1 .C_ON=1'b0;
    defparam \tok.inv_106_i16_1_lut_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i16_1_lut_LC_11_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i16_1_lut_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24846),
            .lcout(\tok.n287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i15_LC_11_11_2 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i15_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i15_LC_11_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.head_i0_i15_LC_11_11_2  (
            .in0(N__24847),
            .in1(N__24703),
            .in2(_gnd_net_),
            .in3(N__25514),
            .lcout(\tok.S_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28544),
            .ce(N__26078),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i15_LC_11_11_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i15_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i15_LC_11_11_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i15_LC_11_11_3  (
            .in0(N__24695),
            .in1(N__26602),
            .in2(_gnd_net_),
            .in3(N__24759),
            .lcout(\tok.A_stk.tail_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28544),
            .ce(N__26078),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i31_LC_11_11_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i31_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i31_LC_11_11_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i31_LC_11_11_4  (
            .in0(N__26603),
            .in1(N__24704),
            .in2(_gnd_net_),
            .in3(N__24686),
            .lcout(\tok.A_stk.tail_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28544),
            .ce(N__26078),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i47_LC_11_11_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i47_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i47_LC_11_11_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.tail_i0_i47_LC_11_11_5  (
            .in0(N__24694),
            .in1(N__26604),
            .in2(_gnd_net_),
            .in3(N__24650),
            .lcout(\tok.A_stk.tail_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28544),
            .ce(N__26078),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i63_LC_11_11_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i63_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i63_LC_11_11_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i63_LC_11_11_6  (
            .in0(N__26605),
            .in1(N__24685),
            .in2(_gnd_net_),
            .in3(N__24634),
            .lcout(\tok.A_stk.tail_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28544),
            .ce(N__26078),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i79_LC_11_11_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i79_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i79_LC_11_11_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i79_LC_11_11_7  (
            .in0(N__24677),
            .in1(N__26606),
            .in2(_gnd_net_),
            .in3(N__24649),
            .lcout(\tok.A_stk.tail_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28544),
            .ce(N__26078),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i90_LC_12_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i90_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i90_LC_12_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i90_LC_12_3_0  (
            .in0(N__25207),
            .in1(N__24982),
            .in2(_gnd_net_),
            .in3(N__26573),
            .lcout(\tok.A_stk.tail_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28521),
            .ce(N__26071),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i42_LC_12_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i42_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i42_LC_12_3_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i42_LC_12_3_1  (
            .in0(N__26570),
            .in1(_gnd_net_),
            .in2(N__24974),
            .in3(N__24952),
            .lcout(\tok.A_stk.tail_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28521),
            .ce(N__26071),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i74_LC_12_3_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i74_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i74_LC_12_3_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i74_LC_12_3_2  (
            .in0(N__25247),
            .in1(N__24970),
            .in2(_gnd_net_),
            .in3(N__26572),
            .lcout(\tok.A_stk.tail_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28521),
            .ce(N__26071),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i58_LC_12_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i58_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i58_LC_12_3_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i58_LC_12_3_3  (
            .in0(N__26571),
            .in1(_gnd_net_),
            .in2(N__24986),
            .in3(N__24961),
            .lcout(\tok.A_stk.tail_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28521),
            .ce(N__26071),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i26_LC_12_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i26_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i26_LC_12_3_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.A_stk.tail_i0_i26_LC_12_3_5  (
            .in0(N__26569),
            .in1(_gnd_net_),
            .in2(N__24944),
            .in3(N__24962),
            .lcout(\tok.A_stk.tail_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28521),
            .ce(N__26071),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i10_LC_12_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i10_LC_12_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i10_LC_12_3_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i10_LC_12_3_6  (
            .in0(N__24953),
            .in1(N__26568),
            .in2(_gnd_net_),
            .in3(N__27414),
            .lcout(\tok.A_stk.tail_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28521),
            .ce(N__26071),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i10_LC_12_3_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i10_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i10_LC_12_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i10_LC_12_3_7  (
            .in0(N__24940),
            .in1(N__25511),
            .in2(_gnd_net_),
            .in3(N__29282),
            .lcout(\tok.S_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28521),
            .ce(N__26071),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i101_LC_12_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i101_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i101_LC_12_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i101_LC_12_4_0  (
            .in0(N__24932),
            .in1(N__24892),
            .in2(_gnd_net_),
            .in3(N__26518),
            .lcout(tail_101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28526),
            .ce(N__25986),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i85_LC_12_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i85_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i85_LC_12_4_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i85_LC_12_4_1  (
            .in0(N__26525),
            .in1(N__24904),
            .in2(_gnd_net_),
            .in3(N__24880),
            .lcout(\tok.A_stk.tail_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28526),
            .ce(N__25986),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i69_LC_12_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i69_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i69_LC_12_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i69_LC_12_4_2  (
            .in0(N__24893),
            .in1(N__25273),
            .in2(_gnd_net_),
            .in3(N__26524),
            .lcout(\tok.A_stk.tail_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28526),
            .ce(N__25986),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i53_LC_12_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i53_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i53_LC_12_4_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i53_LC_12_4_3  (
            .in0(N__26522),
            .in1(N__25264),
            .in2(_gnd_net_),
            .in3(N__24881),
            .lcout(\tok.A_stk.tail_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28526),
            .ce(N__25986),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i37_LC_12_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i37_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i37_LC_12_4_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i37_LC_12_4_4  (
            .in0(N__25255),
            .in1(N__25274),
            .in2(_gnd_net_),
            .in3(N__26521),
            .lcout(\tok.A_stk.tail_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28526),
            .ce(N__25986),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i21_LC_12_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i21_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i21_LC_12_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i21_LC_12_4_5  (
            .in0(N__26520),
            .in1(N__25265),
            .in2(_gnd_net_),
            .in3(N__25390),
            .lcout(\tok.A_stk.tail_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28526),
            .ce(N__25986),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i5_LC_12_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i5_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i5_LC_12_4_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i5_LC_12_4_6  (
            .in0(N__25256),
            .in1(N__26523),
            .in2(_gnd_net_),
            .in3(N__27187),
            .lcout(\tok.A_stk.tail_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28526),
            .ce(N__25986),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i106_LC_12_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i106_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i106_LC_12_4_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i106_LC_12_4_7  (
            .in0(N__26519),
            .in1(N__25246),
            .in2(_gnd_net_),
            .in3(N__25235),
            .lcout(tail_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28526),
            .ce(N__25986),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_LC_12_5_0 .C_ON=1'b0;
    defparam \tok.i7_4_lut_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_LC_12_5_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i7_4_lut_LC_12_5_0  (
            .in0(N__25762),
            .in1(N__25009),
            .in2(N__28837),
            .in3(N__25168),
            .lcout(\tok.n23_adj_642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i15_1_lut_LC_12_5_1 .C_ON=1'b0;
    defparam \tok.inv_106_i15_1_lut_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i15_1_lut_LC_12_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i15_1_lut_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25761),
            .lcout(\tok.n288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i11_LC_12_5_2 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i11_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i11_LC_12_5_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i11_LC_12_5_2  (
            .in0(N__25594),
            .in1(N__25502),
            .in2(_gnd_net_),
            .in3(N__25169),
            .lcout(\tok.S_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28529),
            .ce(N__26060),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i14_LC_12_5_3 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i14_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i14_LC_12_5_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.head_i0_i14_LC_12_5_3  (
            .in0(N__25503),
            .in1(N__25082),
            .in2(_gnd_net_),
            .in3(N__25763),
            .lcout(\tok.S_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28529),
            .ce(N__26060),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i11_LC_12_5_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i11_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i11_LC_12_5_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i11_LC_12_5_4  (
            .in0(N__25586),
            .in1(N__26583),
            .in2(_gnd_net_),
            .in3(N__25010),
            .lcout(\tok.A_stk.tail_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28529),
            .ce(N__26060),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i27_LC_12_5_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i27_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i27_LC_12_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i27_LC_12_5_5  (
            .in0(N__26584),
            .in1(N__25595),
            .in2(_gnd_net_),
            .in3(N__25577),
            .lcout(\tok.A_stk.tail_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28529),
            .ce(N__26060),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i43_LC_12_5_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i43_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i43_LC_12_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i43_LC_12_5_6  (
            .in0(N__25585),
            .in1(N__25549),
            .in2(_gnd_net_),
            .in3(N__26585),
            .lcout(\tok.A_stk.tail_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28529),
            .ce(N__26060),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i59_LC_12_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i59_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i59_LC_12_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i59_LC_12_5_7  (
            .in0(N__26586),
            .in1(N__25576),
            .in2(_gnd_net_),
            .in3(N__25568),
            .lcout(\tok.A_stk.tail_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28529),
            .ce(N__26060),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_31_LC_12_6_0 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_31_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_31_LC_12_6_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \tok.i4_4_lut_adj_31_LC_12_6_0  (
            .in0(N__29733),
            .in1(N__25328),
            .in2(N__27196),
            .in3(N__27290),
            .lcout(\tok.n20_adj_648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i4_1_lut_LC_12_6_1 .C_ON=1'b0;
    defparam \tok.inv_106_i4_1_lut_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i4_1_lut_LC_12_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i4_1_lut_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29732),
            .lcout(\tok.n299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i3_LC_12_6_2 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i3_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i3_LC_12_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.head_i0_i3_LC_12_6_2  (
            .in0(N__29734),
            .in1(N__25282),
            .in2(_gnd_net_),
            .in3(N__25504),
            .lcout(\tok.S_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28534),
            .ce(N__26074),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i5_LC_12_6_3 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i5_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i5_LC_12_6_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \tok.A_stk.head_i0_i5_LC_12_6_3  (
            .in0(N__27291),
            .in1(_gnd_net_),
            .in2(N__25513),
            .in3(N__25394),
            .lcout(\tok.S_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28534),
            .ce(N__26074),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i3_LC_12_6_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i3_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i3_LC_12_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i3_LC_12_6_4  (
            .in0(N__26589),
            .in1(N__26645),
            .in2(_gnd_net_),
            .in3(N__25329),
            .lcout(\tok.A_stk.tail_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28534),
            .ce(N__26074),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i19_LC_12_6_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i19_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i19_LC_12_6_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \tok.A_stk.tail_i0_i19_LC_12_6_5  (
            .in0(N__26636),
            .in1(_gnd_net_),
            .in2(N__25286),
            .in3(N__26587),
            .lcout(\tok.A_stk.tail_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28534),
            .ce(N__26074),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i35_LC_12_6_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i35_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i35_LC_12_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i35_LC_12_6_6  (
            .in0(N__26588),
            .in1(N__26644),
            .in2(_gnd_net_),
            .in3(N__26092),
            .lcout(\tok.A_stk.tail_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28534),
            .ce(N__26074),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i51_LC_12_6_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i51_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i51_LC_12_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i51_LC_12_6_7  (
            .in0(N__26635),
            .in1(N__26627),
            .in2(_gnd_net_),
            .in3(N__26590),
            .lcout(\tok.A_stk.tail_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28534),
            .ce(N__26074),
            .sr(_gnd_net_));
    defparam \tok.i5240_3_lut_LC_12_7_0 .C_ON=1'b0;
    defparam \tok.i5240_3_lut_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5240_3_lut_LC_12_7_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \tok.i5240_3_lut_LC_12_7_0  (
            .in0(N__27886),
            .in1(N__26795),
            .in2(_gnd_net_),
            .in3(N__25742),
            .lcout(\tok.n5412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_112_LC_12_7_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_112_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_112_LC_12_7_1 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i1_4_lut_adj_112_LC_12_7_1  (
            .in0(N__27654),
            .in1(N__25817),
            .in2(N__25764),
            .in3(N__26764),
            .lcout(),
            .ltout(\tok.n13_adj_772_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_113_LC_12_7_2 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_113_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_113_LC_12_7_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i10_4_lut_adj_113_LC_12_7_2  (
            .in0(N__25811),
            .in1(N__25799),
            .in2(N__25784),
            .in3(N__25781),
            .lcout(),
            .ltout(\tok.n22_adj_773_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i15_LC_12_7_3 .C_ON=1'b0;
    defparam \tok.A_i15_LC_12_7_3 .SEQ_MODE=4'b1010;
    defparam \tok.A_i15_LC_12_7_3 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \tok.A_i15_LC_12_7_3  (
            .in0(N__28626),
            .in1(N__28850),
            .in2(N__25775),
            .in3(N__28667),
            .lcout(\tok.A_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28540),
            .ce(N__28301),
            .sr(N__28233));
    defparam \tok.A_i6_LC_12_7_5 .C_ON=1'b0;
    defparam \tok.A_i6_LC_12_7_5 .SEQ_MODE=4'b1010;
    defparam \tok.A_i6_LC_12_7_5 .LUT_INIT=16'b1111110001011100;
    LogicCell40 \tok.A_i6_LC_12_7_5  (
            .in0(N__26796),
            .in1(N__27180),
            .in2(N__28638),
            .in3(N__27002),
            .lcout(\tok.A_low_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28540),
            .ce(N__28301),
            .sr(N__28233));
    defparam \tok.i2_3_lut_adj_189_LC_12_7_6 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_189_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_189_LC_12_7_6 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \tok.i2_3_lut_adj_189_LC_12_7_6  (
            .in0(N__27885),
            .in1(N__27292),
            .in2(_gnd_net_),
            .in3(N__27653),
            .lcout(\tok.n14_adj_856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i5_LC_12_8_0 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i5_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i5_LC_12_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.uart.rx_data_i0_i5_LC_12_8_0  (
            .in0(N__25693),
            .in1(N__25616),
            .in2(_gnd_net_),
            .in3(N__27124),
            .lcout(uart_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28541),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_192_LC_12_8_1 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_192_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_192_LC_12_8_1 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \tok.i6_4_lut_adj_192_LC_12_8_1  (
            .in0(N__27195),
            .in1(N__27957),
            .in2(N__27125),
            .in3(N__28788),
            .lcout(\tok.n18_adj_860 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_4_lut_adj_190_LC_12_8_2 .C_ON=1'b0;
    defparam \tok.i8_4_lut_adj_190_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i8_4_lut_adj_190_LC_12_8_2 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \tok.i8_4_lut_adj_190_LC_12_8_2  (
            .in0(N__27113),
            .in1(N__26995),
            .in2(N__27107),
            .in3(N__27077),
            .lcout(),
            .ltout(\tok.n20_adj_857_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_193_LC_12_8_3 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_193_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_193_LC_12_8_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i10_4_lut_adj_193_LC_12_8_3  (
            .in0(N__27071),
            .in1(N__27056),
            .in2(N__27044),
            .in3(N__27041),
            .lcout(),
            .ltout(\tok.n22_adj_861_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5564_4_lut_LC_12_8_4 .C_ON=1'b0;
    defparam \tok.i5564_4_lut_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5564_4_lut_LC_12_8_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i5564_4_lut_LC_12_8_4  (
            .in0(N__27035),
            .in1(N__27026),
            .in2(N__27011),
            .in3(N__27008),
            .lcout(\tok.n5556 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_LC_12_8_5 .C_ON=1'b0;
    defparam \tok.i3_3_lut_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_LC_12_8_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \tok.i3_3_lut_LC_12_8_5  (
            .in0(N__26996),
            .in1(N__26891),
            .in2(_gnd_net_),
            .in3(N__26882),
            .lcout(\tok.n15_adj_670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5244_3_lut_LC_12_9_0 .C_ON=1'b0;
    defparam \tok.i5244_3_lut_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5244_3_lut_LC_12_9_0 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \tok.i5244_3_lut_LC_12_9_0  (
            .in0(N__27884),
            .in1(_gnd_net_),
            .in2(N__26829),
            .in3(N__29411),
            .lcout(\tok.n5416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_43_LC_12_9_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_43_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_43_LC_12_9_1 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i1_4_lut_adj_43_LC_12_9_1  (
            .in0(N__27656),
            .in1(N__26780),
            .in2(N__29441),
            .in3(N__26753),
            .lcout(),
            .ltout(\tok.n13_adj_674_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_LC_12_9_2 .C_ON=1'b0;
    defparam \tok.i10_4_lut_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_LC_12_9_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i10_4_lut_LC_12_9_2  (
            .in0(N__26660),
            .in1(N__27893),
            .in2(N__26654),
            .in3(N__26651),
            .lcout(),
            .ltout(\tok.n22_adj_676_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i9_LC_12_9_3 .C_ON=1'b0;
    defparam \tok.A_i9_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \tok.A_i9_LC_12_9_3 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \tok.A_i9_LC_12_9_3  (
            .in0(N__28648),
            .in1(N__28072),
            .in2(N__28547),
            .in3(N__27977),
            .lcout(\tok.A_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__28543),
            .ce(N__28292),
            .sr(N__28231));
    defparam \tok.i5496_4_lut_LC_12_9_4 .C_ON=1'b0;
    defparam \tok.i5496_4_lut_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5496_4_lut_LC_12_9_4 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \tok.i5496_4_lut_LC_12_9_4  (
            .in0(N__28071),
            .in1(N__28784),
            .in2(N__27986),
            .in3(N__29477),
            .lcout(\tok.n5542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_41_LC_12_9_5 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_41_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_41_LC_12_9_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i2_3_lut_adj_41_LC_12_9_5  (
            .in0(N__27785),
            .in1(N__27971),
            .in2(_gnd_net_),
            .in3(N__27958),
            .lcout(\tok.n14_adj_668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i45_3_lut_LC_12_9_6 .C_ON=1'b0;
    defparam \tok.i45_3_lut_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i45_3_lut_LC_12_9_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.i45_3_lut_LC_12_9_6  (
            .in0(N__27883),
            .in1(N__27784),
            .in2(_gnd_net_),
            .in3(N__27655),
            .lcout(\tok.n5372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_52_LC_12_10_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_52_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_52_LC_12_10_0 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \tok.i1_4_lut_adj_52_LC_12_10_0  (
            .in0(N__28935),
            .in1(N__28785),
            .in2(N__27554),
            .in3(N__29565),
            .lcout(\tok.n8_adj_689 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_61_LC_12_10_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_61_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_61_LC_12_10_1 .LUT_INIT=16'b0101000001110011;
    LogicCell40 \tok.i1_4_lut_adj_61_LC_12_10_1  (
            .in0(N__28786),
            .in1(N__27297),
            .in2(N__27448),
            .in3(N__28937),
            .lcout(\tok.n8_adj_702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i5_1_lut_LC_12_10_2 .C_ON=1'b0;
    defparam \tok.inv_106_i5_1_lut_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i5_1_lut_LC_12_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i5_1_lut_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29564),
            .lcout(\tok.n298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i6_1_lut_LC_12_10_3 .C_ON=1'b0;
    defparam \tok.inv_106_i6_1_lut_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i6_1_lut_LC_12_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i6_1_lut_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27296),
            .lcout(\tok.n297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5197_2_lut_LC_12_10_4 .C_ON=1'b0;
    defparam \tok.i5197_2_lut_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i5197_2_lut_LC_12_10_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i5197_2_lut_LC_12_10_4  (
            .in0(N__28936),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30032),
            .lcout(\tok.n5366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5225_2_lut_LC_12_10_5 .C_ON=1'b0;
    defparam \tok.i5225_2_lut_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i5225_2_lut_LC_12_10_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i5225_2_lut_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__29703),
            .in2(_gnd_net_),
            .in3(N__28938),
            .lcout(),
            .ltout(\tok.n5396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_4_lut_adj_183_LC_12_10_6 .C_ON=1'b0;
    defparam \tok.i6_4_lut_4_lut_adj_183_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_4_lut_adj_183_LC_12_10_6 .LUT_INIT=16'b0000111111101111;
    LogicCell40 \tok.i6_4_lut_4_lut_adj_183_LC_12_10_6  (
            .in0(N__29353),
            .in1(N__29566),
            .in2(N__29480),
            .in3(N__29179),
            .lcout(\tok.n18_adj_677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i9_1_lut_LC_12_10_7 .C_ON=1'b0;
    defparam \tok.inv_106_i9_1_lut_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i9_1_lut_LC_12_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i9_1_lut_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29407),
            .lcout(\tok.n294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_101_i15_2_lut_LC_12_11_1 .C_ON=1'b0;
    defparam \tok.or_101_i15_2_lut_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.or_101_i15_2_lut_LC_12_11_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.or_101_i15_2_lut_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__29354),
            .in2(_gnd_net_),
            .in3(N__29278),
            .lcout(),
            .ltout(\tok.n202_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_4_lut_LC_12_11_2 .C_ON=1'b0;
    defparam \tok.i6_4_lut_4_lut_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_4_lut_LC_12_11_2 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i6_4_lut_4_lut_LC_12_11_2  (
            .in0(N__29180),
            .in1(N__29066),
            .in2(N__28982),
            .in3(N__28977),
            .lcout(),
            .ltout(\tok.n18_adj_774_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5455_4_lut_LC_12_11_3 .C_ON=1'b0;
    defparam \tok.i5455_4_lut_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5455_4_lut_LC_12_11_3 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \tok.i5455_4_lut_LC_12_11_3  (
            .in0(N__28874),
            .in1(N__28858),
            .in2(N__28793),
            .in3(N__28787),
            .lcout(\tok.n5518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
