-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Dec 31 2020 10:49:40

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    tx : out std_logic;
    rx : in std_logic;
    reset : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__30609\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10130\ : std_logic;
signal \VCCG0\ : std_logic;
signal \tok.A_stk.tail_89\ : std_logic;
signal \tok.A_stk.tail_73\ : std_logic;
signal \tok.A_stk.tail_57\ : std_logic;
signal \tok.A_stk.tail_41\ : std_logic;
signal \tok.A_stk.tail_25\ : std_logic;
signal \tok.A_stk.tail_9\ : std_logic;
signal \tok.A_stk.tail_87\ : std_logic;
signal \tok.A_stk.tail_71\ : std_logic;
signal \tok.A_stk.tail_55\ : std_logic;
signal \tok.A_stk.tail_39\ : std_logic;
signal \tok.A_stk.tail_23\ : std_logic;
signal \tok.A_stk.tail_7\ : std_logic;
signal tail_123 : std_logic;
signal tail_107 : std_logic;
signal \tok.A_stk.tail_91\ : std_logic;
signal \tok.A_stk.tail_75\ : std_logic;
signal \tok.A_stk.tail_59\ : std_logic;
signal \tok.A_stk.tail_43\ : std_logic;
signal \tok.A_stk.tail_27\ : std_logic;
signal \tok.A_stk.tail_11\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \tok.uart.n3955\ : std_logic;
signal \tok.uart.n3956\ : std_logic;
signal \tok.uart.n3957\ : std_logic;
signal \tok.uart.n3958\ : std_logic;
signal \tok.uart.n3959\ : std_logic;
signal \tok.uart.n3960\ : std_logic;
signal \tok.uart.n3961\ : std_logic;
signal \tok.uart.n3962\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \tok.uart.txclkcounter_3\ : std_logic;
signal \tok.uart.txclkcounter_5\ : std_logic;
signal \tok.uart.txclkcounter_0\ : std_logic;
signal \tok.uart.txclkcounter_2\ : std_logic;
signal \tok.uart.txclkcounter_6\ : std_logic;
signal \tok.uart.txclkcounter_1\ : std_logic;
signal \tok.uart.txclkcounter_7\ : std_logic;
signal \tok.uart.txclkcounter_8\ : std_logic;
signal \tok.uart.txclkcounter_4\ : std_logic;
signal \tok.uart.n14_cascade_\ : std_logic;
signal \tok.uart.n15_adj_640\ : std_logic;
signal \txtick_cascade_\ : std_logic;
signal \tok.uart.n1081\ : std_logic;
signal \tok.uart.rxclkcounter_0\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \tok.uart.rxclkcounter_1\ : std_logic;
signal \tok.uart.n3968\ : std_logic;
signal \tok.uart.n3969\ : std_logic;
signal \tok.uart.rxclkcounter_3\ : std_logic;
signal \tok.uart.n3970\ : std_logic;
signal \tok.uart.rxclkcounter_4\ : std_logic;
signal \tok.uart.n3971\ : std_logic;
signal \tok.uart.n3972\ : std_logic;
signal \tok.uart.n3973\ : std_logic;
signal \tok.table_wr_data_8\ : std_logic;
signal \tok.table_wr_data_15\ : std_logic;
signal \tok.table_wr_data_14\ : std_logic;
signal \tok.table_wr_data_13\ : std_logic;
signal \tok.uart.n12\ : std_logic;
signal \tok.uart.rxclkcounter_6\ : std_logic;
signal \tok.uart.rxclkcounter_5\ : std_logic;
signal \tok.uart.rxclkcounter_2\ : std_logic;
signal \n795_cascade_\ : std_logic;
signal \tok.table_wr_data_9\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \tok.uart.n3963\ : std_logic;
signal \tok.uart.n3964\ : std_logic;
signal \tok.uart.n3965\ : std_logic;
signal \tok.uart.n3966\ : std_logic;
signal \tok.uart.n3967\ : std_logic;
signal n940 : std_logic;
signal \tok.A_stk.tail_16\ : std_logic;
signal \tok.A_stk.tail_32\ : std_logic;
signal \tok.A_stk.tail_48\ : std_logic;
signal \tok.A_stk.tail_64\ : std_logic;
signal \tok.A_stk.tail_80\ : std_logic;
signal \tok.A_stk.tail_0\ : std_logic;
signal \tok.A_stk.tail_94\ : std_logic;
signal \tok.A_stk.tail_78\ : std_logic;
signal \tok.A_stk.tail_62\ : std_logic;
signal \tok.A_stk.tail_46\ : std_logic;
signal \tok.A_stk.tail_30\ : std_logic;
signal \tok.A_stk.tail_14\ : std_logic;
signal \tok.A_stk.tail_88\ : std_logic;
signal \tok.A_stk.tail_72\ : std_logic;
signal \tok.A_stk.tail_56\ : std_logic;
signal \tok.A_stk.tail_40\ : std_logic;
signal \tok.A_stk.tail_24\ : std_logic;
signal \tok.A_stk.tail_8\ : std_logic;
signal tail_96 : std_logic;
signal tail_112 : std_logic;
signal tail_105 : std_logic;
signal tail_121 : std_logic;
signal tail_104 : std_logic;
signal tail_120 : std_logic;
signal tail_103 : std_logic;
signal tail_119 : std_logic;
signal \tok.table_wr_data_12\ : std_logic;
signal tail_122 : std_logic;
signal tail_106 : std_logic;
signal \tok.A_stk.tail_90\ : std_logic;
signal \tok.A_stk.tail_74\ : std_logic;
signal \tok.A_stk.tail_58\ : std_logic;
signal \tok.A_stk.tail_42\ : std_logic;
signal \tok.A_stk.tail_26\ : std_logic;
signal \tok.A_stk.tail_10\ : std_logic;
signal \tok.n2_adj_763\ : std_logic;
signal \tok.n13_adj_765_cascade_\ : std_logic;
signal \tok.n18_adj_767_cascade_\ : std_logic;
signal \tok.n20_adj_770_cascade_\ : std_logic;
signal \tok.A_15_N_113_7_cascade_\ : std_logic;
signal \tok.A_15_N_84_7\ : std_logic;
signal \tok.A_15_N_113_7\ : std_logic;
signal \tok.uart.sentbits_3\ : std_logic;
signal \tok.uart.sentbits_2\ : std_logic;
signal \tok.uart.n3994_cascade_\ : std_logic;
signal n795 : std_logic;
signal \tok.uart.n4506_cascade_\ : std_logic;
signal \tok.uart.rxclkcounter_6__N_477\ : std_logic;
signal \tok.uart.n4438\ : std_logic;
signal \tok.uart.n2\ : std_logic;
signal \tok.n16_adj_769\ : std_logic;
signal \tok.uart.bytephase_1\ : std_logic;
signal \tok.uart.bytephase_5\ : std_logic;
signal \tok.uart.bytephase_3\ : std_logic;
signal \tok.uart.bytephase_0\ : std_logic;
signal \tok.uart.bytephase_2\ : std_logic;
signal \tok.uart.n13_cascade_\ : std_logic;
signal \tok.uart.bytephase_4\ : std_logic;
signal \bytephase_5__N_510\ : std_logic;
signal rx_c : std_logic;
signal capture_9 : std_logic;
signal \tok.n4508_cascade_\ : std_logic;
signal \tok.n4680\ : std_logic;
signal \tok.n16_adj_660_cascade_\ : std_logic;
signal \tok.n4\ : std_logic;
signal \tok.n206_cascade_\ : std_logic;
signal \tok.n204_cascade_\ : std_logic;
signal \tok.n16_adj_699_cascade_\ : std_logic;
signal \tok.n4667\ : std_logic;
signal \tok.A_stk.tail_18\ : std_logic;
signal \tok.A_stk.tail_34\ : std_logic;
signal \tok.A_stk.tail_50\ : std_logic;
signal \tok.A_stk.tail_66\ : std_logic;
signal \tok.A_stk.tail_82\ : std_logic;
signal \tok.A_stk.tail_2\ : std_logic;
signal tail_110 : std_logic;
signal tail_126 : std_logic;
signal tail_98 : std_logic;
signal tail_114 : std_logic;
signal tail_125 : std_logic;
signal tail_109 : std_logic;
signal \tok.A_stk.tail_93\ : std_logic;
signal \tok.A_stk.tail_77\ : std_logic;
signal \tok.A_stk.tail_61\ : std_logic;
signal \tok.A_stk.tail_45\ : std_logic;
signal \tok.A_stk.tail_29\ : std_logic;
signal \tok.A_stk.tail_13\ : std_logic;
signal tail_118 : std_logic;
signal tail_102 : std_logic;
signal \tok.A_stk.tail_86\ : std_logic;
signal \tok.A_stk.tail_70\ : std_logic;
signal \tok.A_stk.tail_54\ : std_logic;
signal \tok.A_stk.tail_38\ : std_logic;
signal \tok.A_stk.tail_22\ : std_logic;
signal \tok.A_stk.tail_6\ : std_logic;
signal \tok.n20_adj_803_cascade_\ : std_logic;
signal \tok.key_rd_5\ : std_logic;
signal \tok.key_rd_3\ : std_logic;
signal \tok.key_rd_8\ : std_logic;
signal \tok.n28\ : std_logic;
signal \tok.n25_cascade_\ : std_logic;
signal \tok.n26\ : std_logic;
signal \tok.key_rd_14\ : std_logic;
signal \tok.key_rd_11\ : std_logic;
signal \tok.table_wr_data_11\ : std_logic;
signal \tok.key_rd_15\ : std_logic;
signal \tok.key_rd_9\ : std_logic;
signal \tok.table_wr_data_7\ : std_logic;
signal \tok.table_wr_data_4\ : std_logic;
signal \tok.table_wr_data_1\ : std_logic;
signal \tok.n15_adj_771\ : std_logic;
signal \tok.uart.n6_cascade_\ : std_logic;
signal \n23_cascade_\ : std_logic;
signal \tok.uart.sentbits_0\ : std_logic;
signal \tok.uart.sentbits_1\ : std_logic;
signal \tok.uart.n978\ : std_logic;
signal \tok.uart.n1083\ : std_logic;
signal capture_7 : std_logic;
signal capture_6 : std_logic;
signal txtick : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \tok.n3910\ : std_logic;
signal \tok.n300\ : std_logic;
signal \tok.n3911\ : std_logic;
signal \tok.n3912\ : std_logic;
signal \tok.n3913\ : std_logic;
signal \tok.n3914\ : std_logic;
signal \tok.n3915\ : std_logic;
signal \tok.n295\ : std_logic;
signal \tok.n6_adj_768\ : std_logic;
signal \tok.n3916\ : std_logic;
signal \tok.n3917\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \tok.n3918\ : std_logic;
signal \tok.n3919\ : std_logic;
signal \tok.n291\ : std_logic;
signal \tok.n3920\ : std_logic;
signal \tok.n290\ : std_logic;
signal \tok.n6_adj_701\ : std_logic;
signal \tok.n3921\ : std_logic;
signal \tok.n3922\ : std_logic;
signal \tok.n288\ : std_logic;
signal \tok.n3923\ : std_logic;
signal \GNDG0\ : std_logic;
signal \tok.n3924\ : std_logic;
signal \tok.n3924_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \tok.n292\ : std_logic;
signal \tok.n287\ : std_logic;
signal tail_124 : std_logic;
signal tail_108 : std_logic;
signal \tok.A_stk.tail_92\ : std_logic;
signal \tok.A_stk.tail_76\ : std_logic;
signal \tok.A_stk.tail_60\ : std_logic;
signal \tok.A_stk.tail_44\ : std_logic;
signal \tok.A_stk.tail_28\ : std_logic;
signal \tok.A_stk.tail_12\ : std_logic;
signal \tok.A_stk.tail_17\ : std_logic;
signal \tok.A_stk.tail_33\ : std_logic;
signal \tok.A_stk.tail_49\ : std_logic;
signal \tok.A_stk.tail_65\ : std_logic;
signal \tok.A_stk.tail_81\ : std_logic;
signal \tok.A_stk.tail_1\ : std_logic;
signal tail_115 : std_logic;
signal \tok.A_stk.tail_51\ : std_logic;
signal tail_117 : std_logic;
signal tail_101 : std_logic;
signal \tok.A_stk.tail_67\ : std_logic;
signal tail_99 : std_logic;
signal \tok.A_stk.tail_83\ : std_logic;
signal \tok.A_stk.tail_35\ : std_logic;
signal \tok.A_stk.tail_3\ : std_logic;
signal \tok.A_stk.tail_19\ : std_logic;
signal \tok.A_stk.tail_85\ : std_logic;
signal \tok.A_stk.tail_69\ : std_logic;
signal \tok.A_stk.tail_53\ : std_logic;
signal \tok.A_stk.tail_37\ : std_logic;
signal \tok.A_stk.tail_21\ : std_logic;
signal \tok.A_stk.tail_5\ : std_logic;
signal tail_116 : std_logic;
signal tail_100 : std_logic;
signal \tok.A_stk.tail_84\ : std_logic;
signal \tok.A_stk.tail_68\ : std_logic;
signal \tok.A_stk.tail_52\ : std_logic;
signal \tok.A_stk.tail_36\ : std_logic;
signal \tok.A_stk.tail_20\ : std_logic;
signal \tok.A_stk.tail_4\ : std_logic;
signal \tok.n23_adj_677\ : std_logic;
signal \tok.n24\ : std_logic;
signal \tok.n26_adj_805\ : std_logic;
signal \tok.n30_adj_824_cascade_\ : std_logic;
signal \tok.found_slot_N_145\ : std_logic;
signal \tok.n4642_cascade_\ : std_logic;
signal \tok.key_rd_13\ : std_logic;
signal \tok.n14_adj_804\ : std_logic;
signal \tok.n27_adj_734\ : std_logic;
signal \tok.key_rd_12\ : std_logic;
signal \tok.key_rd_10\ : std_logic;
signal \tok.n21_adj_714\ : std_logic;
signal \tok.key_rd_2\ : std_logic;
signal \tok.key_rd_7\ : std_logic;
signal \tok.n22\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \tok.n3940\ : std_logic;
signal \tok.n3941\ : std_logic;
signal \tok.n3942\ : std_logic;
signal \tok.n3943\ : std_logic;
signal \tok.n3944\ : std_logic;
signal \tok.n3945\ : std_logic;
signal \tok.n10_adj_764\ : std_logic;
signal \tok.n3946\ : std_logic;
signal \tok.n3947\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \tok.n3948\ : std_logic;
signal \tok.n3949\ : std_logic;
signal \tok.n3950\ : std_logic;
signal \tok.n3951\ : std_logic;
signal \tok.n3952\ : std_logic;
signal \tok.n3953\ : std_logic;
signal \tok.n3954\ : std_logic;
signal \tok.n2_adj_739_cascade_\ : std_logic;
signal \tok.n6_adj_753\ : std_logic;
signal \tok.n14_adj_741_cascade_\ : std_logic;
signal \tok.n13_adj_748\ : std_logic;
signal \tok.n4656\ : std_logic;
signal \tok.n20_adj_754_cascade_\ : std_logic;
signal \tok.n9_adj_749\ : std_logic;
signal \tok.table_rd_15\ : std_logic;
signal \tok.n16_adj_751\ : std_logic;
signal \tok.n17_adj_774\ : std_logic;
signal \tok.n10_adj_705\ : std_logic;
signal \tok.n6_adj_692\ : std_logic;
signal \tok.n13_adj_688_cascade_\ : std_logic;
signal \tok.n12_adj_687\ : std_logic;
signal \tok.n4674\ : std_logic;
signal \tok.n20_adj_693_cascade_\ : std_logic;
signal \tok.n6_adj_667\ : std_logic;
signal \tok.n294\ : std_logic;
signal \tok.table_wr_data_3\ : std_logic;
signal \tok.n298\ : std_logic;
signal \tok.n289\ : std_logic;
signal \tok.n6_adj_814\ : std_logic;
signal \tok.n34_cascade_\ : std_logic;
signal \tok.n13\ : std_logic;
signal \tok.n2_adj_685_cascade_\ : std_logic;
signal \tok.n14_adj_686\ : std_logic;
signal sender_1 : std_logic;
signal tx_c : std_logic;
signal reset_c : std_logic;
signal \tok.A_stk.tail_63\ : std_logic;
signal \tok.A_stk.tail_47\ : std_logic;
signal \tok.A_stk.tail_31\ : std_logic;
signal \tok.A_stk.tail_15\ : std_logic;
signal \tok.A_stk.tail_79\ : std_logic;
signal \tok.A_stk.tail_95\ : std_logic;
signal tail_111 : std_logic;
signal tail_127 : std_logic;
signal tail_97 : std_logic;
signal tail_113 : std_logic;
signal n29 : std_logic;
signal \n29_cascade_\ : std_logic;
signal \tok.A_stk.rd_15__N_301\ : std_logic;
signal \tok.n83_adj_735_cascade_\ : std_logic;
signal \tok.n7_cascade_\ : std_logic;
signal \tok.n4516\ : std_logic;
signal capture_0 : std_logic;
signal \tok.n17\ : std_logic;
signal \tok.n4_adj_654_cascade_\ : std_logic;
signal n786 : std_logic;
signal \tok.n83_adj_716_cascade_\ : std_logic;
signal \tok.n12_adj_740_cascade_\ : std_logic;
signal \tok.n12_adj_801_cascade_\ : std_logic;
signal \tok.n284\ : std_logic;
signal \tok.n284_cascade_\ : std_logic;
signal \tok.n182_cascade_\ : std_logic;
signal \tok.n12_adj_766\ : std_logic;
signal \tok.n24_adj_854\ : std_logic;
signal \tok.n21_adj_857\ : std_logic;
signal \tok.n30_adj_862_cascade_\ : std_logic;
signal \tok.n19_adj_860_cascade_\ : std_logic;
signal \tok.n17_adj_861\ : std_logic;
signal \tok.n29_adj_864\ : std_logic;
signal capture_8 : std_logic;
signal uart_rx_data_7 : std_logic;
signal \tok.table_wr_data_10\ : std_logic;
signal \tok.n293\ : std_logic;
signal \tok.n2634\ : std_logic;
signal \tok.write_slot\ : std_logic;
signal \tok.table_wr_data_5\ : std_logic;
signal \tok.key_rd_4\ : std_logic;
signal \tok.key_rd_1\ : std_logic;
signal \tok.n18_adj_756\ : std_logic;
signal \tok.key_rd_0\ : std_logic;
signal \tok.key_rd_6\ : std_logic;
signal \tok.n4645\ : std_logic;
signal \tok.n13_adj_657\ : std_logic;
signal \tok.n10_adj_656\ : std_logic;
signal \tok.table_rd_9\ : std_logic;
signal \tok.n30_cascade_\ : std_logic;
signal \tok.n12_adj_659\ : std_logic;
signal \tok.uart.n922\ : std_logic;
signal \tok.n301\ : std_logic;
signal \tok.n15_cascade_\ : std_logic;
signal \tok.n183\ : std_logic;
signal \tok.table_rd_6\ : std_logic;
signal \tok.n16_adj_778_cascade_\ : std_logic;
signal \tok.n6_adj_780\ : std_logic;
signal \tok.table_rd_13\ : std_logic;
signal \tok.table_rd_10\ : std_logic;
signal \tok.n10_adj_671\ : std_logic;
signal \tok.n14_adj_669_cascade_\ : std_logic;
signal \tok.table_rd_11\ : std_logic;
signal \tok.n16_adj_691\ : std_logic;
signal \tok.n4653\ : std_logic;
signal \tok.n4671\ : std_logic;
signal \tok.n18_adj_672\ : std_logic;
signal \tok.n6_adj_676\ : std_logic;
signal \tok.n20_adj_674_cascade_\ : std_logic;
signal \tok.n16_adj_673\ : std_logic;
signal \tok.n4676_cascade_\ : std_logic;
signal \tok.n12_adj_744\ : std_logic;
signal \tok.n4524\ : std_logic;
signal \tok.n12_adj_670\ : std_logic;
signal \tok.n2_adj_720_cascade_\ : std_logic;
signal \tok.n14_adj_722\ : std_logic;
signal \tok.n6_adj_731\ : std_logic;
signal \tok.n13_adj_726_cascade_\ : std_logic;
signal \tok.n12_adj_723\ : std_logic;
signal \tok.n4661\ : std_logic;
signal \tok.n20_adj_732_cascade_\ : std_logic;
signal \tok.n4658\ : std_logic;
signal \tok.n9_adj_728\ : std_logic;
signal \tok.n184\ : std_logic;
signal uart_rx_data_5 : std_logic;
signal \tok.n12_adj_815_cascade_\ : std_logic;
signal \tok.n16_adj_820\ : std_logic;
signal \tok.n20_adj_822_cascade_\ : std_logic;
signal \tok.A_15_N_113_5_cascade_\ : std_logic;
signal \tok.n297\ : std_logic;
signal \tok.n208\ : std_logic;
signal \tok.n20_adj_858\ : std_logic;
signal \tok.n299\ : std_logic;
signal \tok.n27_adj_644_cascade_\ : std_logic;
signal \tok.tail_9\ : std_logic;
signal \tok.C_stk.tail_17\ : std_logic;
signal \tok.tail_25\ : std_logic;
signal \tok.C_stk.tail_33\ : std_logic;
signal \tok.tail_57\ : std_logic;
signal \tok.tail_41\ : std_logic;
signal \tok.tail_49\ : std_logic;
signal \tok.tail_58\ : std_logic;
signal \tok.n875_cascade_\ : std_logic;
signal \tok.n2562\ : std_logic;
signal \tok.n2503\ : std_logic;
signal \tok.n2562_cascade_\ : std_logic;
signal \tok.n4474_cascade_\ : std_logic;
signal \tok.n875\ : std_logic;
signal \tok.n20_adj_772_cascade_\ : std_logic;
signal \tok.n63\ : std_logic;
signal \tok.A_stk_delta_1__N_4_cascade_\ : std_logic;
signal \tok.n61\ : std_logic;
signal \tok.n4_adj_809_cascade_\ : std_logic;
signal \tok.depth_3_cascade_\ : std_logic;
signal \tok.depth_1\ : std_logic;
signal \tok.n4554_cascade_\ : std_logic;
signal \tok.n237\ : std_logic;
signal \tok.n6_adj_832\ : std_logic;
signal \tok.n4504\ : std_logic;
signal \tok.n4432_cascade_\ : std_logic;
signal \tok.A_stk_delta_1__N_4\ : std_logic;
signal \tok.n1_adj_802_cascade_\ : std_logic;
signal \tok.n189\ : std_logic;
signal \tok.n62\ : std_logic;
signal \tok.n189_cascade_\ : std_logic;
signal \tok.n4_adj_809\ : std_logic;
signal \tok.n27_adj_793_cascade_\ : std_logic;
signal \tok.n25_adj_794\ : std_logic;
signal \tok.n26_adj_792\ : std_logic;
signal \tok.n28_adj_791\ : std_logic;
signal \tok.n18_adj_859\ : std_logic;
signal \tok.n22_adj_855\ : std_logic;
signal \tok.n880\ : std_logic;
signal \tok.n23_cascade_\ : std_logic;
signal \tok.n23_adj_856\ : std_logic;
signal \tok.n64\ : std_logic;
signal \tok.n1_adj_802\ : std_logic;
signal \tok.depth_2\ : std_logic;
signal \tok.depth_0_cascade_\ : std_logic;
signal \tok.n6_adj_853\ : std_logic;
signal \tok.A__15__N_129_cascade_\ : std_logic;
signal \tok.n27_adj_867_cascade_\ : std_logic;
signal \tok.n1\ : std_logic;
signal \tok.n14_adj_678_cascade_\ : std_logic;
signal \tok.n2\ : std_logic;
signal \tok.n19_cascade_\ : std_logic;
signal \tok.n6_adj_684\ : std_logic;
signal \tok.n22_adj_683_cascade_\ : std_logic;
signal \tok.n4544\ : std_logic;
signal \tok.A_15_N_113_0_cascade_\ : std_logic;
signal \tok.n4520\ : std_logic;
signal \tok.n46_cascade_\ : std_logic;
signal \tok.A_15_N_113_1\ : std_logic;
signal \tok.A_15_N_113_1_cascade_\ : std_logic;
signal \tok.A_1_cascade_\ : std_logic;
signal \tok.uart.sender_3\ : std_logic;
signal \tok.A_0\ : std_logic;
signal sender_2 : std_logic;
signal \tok.A_2\ : std_logic;
signal \tok.uart.sender_4\ : std_logic;
signal \tok.n10_adj_783\ : std_logic;
signal \tok.n14_adj_779_cascade_\ : std_logic;
signal \tok.n20_adj_781\ : std_logic;
signal \tok.n22_adj_784_cascade_\ : std_logic;
signal \tok.A_15_N_113_6_cascade_\ : std_logic;
signal \tok.A_6_cascade_\ : std_logic;
signal \tok.uart.sender_9\ : std_logic;
signal \tok.uart.sender_8\ : std_logic;
signal \tok.A_5\ : std_logic;
signal \tok.uart.sender_7\ : std_logic;
signal \tok.uart.sender_6\ : std_logic;
signal n23 : std_logic;
signal \tok.uart.sender_5\ : std_logic;
signal \tok.uart.n964\ : std_logic;
signal \tok.n16_adj_706\ : std_logic;
signal \tok.n14_adj_707\ : std_logic;
signal \tok.n20_adj_708_cascade_\ : std_logic;
signal \tok.n22_adj_709_cascade_\ : std_logic;
signal \tok.A_15_N_113_5\ : std_logic;
signal \tok.n10_adj_806\ : std_logic;
signal \tok.n13_adj_813_cascade_\ : std_logic;
signal \tok.n18_adj_819\ : std_logic;
signal \tok.n15_adj_823\ : std_logic;
signal \tok.n27_adj_863_cascade_\ : std_logic;
signal \tok.n27_adj_865_cascade_\ : std_logic;
signal \tok.n27_adj_664\ : std_logic;
signal \tok.n27_adj_866\ : std_logic;
signal \tok.tail_50\ : std_logic;
signal \tok.C_stk.tail_34\ : std_logic;
signal \tok.tail_42\ : std_logic;
signal \tok.tail_28\ : std_logic;
signal \tok.n127_cascade_\ : std_logic;
signal \tok.n4446\ : std_logic;
signal \tok.n4394_cascade_\ : std_logic;
signal \tok.n28_adj_834_cascade_\ : std_logic;
signal \tok.n4604_cascade_\ : std_logic;
signal \tok.n34_adj_719\ : std_logic;
signal \tok.n4610_cascade_\ : std_logic;
signal \tok.n37\ : std_logic;
signal \tok.table_rd_7\ : std_logic;
signal \tok.n83_adj_796_cascade_\ : std_logic;
signal capture_3 : std_logic;
signal \tok.n847\ : std_logic;
signal \tok.n31\ : std_logic;
signal \tok.C_stk.n4906_cascade_\ : std_logic;
signal \tok.ram.n4699_cascade_\ : std_logic;
signal \tok.n4649\ : std_logic;
signal \tok.n1_adj_760_cascade_\ : std_logic;
signal \tok.n13_adj_761_cascade_\ : std_logic;
signal \tok.tc_7\ : std_logic;
signal \tok.C_stk.tail_1\ : std_logic;
signal \tok.C_stk.n4870_cascade_\ : std_logic;
signal \tok.ram.n4714_cascade_\ : std_logic;
signal \tok.c_stk_r_1\ : std_logic;
signal \tok.n4690\ : std_logic;
signal \tok.n1_adj_717_cascade_\ : std_logic;
signal \tok.n5_adj_718_cascade_\ : std_logic;
signal \n92_cascade_\ : std_logic;
signal \tok.tc_1\ : std_logic;
signal \tok.n28_adj_821\ : std_logic;
signal \tok.n10_adj_786\ : std_logic;
signal \tok.n6_adj_848_cascade_\ : std_logic;
signal \tok.n32_cascade_\ : std_logic;
signal uart_rx_data_1 : std_logic;
signal \tok.table_wr_data_6\ : std_logic;
signal capture_2 : std_logic;
signal n4005 : std_logic;
signal \tok.table_wr_data_2\ : std_logic;
signal \tok.n18_adj_844_cascade_\ : std_logic;
signal \tok.n16_adj_845\ : std_logic;
signal \tok.n20_adj_846_cascade_\ : std_logic;
signal \tok.A_15_N_113_2\ : std_logic;
signal \tok.n15_adj_847\ : std_logic;
signal uart_rx_data_2 : std_logic;
signal \tok.n12_adj_843\ : std_logic;
signal capture_1 : std_logic;
signal uart_rx_data_0 : std_logic;
signal \tok.table_rd_14\ : std_logic;
signal \tok.n16_adj_730\ : std_logic;
signal \tok.n400\ : std_logic;
signal \tok.table_wr_data_0\ : std_logic;
signal \tok.n2614\ : std_logic;
signal \tok.n2614_cascade_\ : std_logic;
signal \tok.n2616_cascade_\ : std_logic;
signal \tok.n10_adj_849\ : std_logic;
signal \tok.n12_adj_851\ : std_logic;
signal \tok.table_rd_1\ : std_logic;
signal \tok.n8_adj_850\ : std_logic;
signal \tok.A_4\ : std_logic;
signal \tok.n4051\ : std_logic;
signal \tok.A_15_N_113_4\ : std_logic;
signal \tok.A_15_N_113_4_cascade_\ : std_logic;
signal \tok.A_15_N_113_0\ : std_logic;
signal \tok.A_15_N_113_6\ : std_logic;
signal \tok.n23\ : std_logic;
signal \tok.n950\ : std_logic;
signal \tok.A__15__N_129\ : std_logic;
signal \tok.A_15_N_113_3\ : std_logic;
signal \tok.A_3\ : std_logic;
signal \tok.n4528_cascade_\ : std_logic;
signal \tok.n892_cascade_\ : std_logic;
signal \tok.n10_adj_818\ : std_logic;
signal \tok.n13_adj_842\ : std_logic;
signal \tok.n8_adj_666\ : std_logic;
signal \tok.n8_adj_777\ : std_logic;
signal \tok.n4502_cascade_\ : std_logic;
signal \tok.n12_adj_830\ : std_logic;
signal \tok.n4607\ : std_logic;
signal \tok.n9_adj_689\ : std_logic;
signal \tok.n181_cascade_\ : std_logic;
signal \tok.n12_cascade_\ : std_logic;
signal \tok.n6_adj_653\ : std_logic;
signal \tok.n20_cascade_\ : std_logic;
signal \tok.n16\ : std_logic;
signal \tok.n4684\ : std_logic;
signal \tok.n892\ : std_logic;
signal \tok.n177_cascade_\ : std_logic;
signal \tok.n12_adj_696_cascade_\ : std_logic;
signal \tok.n20_adj_700\ : std_logic;
signal \tok.n52\ : std_logic;
signal \tok.n33_adj_663\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \tok.n50\ : std_logic;
signal \tok.n33_adj_841\ : std_logic;
signal \tok.n3888\ : std_logic;
signal \tok.n49\ : std_logic;
signal \tok.n33_adj_665\ : std_logic;
signal \tok.n3889\ : std_logic;
signal \tok.n47\ : std_logic;
signal \tok.n33_adj_755\ : std_logic;
signal \tok.n3890\ : std_logic;
signal \tok.n45\ : std_logic;
signal \tok.n33_adj_852\ : std_logic;
signal \tok.n3891\ : std_logic;
signal \tok.n44\ : std_logic;
signal \tok.n3892\ : std_logic;
signal \tok.n3893\ : std_logic;
signal \tok.n39\ : std_logic;
signal \tok.n3894\ : std_logic;
signal \tok.n33_adj_643\ : std_logic;
signal \tok.C_stk.tail_20\ : std_logic;
signal \tok.tail_26\ : std_logic;
signal \tok.tail_12\ : std_logic;
signal \tok.C_stk.tail_36\ : std_logic;
signal \tok.tail_56\ : std_logic;
signal \tok.tail_40\ : std_logic;
signal \tok.tail_48\ : std_logic;
signal \tok.n83_adj_704\ : std_logic;
signal \tok.n4694_cascade_\ : std_logic;
signal \tok.n13_adj_713_cascade_\ : std_logic;
signal \tok.C_stk.n4894_cascade_\ : std_logic;
signal \tok.c_stk_r_0\ : std_logic;
signal \tok.ram.n4717_cascade_\ : std_logic;
signal \tok.n1_adj_712\ : std_logic;
signal \tok.C_stk.tail_7\ : std_logic;
signal \tok.C_stk.n4912_cascade_\ : std_logic;
signal \tok.tc_6\ : std_logic;
signal \tok.c_stk_r_7\ : std_logic;
signal \tok.ram.n4696_cascade_\ : std_logic;
signal \tok.n4602\ : std_logic;
signal \tok.n1_adj_798_cascade_\ : std_logic;
signal \tok.n13_adj_799\ : std_logic;
signal \tok.tc_0\ : std_logic;
signal \tok.tc_plus_1_0\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \tok.tc_plus_1_1\ : std_logic;
signal \tok.n3895\ : std_logic;
signal \tok.n3896\ : std_logic;
signal \tok.n3897\ : std_logic;
signal \tok.n3898\ : std_logic;
signal \tok.n3899\ : std_logic;
signal \tok.tc_plus_1_6\ : std_logic;
signal \tok.n3900\ : std_logic;
signal \tok.n3901\ : std_logic;
signal \tok.tc_plus_1_7\ : std_logic;
signal n92_adj_872 : std_logic;
signal \c_stk_w_7_N_18_7\ : std_logic;
signal n92_adj_871 : std_logic;
signal \c_stk_w_7_N_18_6\ : std_logic;
signal n92 : std_logic;
signal \c_stk_w_7_N_18_1\ : std_logic;
signal n10_adj_875 : std_logic;
signal \c_stk_w_7_N_18_0\ : std_logic;
signal \tok.found_slot\ : std_logic;
signal \tok.n5_adj_655_cascade_\ : std_logic;
signal \tok.uart_tx_busy\ : std_logic;
signal \tok.uart_rx_valid\ : std_logic;
signal \tok.uart_stall_cascade_\ : std_logic;
signal \tok.n2732\ : std_logic;
signal \tok.n2732_cascade_\ : std_logic;
signal \tok.n43\ : std_logic;
signal \tok.n5_adj_655\ : std_logic;
signal \tok.reset_N_2\ : std_logic;
signal \tok.uart_stall\ : std_logic;
signal \tok.n2724\ : std_logic;
signal \tok.n4431\ : std_logic;
signal \tok.n5_adj_682\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \tok.S_1\ : std_logic;
signal \tok.n4_adj_790\ : std_logic;
signal \tok.n3925\ : std_logic;
signal \tok.S_2\ : std_logic;
signal \tok.n5_adj_789\ : std_logic;
signal \tok.n3926\ : std_logic;
signal \tok.n3927\ : std_logic;
signal \tok.n3928\ : std_logic;
signal \tok.S_5\ : std_logic;
signal \tok.n5_adj_775\ : std_logic;
signal \tok.n3929\ : std_logic;
signal \tok.n5_adj_773\ : std_logic;
signal \tok.n3930\ : std_logic;
signal \tok.A_low_7\ : std_logic;
signal \tok.S_7\ : std_logic;
signal \tok.n5_adj_752\ : std_logic;
signal \tok.n3931\ : std_logic;
signal \tok.n3932\ : std_logic;
signal \tok.S_8\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \tok.S_9\ : std_logic;
signal \tok.n21\ : std_logic;
signal \tok.n3933\ : std_logic;
signal \tok.n58\ : std_logic;
signal \tok.S_10\ : std_logic;
signal \tok.n5_adj_668\ : std_logic;
signal \tok.n3934\ : std_logic;
signal \tok.S_11\ : std_logic;
signal \tok.n5_adj_690\ : std_logic;
signal \tok.n3935\ : std_logic;
signal \tok.S_12\ : std_logic;
signal \tok.n3936\ : std_logic;
signal \tok.n55\ : std_logic;
signal \tok.S_13\ : std_logic;
signal \tok.n3937\ : std_logic;
signal \tok.S_14\ : std_logic;
signal \tok.n5_adj_729\ : std_logic;
signal \tok.n3938\ : std_logic;
signal \tok.S_15\ : std_logic;
signal \tok.n53\ : std_logic;
signal \tok.n3939\ : std_logic;
signal \tok.n5_adj_750\ : std_logic;
signal \tok.n6_adj_812\ : std_logic;
signal \tok.n9_adj_836\ : std_logic;
signal \tok.n5_adj_837_cascade_\ : std_logic;
signal \tok.S_3\ : std_logic;
signal \tok.n23_adj_788\ : std_logic;
signal \tok.n10_adj_838_cascade_\ : std_logic;
signal \tok.n12_adj_840\ : std_logic;
signal \tok.n57\ : std_logic;
signal \tok.n6_adj_835\ : std_logic;
signal uart_rx_data_6 : std_logic;
signal \tok.n109_cascade_\ : std_logic;
signal \tok.S_6\ : std_logic;
signal \tok.n18_adj_782\ : std_logic;
signal capture_4 : std_logic;
signal uart_rx_data_3 : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \tok.n13_adj_816\ : std_logic;
signal \tok.n3902\ : std_logic;
signal \tok.n2_adj_811\ : std_logic;
signal \tok.n3903\ : std_logic;
signal \tok.n26_adj_808\ : std_logic;
signal \tok.n3904\ : std_logic;
signal \tok.n3905\ : std_logic;
signal \tok.n3906\ : std_logic;
signal \tok.A_low_2\ : std_logic;
signal \tok.n210\ : std_logic;
signal \tok.n3907\ : std_logic;
signal \tok.A_low_3\ : std_logic;
signal \tok.n209\ : std_logic;
signal \tok.n3908\ : std_logic;
signal \tok.n3909\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \tok.n2598\ : std_logic;
signal \tok.n211\ : std_logic;
signal \tok.n2_adj_810\ : std_logic;
signal \tok.n5_adj_710\ : std_logic;
signal \tok.n6_adj_711\ : std_logic;
signal \tok.n4664\ : std_logic;
signal \tok.n4663\ : std_logic;
signal \tok.n33\ : std_logic;
signal \tok.n27\ : std_logic;
signal \tok.n296\ : std_logic;
signal \tok.n191\ : std_logic;
signal \tok.n59\ : std_logic;
signal \tok.n2_adj_703\ : std_logic;
signal \tok.stall\ : std_logic;
signal \tok.A_low_5\ : std_logic;
signal \tok.search_clk\ : std_logic;
signal \tok.n33_adj_817\ : std_logic;
signal \tok.n27_adj_868\ : std_logic;
signal \tok.n82\ : std_logic;
signal capture_5 : std_logic;
signal \rx_data_7__N_511\ : std_logic;
signal \tok.n9_adj_807\ : std_logic;
signal uart_rx_data_4 : std_logic;
signal \tok.n3_adj_826\ : std_logic;
signal \tok.n6_adj_827_cascade_\ : std_logic;
signal \tok.n36\ : std_logic;
signal \tok.n33_adj_828_cascade_\ : std_logic;
signal \tok.n11_adj_831\ : std_logic;
signal \tok.n56\ : std_logic;
signal \tok.n2514\ : std_logic;
signal \tok.C_stk.tail_0\ : std_logic;
signal \tok.tail_8\ : std_logic;
signal \tok.tail_15\ : std_logic;
signal \tok.C_stk.tail_23\ : std_logic;
signal \tok.tail_31\ : std_logic;
signal \tok.C_stk.tail_39\ : std_logic;
signal \tok.tail_47\ : std_logic;
signal \tok.C_stk.tail_16\ : std_logic;
signal \tok.C_stk.tail_32\ : std_logic;
signal \tok.tail_24\ : std_logic;
signal \tok.tail_30\ : std_logic;
signal \tok.C_stk.tail_38\ : std_logic;
signal \tok.tail_46\ : std_logic;
signal \tok.c_stk_r_6\ : std_logic;
signal \tok.tail_44\ : std_logic;
signal \tok.C_stk.tail_18\ : std_logic;
signal \tok.n240\ : std_logic;
signal \tok.tail_55\ : std_logic;
signal \tok.tail_63\ : std_logic;
signal \tok.tail_54\ : std_logic;
signal \tok.tail_62\ : std_logic;
signal \tok.tail_52\ : std_logic;
signal \tok.tail_60\ : std_logic;
signal \tok.C_stk.n4900_cascade_\ : std_logic;
signal \tok.table_rd_5\ : std_logic;
signal \tok.n83_adj_742_cascade_\ : std_logic;
signal \tok.n4651_cascade_\ : std_logic;
signal \tok.ram.n4702_cascade_\ : std_logic;
signal \tok.n1_adj_757\ : std_logic;
signal \tok.tc_plus_1_5\ : std_logic;
signal \tok.n13_adj_758\ : std_logic;
signal n10_adj_873 : std_logic;
signal \n10_adj_873_cascade_\ : std_logic;
signal \c_stk_w_7_N_18_5\ : std_logic;
signal \tok.tc_5\ : std_logic;
signal n10_adj_874 : std_logic;
signal \n10_adj_874_cascade_\ : std_logic;
signal \tok.tc_2\ : std_logic;
signal \tok.tc_plus_1_3\ : std_logic;
signal n92_adj_870 : std_logic;
signal \n92_adj_870_cascade_\ : std_logic;
signal \c_stk_w_7_N_18_3\ : std_logic;
signal \tok.tc_3\ : std_logic;
signal \stall_\ : std_logic;
signal \tok.tc_4\ : std_logic;
signal \tok.n9_adj_797\ : std_logic;
signal \tok.n11_adj_647\ : std_logic;
signal \tok.n4575_cascade_\ : std_logic;
signal \tok.n83_cascade_\ : std_logic;
signal \tok.n40\ : std_logic;
signal \tok.n4571_cascade_\ : std_logic;
signal \tok.n4393\ : std_logic;
signal \tok.n4460_cascade_\ : std_logic;
signal \tok.n2726\ : std_logic;
signal \tok.S_4\ : std_logic;
signal \tok.n13_adj_787\ : std_logic;
signal \tok.n10_adj_829_cascade_\ : std_logic;
signal \tok.n13_adj_833\ : std_logic;
signal \tok.n2746\ : std_logic;
signal \tok.n8_adj_839\ : std_logic;
signal \tok.table_rd_0\ : std_logic;
signal \tok.n18_adj_681\ : std_logic;
signal \tok.A_low_1\ : std_logic;
signal \tok.n101\ : std_logic;
signal \tok.n54\ : std_logic;
signal \tok.n244_cascade_\ : std_logic;
signal \tok.n17_adj_785\ : std_logic;
signal \tok.n60\ : std_logic;
signal \tok.n83\ : std_logic;
signal \tok.n3\ : std_logic;
signal \tok.n4478\ : std_logic;
signal \tok.c_stk_r_5\ : std_logic;
signal \tok.C_stk.tail_5\ : std_logic;
signal \tok.tail_13\ : std_logic;
signal \tok.C_stk.tail_21\ : std_logic;
signal \tok.tail_29\ : std_logic;
signal \tok.C_stk.tail_37\ : std_logic;
signal \tok.tail_61\ : std_logic;
signal \tok.tail_45\ : std_logic;
signal \tok.tail_53\ : std_logic;
signal \tok.C_stk.tail_22\ : std_logic;
signal \tok.C_stk.tail_6\ : std_logic;
signal \tok.tail_14\ : std_logic;
signal \tok.tail_11\ : std_logic;
signal \tok.C_stk.tail_19\ : std_logic;
signal \tok.tail_27\ : std_logic;
signal \tok.C_stk.tail_35\ : std_logic;
signal \tok.tail_59\ : std_logic;
signal \tok.tail_43\ : std_logic;
signal \tok.tail_51\ : std_logic;
signal \tok.tail_10\ : std_logic;
signal \tok.C_stk_delta_1\ : std_logic;
signal \tok.rd_7__N_374\ : std_logic;
signal \c_stk_w_7_N_18_4\ : std_logic;
signal \tok.C_stk.tail_4\ : std_logic;
signal \tok.C_stk.n4888_cascade_\ : std_logic;
signal \tok.ram.n4705_cascade_\ : std_logic;
signal \tok.n1_adj_745_cascade_\ : std_logic;
signal \tok.tc_plus_1_4\ : std_logic;
signal \tok.n802\ : std_logic;
signal \tok.n13_adj_746_cascade_\ : std_logic;
signal \tok.n86\ : std_logic;
signal n10 : std_logic;
signal \tok.C_stk.tail_3\ : std_logic;
signal \tok.C_stk.n4882\ : std_logic;
signal \tok.n602\ : std_logic;
signal \c_stk_w_7_N_18_2\ : std_logic;
signal \tok.C_stk.tail_2\ : std_logic;
signal \tok.C_stk.n4876_cascade_\ : std_logic;
signal \tok.C_stk.n600\ : std_logic;
signal clk : std_logic;
signal \tok.tc_plus_1_2\ : std_logic;
signal \tok.tc__7__N_134\ : std_logic;
signal \tok.ram.n4711_cascade_\ : std_logic;
signal \tok.n1_adj_724_cascade_\ : std_logic;
signal \tok.n13_adj_725\ : std_logic;
signal \tok.n101_adj_776\ : std_logic;
signal \tok.ram.n4708\ : std_logic;
signal \tok.n1_adj_736\ : std_logic;
signal \tok.n5_adj_737\ : std_logic;
signal \tok.c_stk_r_2\ : std_logic;
signal \tok.table_rd_2\ : std_logic;
signal \tok.n83_adj_721_cascade_\ : std_logic;
signal \tok.n4692\ : std_logic;
signal \tok.ram.n14_adj_631_cascade_\ : std_logic;
signal \tok.n2635\ : std_logic;
signal \tok.n4_adj_795\ : std_logic;
signal \tok.n41_cascade_\ : std_logic;
signal \tok.n884\ : std_logic;
signal \tok.n14_adj_702\ : std_logic;
signal \tok.n15_adj_662\ : std_logic;
signal \tok.n4464\ : std_logic;
signal \tok.n4573\ : std_logic;
signal \tok.n9_adj_645\ : std_logic;
signal \tok.n11\ : std_logic;
signal \tok.n6_cascade_\ : std_logic;
signal \tok.n14\ : std_logic;
signal \tok.n4422_cascade_\ : std_logic;
signal \tok.n11_adj_648\ : std_logic;
signal \tok.n4558\ : std_logic;
signal \tok.n14_adj_650\ : std_logic;
signal \tok.n51_cascade_\ : std_logic;
signal \tok.n4424\ : std_logic;
signal \tok.n48\ : std_logic;
signal \tok.table_rd_12\ : std_logic;
signal \tok.n5_adj_694\ : std_logic;
signal \tok.n10_adj_697\ : std_logic;
signal \tok.n14_adj_695_cascade_\ : std_logic;
signal \tok.A_low_4\ : std_logic;
signal \tok.n18_adj_698\ : std_logic;
signal \tok.n2177\ : std_logic;
signal \tok.n14_adj_825\ : std_logic;
signal \tok.n2177_cascade_\ : std_logic;
signal \tok.n10_adj_646\ : std_logic;
signal \tok.n132\ : std_logic;
signal \tok.table_rd_8\ : std_logic;
signal \tok.n132_cascade_\ : std_logic;
signal \tok.n5\ : std_logic;
signal \tok.n10_adj_652\ : std_logic;
signal \tok.n14_adj_651\ : std_logic;
signal \tok.n109\ : std_logic;
signal \tok.A_low_0\ : std_logic;
signal \tok.n18\ : std_logic;
signal \tok.A_low_6\ : std_logic;
signal \tok.n179\ : std_logic;
signal \tok.n10_adj_675\ : std_logic;
signal \tok.n9\ : std_logic;
signal \tok.n10_adj_675_cascade_\ : std_logic;
signal \tok.n2586\ : std_logic;
signal \tok.T_3\ : std_logic;
signal \tok.n2178\ : std_logic;
signal \tok.n41\ : std_logic;
signal \tok.n4484\ : std_logic;
signal \tok.n40_adj_661\ : std_logic;
signal \tok.n42\ : std_logic;
signal \tok.n4688\ : std_logic;
signal \tok.n10\ : std_logic;
signal \tok.n14_adj_658_cascade_\ : std_logic;
signal \tok.n399\ : std_logic;
signal \tok.table_rd_4\ : std_logic;
signal \tok.c_stk_r_4\ : std_logic;
signal \tok.n83_adj_743\ : std_logic;
signal \tok.c_stk_r_3\ : std_logic;
signal \tok.T_1\ : std_logic;
signal \tok.table_rd_3\ : std_logic;
signal \tok.T_0\ : std_logic;
signal \tok.n83_adj_733_cascade_\ : std_logic;
signal \tok.T_2\ : std_logic;
signal \tok.n4627\ : std_logic;
signal \tok.n883\ : std_logic;
signal \tok.n10_adj_679\ : std_logic;
signal \tok.S_0\ : std_logic;
signal \tok.n2616\ : std_logic;
signal \tok.n15_adj_680\ : std_logic;
signal \tok.n14_adj_658\ : std_logic;
signal \tok.n11_adj_649\ : std_logic;
signal \tok.write_flag\ : std_logic;
signal \tok.T_4\ : std_logic;
signal \tok.T_7\ : std_logic;
signal \tok.T_5\ : std_logic;
signal \tok.T_6\ : std_logic;
signal \tok.n8\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal rx_wire : std_logic;
signal tx_wire : std_logic;
signal reset_wire : std_logic;
signal \tok.vals.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.vals.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.vals.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.vals.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \tok.vals.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.keys.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.keys.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.keys.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.keys.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \tok.keys.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.ram.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.ram.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.ram.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.ram.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \tok.ram.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    rx_wire <= rx;
    tx <= tx_wire;
    reset_wire <= reset;
    \tok.table_rd_15\ <= \tok.vals.mem1_physical_RDATA_wire\(15);
    \tok.table_rd_14\ <= \tok.vals.mem1_physical_RDATA_wire\(14);
    \tok.table_rd_13\ <= \tok.vals.mem1_physical_RDATA_wire\(13);
    \tok.table_rd_12\ <= \tok.vals.mem1_physical_RDATA_wire\(12);
    \tok.table_rd_11\ <= \tok.vals.mem1_physical_RDATA_wire\(11);
    \tok.table_rd_10\ <= \tok.vals.mem1_physical_RDATA_wire\(10);
    \tok.table_rd_9\ <= \tok.vals.mem1_physical_RDATA_wire\(9);
    \tok.table_rd_8\ <= \tok.vals.mem1_physical_RDATA_wire\(8);
    \tok.table_rd_7\ <= \tok.vals.mem1_physical_RDATA_wire\(7);
    \tok.table_rd_6\ <= \tok.vals.mem1_physical_RDATA_wire\(6);
    \tok.table_rd_5\ <= \tok.vals.mem1_physical_RDATA_wire\(5);
    \tok.table_rd_4\ <= \tok.vals.mem1_physical_RDATA_wire\(4);
    \tok.table_rd_3\ <= \tok.vals.mem1_physical_RDATA_wire\(3);
    \tok.table_rd_2\ <= \tok.vals.mem1_physical_RDATA_wire\(2);
    \tok.table_rd_1\ <= \tok.vals.mem1_physical_RDATA_wire\(1);
    \tok.table_rd_0\ <= \tok.vals.mem1_physical_RDATA_wire\(0);
    \tok.vals.mem1_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__18058\&\N__19219\&\N__18127\&\N__18209\&\N__18286\&\N__18352\&\N__18427\&\N__17809\;
    \tok.vals.mem1_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__18055\&\N__19216\&\N__18124\&\N__18206\&\N__18283\&\N__18355\&\N__18424\&\N__17806\;
    \tok.vals.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \tok.vals.mem1_physical_WDATA_wire\ <= \N__10730\&\N__10718\&\N__10703\&\N__11000\&\N__12050\&\N__14888\&\N__10643\&\N__10739\&\N__12014\&\N__17000\&\N__14822\&\N__12005\&\N__13238\&\N__16892\&\N__11993\&\N__17054\;
    \tok.key_rd_15\ <= \tok.keys.mem0_physical_RDATA_wire\(15);
    \tok.key_rd_14\ <= \tok.keys.mem0_physical_RDATA_wire\(14);
    \tok.key_rd_13\ <= \tok.keys.mem0_physical_RDATA_wire\(13);
    \tok.key_rd_12\ <= \tok.keys.mem0_physical_RDATA_wire\(12);
    \tok.key_rd_11\ <= \tok.keys.mem0_physical_RDATA_wire\(11);
    \tok.key_rd_10\ <= \tok.keys.mem0_physical_RDATA_wire\(10);
    \tok.key_rd_9\ <= \tok.keys.mem0_physical_RDATA_wire\(9);
    \tok.key_rd_8\ <= \tok.keys.mem0_physical_RDATA_wire\(8);
    \tok.key_rd_7\ <= \tok.keys.mem0_physical_RDATA_wire\(7);
    \tok.key_rd_6\ <= \tok.keys.mem0_physical_RDATA_wire\(6);
    \tok.key_rd_5\ <= \tok.keys.mem0_physical_RDATA_wire\(5);
    \tok.key_rd_4\ <= \tok.keys.mem0_physical_RDATA_wire\(4);
    \tok.key_rd_3\ <= \tok.keys.mem0_physical_RDATA_wire\(3);
    \tok.key_rd_2\ <= \tok.keys.mem0_physical_RDATA_wire\(2);
    \tok.key_rd_1\ <= \tok.keys.mem0_physical_RDATA_wire\(1);
    \tok.key_rd_0\ <= \tok.keys.mem0_physical_RDATA_wire\(0);
    \tok.keys.mem0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__18068\&\N__19229\&\N__18137\&\N__18221\&\N__18296\&\N__18364\&\N__18437\&\N__17819\;
    \tok.keys.mem0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__18067\&\N__19228\&\N__18136\&\N__18220\&\N__18295\&\N__18365\&\N__18436\&\N__17818\;
    \tok.keys.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \tok.keys.mem0_physical_WDATA_wire\ <= \N__20314\&\N__24004\&\N__20681\&\N__22995\&\N__21436\&\N__21067\&\N__22640\&\N__24839\&\N__19762\&\N__28269\&\N__22400\&\N__27447\&\N__21850\&\N__21988\&\N__24187\&\N__26941\;
    \tok.T_7\ <= \tok.ram.mem2_physical_RDATA_wire\(14);
    \tok.T_6\ <= \tok.ram.mem2_physical_RDATA_wire\(12);
    \tok.T_5\ <= \tok.ram.mem2_physical_RDATA_wire\(10);
    \tok.T_4\ <= \tok.ram.mem2_physical_RDATA_wire\(8);
    \tok.T_3\ <= \tok.ram.mem2_physical_RDATA_wire\(6);
    \tok.T_2\ <= \tok.ram.mem2_physical_RDATA_wire\(4);
    \tok.T_1\ <= \tok.ram.mem2_physical_RDATA_wire\(2);
    \tok.T_0\ <= \tok.ram.mem2_physical_RDATA_wire\(0);
    \tok.ram.mem2_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__16844\&\N__18548\&\N__23663\&\N__23447\&\N__23534\&\N__23639\&\N__16745\&\N__18692\;
    \tok.ram.mem2_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__19690\&\N__21322\&\N__19952\&\N__24395\&\N__21551\&\N__20068\&\N__20171\&\N__29575\;
    \tok.ram.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \tok.ram.mem2_physical_WDATA_wire\ <= '0'&\N__19824\&'0'&\N__28268\&'0'&\N__22401\&'0'&\N__27452\&'0'&\N__21845\&'0'&\N__21985\&'0'&\N__24181\&'0'&\N__26934\;

    \tok.vals.mem1_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \tok.vals.mem1_physical_RDATA_wire\,
            RADDR => \tok.vals.mem1_physical_RADDR_wire\,
            WADDR => \tok.vals.mem1_physical_WADDR_wire\,
            MASK => \tok.vals.mem1_physical_MASK_wire\,
            WDATA => \tok.vals.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__26234\,
            RE => \N__21681\,
            WCLKE => 'H',
            WCLK => \N__26233\,
            WE => \N__14846\
        );

    \tok.keys.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \tok.keys.mem0_physical_RDATA_wire\,
            RADDR => \tok.keys.mem0_physical_RADDR_wire\,
            WADDR => \tok.keys.mem0_physical_WADDR_wire\,
            MASK => \tok.keys.mem0_physical_MASK_wire\,
            WDATA => \tok.keys.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__26221\,
            RE => \N__21698\,
            WCLKE => 'H',
            WCLK => \N__26222\,
            WE => \N__14845\
        );

    \tok.ram.mem2_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000001000000010000000101010000000000010100000100000001000000000000000100000001000000010100010101000001010000010000000100000000000000010000000100000001010001010000000101000001000000010000000000000001000000010000000101000100010000010100000100",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \tok.ram.mem2_physical_RDATA_wire\,
            RADDR => \tok.ram.mem2_physical_RADDR_wire\,
            WADDR => \tok.ram.mem2_physical_WADDR_wire\,
            MASK => \tok.ram.mem2_physical_MASK_wire\,
            WDATA => \tok.ram.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__26258\,
            RE => \N__21699\,
            WCLKE => 'H',
            WCLK => \N__26259\,
            WE => \N__29101\
        );

    \rx_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30609\,
            DIN => \N__30608\,
            DOUT => \N__30607\,
            PACKAGEPIN => rx_wire
        );

    \rx_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30609\,
            PADOUT => \N__30608\,
            PADIN => \N__30607\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => rx_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \tx_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30600\,
            DIN => \N__30599\,
            DOUT => \N__30598\,
            PACKAGEPIN => tx_wire
        );

    \tx_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30600\,
            PADOUT => \N__30599\,
            PADIN => \N__30598\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13289\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \reset_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30591\,
            DIN => \N__30590\,
            DOUT => \N__30589\,
            PACKAGEPIN => reset_wire
        );

    \reset_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30591\,
            PADOUT => \N__30590\,
            PADIN => \N__30589\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => reset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__7643\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30568\
        );

    \I__7642\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30565\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__30568\,
            I => \N__30562\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__30565\,
            I => \N__30559\
        );

    \I__7639\ : Span4Mux_v
    port map (
            O => \N__30562\,
            I => \N__30556\
        );

    \I__7638\ : Span4Mux_v
    port map (
            O => \N__30559\,
            I => \N__30553\
        );

    \I__7637\ : Span4Mux_h
    port map (
            O => \N__30556\,
            I => \N__30550\
        );

    \I__7636\ : Sp12to4
    port map (
            O => \N__30553\,
            I => \N__30545\
        );

    \I__7635\ : Sp12to4
    port map (
            O => \N__30550\,
            I => \N__30545\
        );

    \I__7634\ : Span12Mux_s10_h
    port map (
            O => \N__30545\,
            I => \N__30542\
        );

    \I__7633\ : Odrv12
    port map (
            O => \N__30542\,
            I => \tok.table_rd_4\
        );

    \I__7632\ : CascadeMux
    port map (
            O => \N__30539\,
            I => \N__30532\
        );

    \I__7631\ : InMux
    port map (
            O => \N__30538\,
            I => \N__30529\
        );

    \I__7630\ : InMux
    port map (
            O => \N__30537\,
            I => \N__30526\
        );

    \I__7629\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30519\
        );

    \I__7628\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30519\
        );

    \I__7627\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30519\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__30529\,
            I => \N__30516\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__30526\,
            I => \N__30513\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__30519\,
            I => \N__30510\
        );

    \I__7623\ : Span4Mux_h
    port map (
            O => \N__30516\,
            I => \N__30505\
        );

    \I__7622\ : Span4Mux_v
    port map (
            O => \N__30513\,
            I => \N__30505\
        );

    \I__7621\ : Odrv4
    port map (
            O => \N__30510\,
            I => \tok.c_stk_r_4\
        );

    \I__7620\ : Odrv4
    port map (
            O => \N__30505\,
            I => \tok.c_stk_r_4\
        );

    \I__7619\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30497\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__30497\,
            I => \tok.n83_adj_743\
        );

    \I__7617\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30490\
        );

    \I__7616\ : CascadeMux
    port map (
            O => \N__30493\,
            I => \N__30484\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__30490\,
            I => \N__30481\
        );

    \I__7614\ : CascadeMux
    port map (
            O => \N__30489\,
            I => \N__30478\
        );

    \I__7613\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30475\
        );

    \I__7612\ : InMux
    port map (
            O => \N__30487\,
            I => \N__30472\
        );

    \I__7611\ : InMux
    port map (
            O => \N__30484\,
            I => \N__30469\
        );

    \I__7610\ : Span4Mux_v
    port map (
            O => \N__30481\,
            I => \N__30466\
        );

    \I__7609\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30463\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__30475\,
            I => \tok.c_stk_r_3\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__30472\,
            I => \tok.c_stk_r_3\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__30469\,
            I => \tok.c_stk_r_3\
        );

    \I__7605\ : Odrv4
    port map (
            O => \N__30466\,
            I => \tok.c_stk_r_3\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__30463\,
            I => \tok.c_stk_r_3\
        );

    \I__7603\ : CascadeMux
    port map (
            O => \N__30452\,
            I => \N__30449\
        );

    \I__7602\ : InMux
    port map (
            O => \N__30449\,
            I => \N__30438\
        );

    \I__7601\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30433\
        );

    \I__7600\ : InMux
    port map (
            O => \N__30447\,
            I => \N__30433\
        );

    \I__7599\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30424\
        );

    \I__7598\ : InMux
    port map (
            O => \N__30445\,
            I => \N__30424\
        );

    \I__7597\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30424\
        );

    \I__7596\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30424\
        );

    \I__7595\ : CascadeMux
    port map (
            O => \N__30442\,
            I => \N__30420\
        );

    \I__7594\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30413\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__30438\,
            I => \N__30405\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__30433\,
            I => \N__30405\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30402\
        );

    \I__7590\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30395\
        );

    \I__7589\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30395\
        );

    \I__7588\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30395\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__30418\,
            I => \N__30386\
        );

    \I__7586\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30375\
        );

    \I__7585\ : InMux
    port map (
            O => \N__30416\,
            I => \N__30375\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__30413\,
            I => \N__30372\
        );

    \I__7583\ : InMux
    port map (
            O => \N__30412\,
            I => \N__30369\
        );

    \I__7582\ : InMux
    port map (
            O => \N__30411\,
            I => \N__30366\
        );

    \I__7581\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30363\
        );

    \I__7580\ : Span4Mux_h
    port map (
            O => \N__30405\,
            I => \N__30356\
        );

    \I__7579\ : Span4Mux_s3_v
    port map (
            O => \N__30402\,
            I => \N__30356\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__30395\,
            I => \N__30356\
        );

    \I__7577\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30353\
        );

    \I__7576\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30349\
        );

    \I__7575\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30346\
        );

    \I__7574\ : InMux
    port map (
            O => \N__30391\,
            I => \N__30340\
        );

    \I__7573\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30340\
        );

    \I__7572\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30333\
        );

    \I__7571\ : InMux
    port map (
            O => \N__30386\,
            I => \N__30333\
        );

    \I__7570\ : InMux
    port map (
            O => \N__30385\,
            I => \N__30333\
        );

    \I__7569\ : InMux
    port map (
            O => \N__30384\,
            I => \N__30324\
        );

    \I__7568\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30324\
        );

    \I__7567\ : InMux
    port map (
            O => \N__30382\,
            I => \N__30324\
        );

    \I__7566\ : InMux
    port map (
            O => \N__30381\,
            I => \N__30324\
        );

    \I__7565\ : InMux
    port map (
            O => \N__30380\,
            I => \N__30319\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__30375\,
            I => \N__30316\
        );

    \I__7563\ : Span4Mux_v
    port map (
            O => \N__30372\,
            I => \N__30313\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__30369\,
            I => \N__30310\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__30366\,
            I => \N__30301\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__30363\,
            I => \N__30301\
        );

    \I__7559\ : Span4Mux_h
    port map (
            O => \N__30356\,
            I => \N__30301\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30301\
        );

    \I__7557\ : InMux
    port map (
            O => \N__30352\,
            I => \N__30298\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__30349\,
            I => \N__30295\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__30346\,
            I => \N__30292\
        );

    \I__7554\ : CascadeMux
    port map (
            O => \N__30345\,
            I => \N__30283\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__30340\,
            I => \N__30276\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__30333\,
            I => \N__30271\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__30324\,
            I => \N__30271\
        );

    \I__7550\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30266\
        );

    \I__7549\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30266\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__30319\,
            I => \N__30263\
        );

    \I__7547\ : Span4Mux_v
    port map (
            O => \N__30316\,
            I => \N__30260\
        );

    \I__7546\ : Span4Mux_h
    port map (
            O => \N__30313\,
            I => \N__30253\
        );

    \I__7545\ : Span4Mux_v
    port map (
            O => \N__30310\,
            I => \N__30253\
        );

    \I__7544\ : Span4Mux_v
    port map (
            O => \N__30301\,
            I => \N__30253\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__30298\,
            I => \N__30250\
        );

    \I__7542\ : Span4Mux_v
    port map (
            O => \N__30295\,
            I => \N__30245\
        );

    \I__7541\ : Span4Mux_s2_h
    port map (
            O => \N__30292\,
            I => \N__30245\
        );

    \I__7540\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30238\
        );

    \I__7539\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30238\
        );

    \I__7538\ : InMux
    port map (
            O => \N__30289\,
            I => \N__30238\
        );

    \I__7537\ : InMux
    port map (
            O => \N__30288\,
            I => \N__30231\
        );

    \I__7536\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30231\
        );

    \I__7535\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30231\
        );

    \I__7534\ : InMux
    port map (
            O => \N__30283\,
            I => \N__30220\
        );

    \I__7533\ : InMux
    port map (
            O => \N__30282\,
            I => \N__30220\
        );

    \I__7532\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30220\
        );

    \I__7531\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30220\
        );

    \I__7530\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30220\
        );

    \I__7529\ : Span4Mux_h
    port map (
            O => \N__30276\,
            I => \N__30213\
        );

    \I__7528\ : Span4Mux_s3_h
    port map (
            O => \N__30271\,
            I => \N__30213\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__30266\,
            I => \N__30213\
        );

    \I__7526\ : Odrv4
    port map (
            O => \N__30263\,
            I => \tok.T_1\
        );

    \I__7525\ : Odrv4
    port map (
            O => \N__30260\,
            I => \tok.T_1\
        );

    \I__7524\ : Odrv4
    port map (
            O => \N__30253\,
            I => \tok.T_1\
        );

    \I__7523\ : Odrv4
    port map (
            O => \N__30250\,
            I => \tok.T_1\
        );

    \I__7522\ : Odrv4
    port map (
            O => \N__30245\,
            I => \tok.T_1\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__30238\,
            I => \tok.T_1\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__30231\,
            I => \tok.T_1\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__30220\,
            I => \tok.T_1\
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__30213\,
            I => \tok.T_1\
        );

    \I__7517\ : CascadeMux
    port map (
            O => \N__30194\,
            I => \N__30191\
        );

    \I__7516\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30188\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__30188\,
            I => \N__30185\
        );

    \I__7514\ : Span4Mux_v
    port map (
            O => \N__30185\,
            I => \N__30181\
        );

    \I__7513\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30178\
        );

    \I__7512\ : Span4Mux_h
    port map (
            O => \N__30181\,
            I => \N__30175\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__30178\,
            I => \N__30172\
        );

    \I__7510\ : Span4Mux_h
    port map (
            O => \N__30175\,
            I => \N__30169\
        );

    \I__7509\ : Odrv12
    port map (
            O => \N__30172\,
            I => \tok.table_rd_3\
        );

    \I__7508\ : Odrv4
    port map (
            O => \N__30169\,
            I => \tok.table_rd_3\
        );

    \I__7507\ : InMux
    port map (
            O => \N__30164\,
            I => \N__30138\
        );

    \I__7506\ : InMux
    port map (
            O => \N__30163\,
            I => \N__30138\
        );

    \I__7505\ : InMux
    port map (
            O => \N__30162\,
            I => \N__30138\
        );

    \I__7504\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30131\
        );

    \I__7503\ : InMux
    port map (
            O => \N__30160\,
            I => \N__30128\
        );

    \I__7502\ : InMux
    port map (
            O => \N__30159\,
            I => \N__30121\
        );

    \I__7501\ : InMux
    port map (
            O => \N__30158\,
            I => \N__30121\
        );

    \I__7500\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30121\
        );

    \I__7499\ : InMux
    port map (
            O => \N__30156\,
            I => \N__30114\
        );

    \I__7498\ : InMux
    port map (
            O => \N__30155\,
            I => \N__30114\
        );

    \I__7497\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30114\
        );

    \I__7496\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30099\
        );

    \I__7495\ : InMux
    port map (
            O => \N__30152\,
            I => \N__30094\
        );

    \I__7494\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30094\
        );

    \I__7493\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30089\
        );

    \I__7492\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30089\
        );

    \I__7491\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30086\
        );

    \I__7490\ : InMux
    port map (
            O => \N__30147\,
            I => \N__30083\
        );

    \I__7489\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30078\
        );

    \I__7488\ : InMux
    port map (
            O => \N__30145\,
            I => \N__30078\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__30138\,
            I => \N__30075\
        );

    \I__7486\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30072\
        );

    \I__7485\ : InMux
    port map (
            O => \N__30136\,
            I => \N__30069\
        );

    \I__7484\ : InMux
    port map (
            O => \N__30135\,
            I => \N__30066\
        );

    \I__7483\ : InMux
    port map (
            O => \N__30134\,
            I => \N__30063\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__30131\,
            I => \N__30056\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__30128\,
            I => \N__30056\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__30121\,
            I => \N__30056\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__30114\,
            I => \N__30053\
        );

    \I__7478\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30050\
        );

    \I__7477\ : InMux
    port map (
            O => \N__30112\,
            I => \N__30045\
        );

    \I__7476\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30045\
        );

    \I__7475\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30041\
        );

    \I__7474\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30037\
        );

    \I__7473\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30030\
        );

    \I__7472\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30030\
        );

    \I__7471\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30030\
        );

    \I__7470\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30021\
        );

    \I__7469\ : InMux
    port map (
            O => \N__30104\,
            I => \N__30021\
        );

    \I__7468\ : InMux
    port map (
            O => \N__30103\,
            I => \N__30021\
        );

    \I__7467\ : InMux
    port map (
            O => \N__30102\,
            I => \N__30021\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__30099\,
            I => \N__30015\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__30094\,
            I => \N__30015\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__30089\,
            I => \N__30010\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__30086\,
            I => \N__30010\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__30083\,
            I => \N__30001\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__30078\,
            I => \N__30001\
        );

    \I__7460\ : Span4Mux_v
    port map (
            O => \N__30075\,
            I => \N__30001\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__30072\,
            I => \N__30001\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__30069\,
            I => \N__29998\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__30066\,
            I => \N__29995\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__30063\,
            I => \N__29988\
        );

    \I__7455\ : Span4Mux_s3_v
    port map (
            O => \N__30056\,
            I => \N__29988\
        );

    \I__7454\ : Span4Mux_h
    port map (
            O => \N__30053\,
            I => \N__29988\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__30050\,
            I => \N__29985\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__30045\,
            I => \N__29982\
        );

    \I__7451\ : InMux
    port map (
            O => \N__30044\,
            I => \N__29979\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__30041\,
            I => \N__29976\
        );

    \I__7449\ : CascadeMux
    port map (
            O => \N__30040\,
            I => \N__29970\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__30037\,
            I => \N__29959\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__30030\,
            I => \N__29954\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__30021\,
            I => \N__29954\
        );

    \I__7445\ : InMux
    port map (
            O => \N__30020\,
            I => \N__29951\
        );

    \I__7444\ : Span4Mux_s3_h
    port map (
            O => \N__30015\,
            I => \N__29944\
        );

    \I__7443\ : Span4Mux_h
    port map (
            O => \N__30010\,
            I => \N__29944\
        );

    \I__7442\ : Span4Mux_h
    port map (
            O => \N__30001\,
            I => \N__29944\
        );

    \I__7441\ : Span4Mux_v
    port map (
            O => \N__29998\,
            I => \N__29931\
        );

    \I__7440\ : Span4Mux_h
    port map (
            O => \N__29995\,
            I => \N__29931\
        );

    \I__7439\ : Span4Mux_v
    port map (
            O => \N__29988\,
            I => \N__29931\
        );

    \I__7438\ : Span4Mux_v
    port map (
            O => \N__29985\,
            I => \N__29931\
        );

    \I__7437\ : Span4Mux_v
    port map (
            O => \N__29982\,
            I => \N__29931\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__29979\,
            I => \N__29931\
        );

    \I__7435\ : Span4Mux_s2_h
    port map (
            O => \N__29976\,
            I => \N__29928\
        );

    \I__7434\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29921\
        );

    \I__7433\ : InMux
    port map (
            O => \N__29974\,
            I => \N__29921\
        );

    \I__7432\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29921\
        );

    \I__7431\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29914\
        );

    \I__7430\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29914\
        );

    \I__7429\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29914\
        );

    \I__7428\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29911\
        );

    \I__7427\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29900\
        );

    \I__7426\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29900\
        );

    \I__7425\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29900\
        );

    \I__7424\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29900\
        );

    \I__7423\ : InMux
    port map (
            O => \N__29962\,
            I => \N__29900\
        );

    \I__7422\ : Span4Mux_s3_h
    port map (
            O => \N__29959\,
            I => \N__29893\
        );

    \I__7421\ : Span4Mux_s3_h
    port map (
            O => \N__29954\,
            I => \N__29893\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__29951\,
            I => \N__29893\
        );

    \I__7419\ : Odrv4
    port map (
            O => \N__29944\,
            I => \tok.T_0\
        );

    \I__7418\ : Odrv4
    port map (
            O => \N__29931\,
            I => \tok.T_0\
        );

    \I__7417\ : Odrv4
    port map (
            O => \N__29928\,
            I => \tok.T_0\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__29921\,
            I => \tok.T_0\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__29914\,
            I => \tok.T_0\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__29911\,
            I => \tok.T_0\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__29900\,
            I => \tok.T_0\
        );

    \I__7412\ : Odrv4
    port map (
            O => \N__29893\,
            I => \tok.T_0\
        );

    \I__7411\ : CascadeMux
    port map (
            O => \N__29876\,
            I => \tok.n83_adj_733_cascade_\
        );

    \I__7410\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29844\
        );

    \I__7409\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29837\
        );

    \I__7408\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29837\
        );

    \I__7407\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29837\
        );

    \I__7406\ : InMux
    port map (
            O => \N__29869\,
            I => \N__29832\
        );

    \I__7405\ : InMux
    port map (
            O => \N__29868\,
            I => \N__29832\
        );

    \I__7404\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29825\
        );

    \I__7403\ : InMux
    port map (
            O => \N__29866\,
            I => \N__29825\
        );

    \I__7402\ : InMux
    port map (
            O => \N__29865\,
            I => \N__29825\
        );

    \I__7401\ : CascadeMux
    port map (
            O => \N__29864\,
            I => \N__29821\
        );

    \I__7400\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29814\
        );

    \I__7399\ : InMux
    port map (
            O => \N__29862\,
            I => \N__29814\
        );

    \I__7398\ : InMux
    port map (
            O => \N__29861\,
            I => \N__29811\
        );

    \I__7397\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29808\
        );

    \I__7396\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29803\
        );

    \I__7395\ : InMux
    port map (
            O => \N__29858\,
            I => \N__29803\
        );

    \I__7394\ : InMux
    port map (
            O => \N__29857\,
            I => \N__29794\
        );

    \I__7393\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29794\
        );

    \I__7392\ : InMux
    port map (
            O => \N__29855\,
            I => \N__29791\
        );

    \I__7391\ : InMux
    port map (
            O => \N__29854\,
            I => \N__29786\
        );

    \I__7390\ : InMux
    port map (
            O => \N__29853\,
            I => \N__29786\
        );

    \I__7389\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29783\
        );

    \I__7388\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29779\
        );

    \I__7387\ : InMux
    port map (
            O => \N__29850\,
            I => \N__29774\
        );

    \I__7386\ : InMux
    port map (
            O => \N__29849\,
            I => \N__29774\
        );

    \I__7385\ : InMux
    port map (
            O => \N__29848\,
            I => \N__29771\
        );

    \I__7384\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29768\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__29844\,
            I => \N__29765\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__29837\,
            I => \N__29762\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29757\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__29825\,
            I => \N__29757\
        );

    \I__7379\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29754\
        );

    \I__7378\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29747\
        );

    \I__7377\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29747\
        );

    \I__7376\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29747\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__29814\,
            I => \N__29738\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__29811\,
            I => \N__29738\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__29808\,
            I => \N__29738\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__29803\,
            I => \N__29738\
        );

    \I__7371\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29733\
        );

    \I__7370\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29733\
        );

    \I__7369\ : InMux
    port map (
            O => \N__29800\,
            I => \N__29728\
        );

    \I__7368\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29728\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__29794\,
            I => \N__29725\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__29791\,
            I => \N__29718\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__29786\,
            I => \N__29718\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__29783\,
            I => \N__29718\
        );

    \I__7363\ : InMux
    port map (
            O => \N__29782\,
            I => \N__29715\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__29779\,
            I => \N__29712\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__29774\,
            I => \N__29709\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__29771\,
            I => \N__29706\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__29768\,
            I => \N__29697\
        );

    \I__7358\ : Span4Mux_h
    port map (
            O => \N__29765\,
            I => \N__29697\
        );

    \I__7357\ : Span4Mux_s3_v
    port map (
            O => \N__29762\,
            I => \N__29697\
        );

    \I__7356\ : Span4Mux_h
    port map (
            O => \N__29757\,
            I => \N__29697\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__29754\,
            I => \N__29692\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__29747\,
            I => \N__29692\
        );

    \I__7353\ : Span4Mux_v
    port map (
            O => \N__29738\,
            I => \N__29689\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__29733\,
            I => \N__29686\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__29728\,
            I => \N__29671\
        );

    \I__7350\ : Span4Mux_v
    port map (
            O => \N__29725\,
            I => \N__29666\
        );

    \I__7349\ : Span4Mux_h
    port map (
            O => \N__29718\,
            I => \N__29666\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29663\
        );

    \I__7347\ : Span4Mux_v
    port map (
            O => \N__29712\,
            I => \N__29648\
        );

    \I__7346\ : Span4Mux_h
    port map (
            O => \N__29709\,
            I => \N__29648\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__29706\,
            I => \N__29648\
        );

    \I__7344\ : Span4Mux_v
    port map (
            O => \N__29697\,
            I => \N__29648\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__29692\,
            I => \N__29648\
        );

    \I__7342\ : Span4Mux_s0_h
    port map (
            O => \N__29689\,
            I => \N__29648\
        );

    \I__7341\ : Span4Mux_v
    port map (
            O => \N__29686\,
            I => \N__29648\
        );

    \I__7340\ : InMux
    port map (
            O => \N__29685\,
            I => \N__29643\
        );

    \I__7339\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29643\
        );

    \I__7338\ : InMux
    port map (
            O => \N__29683\,
            I => \N__29636\
        );

    \I__7337\ : InMux
    port map (
            O => \N__29682\,
            I => \N__29636\
        );

    \I__7336\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29636\
        );

    \I__7335\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29621\
        );

    \I__7334\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29621\
        );

    \I__7333\ : InMux
    port map (
            O => \N__29678\,
            I => \N__29621\
        );

    \I__7332\ : InMux
    port map (
            O => \N__29677\,
            I => \N__29621\
        );

    \I__7331\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29621\
        );

    \I__7330\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29621\
        );

    \I__7329\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29621\
        );

    \I__7328\ : Odrv4
    port map (
            O => \N__29671\,
            I => \tok.T_2\
        );

    \I__7327\ : Odrv4
    port map (
            O => \N__29666\,
            I => \tok.T_2\
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__29663\,
            I => \tok.T_2\
        );

    \I__7325\ : Odrv4
    port map (
            O => \N__29648\,
            I => \tok.T_2\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__29643\,
            I => \tok.T_2\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__29636\,
            I => \tok.T_2\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__29621\,
            I => \tok.T_2\
        );

    \I__7321\ : CascadeMux
    port map (
            O => \N__29606\,
            I => \N__29603\
        );

    \I__7320\ : InMux
    port map (
            O => \N__29603\,
            I => \N__29600\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__29600\,
            I => \tok.n4627\
        );

    \I__7318\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29594\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__29594\,
            I => \tok.n883\
        );

    \I__7316\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29588\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__7314\ : Sp12to4
    port map (
            O => \N__29585\,
            I => \N__29582\
        );

    \I__7313\ : Span12Mux_s7_v
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__7312\ : Odrv12
    port map (
            O => \N__29579\,
            I => \tok.n10_adj_679\
        );

    \I__7311\ : CascadeMux
    port map (
            O => \N__29576\,
            I => \N__29568\
        );

    \I__7310\ : CascadeMux
    port map (
            O => \N__29575\,
            I => \N__29565\
        );

    \I__7309\ : CascadeMux
    port map (
            O => \N__29574\,
            I => \N__29562\
        );

    \I__7308\ : InMux
    port map (
            O => \N__29573\,
            I => \N__29559\
        );

    \I__7307\ : InMux
    port map (
            O => \N__29572\,
            I => \N__29556\
        );

    \I__7306\ : CascadeMux
    port map (
            O => \N__29571\,
            I => \N__29553\
        );

    \I__7305\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29550\
        );

    \I__7304\ : InMux
    port map (
            O => \N__29565\,
            I => \N__29545\
        );

    \I__7303\ : InMux
    port map (
            O => \N__29562\,
            I => \N__29542\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__29559\,
            I => \N__29539\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__29556\,
            I => \N__29536\
        );

    \I__7300\ : InMux
    port map (
            O => \N__29553\,
            I => \N__29533\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__29550\,
            I => \N__29530\
        );

    \I__7298\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29527\
        );

    \I__7297\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29524\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__29545\,
            I => \N__29519\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__29542\,
            I => \N__29519\
        );

    \I__7294\ : Span4Mux_v
    port map (
            O => \N__29539\,
            I => \N__29515\
        );

    \I__7293\ : Span4Mux_v
    port map (
            O => \N__29536\,
            I => \N__29512\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__29533\,
            I => \N__29509\
        );

    \I__7291\ : Span4Mux_h
    port map (
            O => \N__29530\,
            I => \N__29506\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__29527\,
            I => \N__29501\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29501\
        );

    \I__7288\ : Span4Mux_v
    port map (
            O => \N__29519\,
            I => \N__29498\
        );

    \I__7287\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29495\
        );

    \I__7286\ : Span4Mux_h
    port map (
            O => \N__29515\,
            I => \N__29492\
        );

    \I__7285\ : Span4Mux_h
    port map (
            O => \N__29512\,
            I => \N__29487\
        );

    \I__7284\ : Span4Mux_v
    port map (
            O => \N__29509\,
            I => \N__29487\
        );

    \I__7283\ : Span4Mux_v
    port map (
            O => \N__29506\,
            I => \N__29480\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__29501\,
            I => \N__29480\
        );

    \I__7281\ : Span4Mux_h
    port map (
            O => \N__29498\,
            I => \N__29480\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29473\
        );

    \I__7279\ : Span4Mux_h
    port map (
            O => \N__29492\,
            I => \N__29473\
        );

    \I__7278\ : Span4Mux_v
    port map (
            O => \N__29487\,
            I => \N__29473\
        );

    \I__7277\ : Span4Mux_h
    port map (
            O => \N__29480\,
            I => \N__29470\
        );

    \I__7276\ : Odrv4
    port map (
            O => \N__29473\,
            I => \tok.S_0\
        );

    \I__7275\ : Odrv4
    port map (
            O => \N__29470\,
            I => \tok.S_0\
        );

    \I__7274\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29462\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__29462\,
            I => \N__29454\
        );

    \I__7272\ : InMux
    port map (
            O => \N__29461\,
            I => \N__29451\
        );

    \I__7271\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29446\
        );

    \I__7270\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29446\
        );

    \I__7269\ : InMux
    port map (
            O => \N__29458\,
            I => \N__29441\
        );

    \I__7268\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29437\
        );

    \I__7267\ : Span4Mux_h
    port map (
            O => \N__29454\,
            I => \N__29431\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__29451\,
            I => \N__29431\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__29446\,
            I => \N__29428\
        );

    \I__7264\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29425\
        );

    \I__7263\ : InMux
    port map (
            O => \N__29444\,
            I => \N__29422\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__29441\,
            I => \N__29418\
        );

    \I__7261\ : InMux
    port map (
            O => \N__29440\,
            I => \N__29415\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29412\
        );

    \I__7259\ : InMux
    port map (
            O => \N__29436\,
            I => \N__29408\
        );

    \I__7258\ : Span4Mux_v
    port map (
            O => \N__29431\,
            I => \N__29405\
        );

    \I__7257\ : Span4Mux_h
    port map (
            O => \N__29428\,
            I => \N__29398\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__29425\,
            I => \N__29398\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__29422\,
            I => \N__29398\
        );

    \I__7254\ : InMux
    port map (
            O => \N__29421\,
            I => \N__29395\
        );

    \I__7253\ : Span4Mux_h
    port map (
            O => \N__29418\,
            I => \N__29387\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__29415\,
            I => \N__29387\
        );

    \I__7251\ : Span4Mux_s0_h
    port map (
            O => \N__29412\,
            I => \N__29384\
        );

    \I__7250\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29381\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__29408\,
            I => \N__29378\
        );

    \I__7248\ : Span4Mux_h
    port map (
            O => \N__29405\,
            I => \N__29371\
        );

    \I__7247\ : Span4Mux_h
    port map (
            O => \N__29398\,
            I => \N__29371\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__29395\,
            I => \N__29371\
        );

    \I__7245\ : InMux
    port map (
            O => \N__29394\,
            I => \N__29368\
        );

    \I__7244\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29363\
        );

    \I__7243\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29363\
        );

    \I__7242\ : Span4Mux_h
    port map (
            O => \N__29387\,
            I => \N__29358\
        );

    \I__7241\ : Span4Mux_h
    port map (
            O => \N__29384\,
            I => \N__29358\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__29381\,
            I => \N__29353\
        );

    \I__7239\ : Span12Mux_s5_v
    port map (
            O => \N__29378\,
            I => \N__29353\
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__29371\,
            I => \tok.n2616\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__29368\,
            I => \tok.n2616\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__29363\,
            I => \tok.n2616\
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__29358\,
            I => \tok.n2616\
        );

    \I__7234\ : Odrv12
    port map (
            O => \N__29353\,
            I => \tok.n2616\
        );

    \I__7233\ : InMux
    port map (
            O => \N__29342\,
            I => \N__29339\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__29339\,
            I => \N__29336\
        );

    \I__7231\ : Span4Mux_h
    port map (
            O => \N__29336\,
            I => \N__29333\
        );

    \I__7230\ : Span4Mux_h
    port map (
            O => \N__29333\,
            I => \N__29330\
        );

    \I__7229\ : Odrv4
    port map (
            O => \N__29330\,
            I => \tok.n15_adj_680\
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__29327\,
            I => \N__29323\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__29326\,
            I => \N__29318\
        );

    \I__7226\ : InMux
    port map (
            O => \N__29323\,
            I => \N__29306\
        );

    \I__7225\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29306\
        );

    \I__7224\ : InMux
    port map (
            O => \N__29321\,
            I => \N__29306\
        );

    \I__7223\ : InMux
    port map (
            O => \N__29318\,
            I => \N__29306\
        );

    \I__7222\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29306\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__29306\,
            I => \N__29301\
        );

    \I__7220\ : InMux
    port map (
            O => \N__29305\,
            I => \N__29298\
        );

    \I__7219\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29295\
        );

    \I__7218\ : Span4Mux_h
    port map (
            O => \N__29301\,
            I => \N__29286\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__29298\,
            I => \N__29286\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__29295\,
            I => \N__29275\
        );

    \I__7215\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29268\
        );

    \I__7214\ : InMux
    port map (
            O => \N__29293\,
            I => \N__29268\
        );

    \I__7213\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29268\
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__29291\,
            I => \N__29262\
        );

    \I__7211\ : Span4Mux_v
    port map (
            O => \N__29286\,
            I => \N__29255\
        );

    \I__7210\ : InMux
    port map (
            O => \N__29285\,
            I => \N__29252\
        );

    \I__7209\ : CascadeMux
    port map (
            O => \N__29284\,
            I => \N__29248\
        );

    \I__7208\ : InMux
    port map (
            O => \N__29283\,
            I => \N__29236\
        );

    \I__7207\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29236\
        );

    \I__7206\ : InMux
    port map (
            O => \N__29281\,
            I => \N__29236\
        );

    \I__7205\ : InMux
    port map (
            O => \N__29280\,
            I => \N__29236\
        );

    \I__7204\ : InMux
    port map (
            O => \N__29279\,
            I => \N__29236\
        );

    \I__7203\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29233\
        );

    \I__7202\ : Span4Mux_h
    port map (
            O => \N__29275\,
            I => \N__29230\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__29268\,
            I => \N__29227\
        );

    \I__7200\ : CascadeMux
    port map (
            O => \N__29267\,
            I => \N__29223\
        );

    \I__7199\ : CascadeMux
    port map (
            O => \N__29266\,
            I => \N__29218\
        );

    \I__7198\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29209\
        );

    \I__7197\ : InMux
    port map (
            O => \N__29262\,
            I => \N__29209\
        );

    \I__7196\ : InMux
    port map (
            O => \N__29261\,
            I => \N__29209\
        );

    \I__7195\ : InMux
    port map (
            O => \N__29260\,
            I => \N__29209\
        );

    \I__7194\ : InMux
    port map (
            O => \N__29259\,
            I => \N__29204\
        );

    \I__7193\ : InMux
    port map (
            O => \N__29258\,
            I => \N__29204\
        );

    \I__7192\ : Span4Mux_h
    port map (
            O => \N__29255\,
            I => \N__29199\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__29252\,
            I => \N__29199\
        );

    \I__7190\ : InMux
    port map (
            O => \N__29251\,
            I => \N__29192\
        );

    \I__7189\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29192\
        );

    \I__7188\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29192\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__29236\,
            I => \N__29189\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__29233\,
            I => \N__29186\
        );

    \I__7185\ : Span4Mux_h
    port map (
            O => \N__29230\,
            I => \N__29181\
        );

    \I__7184\ : Span4Mux_h
    port map (
            O => \N__29227\,
            I => \N__29181\
        );

    \I__7183\ : InMux
    port map (
            O => \N__29226\,
            I => \N__29170\
        );

    \I__7182\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29170\
        );

    \I__7181\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29170\
        );

    \I__7180\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29170\
        );

    \I__7179\ : InMux
    port map (
            O => \N__29218\,
            I => \N__29170\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__29209\,
            I => \N__29165\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__29204\,
            I => \N__29165\
        );

    \I__7176\ : Span4Mux_h
    port map (
            O => \N__29199\,
            I => \N__29162\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__29192\,
            I => \N__29155\
        );

    \I__7174\ : Span4Mux_h
    port map (
            O => \N__29189\,
            I => \N__29155\
        );

    \I__7173\ : Span4Mux_v
    port map (
            O => \N__29186\,
            I => \N__29155\
        );

    \I__7172\ : Sp12to4
    port map (
            O => \N__29181\,
            I => \N__29150\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__29170\,
            I => \N__29150\
        );

    \I__7170\ : Span12Mux_h
    port map (
            O => \N__29165\,
            I => \N__29146\
        );

    \I__7169\ : Span4Mux_v
    port map (
            O => \N__29162\,
            I => \N__29143\
        );

    \I__7168\ : Sp12to4
    port map (
            O => \N__29155\,
            I => \N__29138\
        );

    \I__7167\ : Span12Mux_s7_v
    port map (
            O => \N__29150\,
            I => \N__29138\
        );

    \I__7166\ : InMux
    port map (
            O => \N__29149\,
            I => \N__29135\
        );

    \I__7165\ : Odrv12
    port map (
            O => \N__29146\,
            I => \tok.n14_adj_658\
        );

    \I__7164\ : Odrv4
    port map (
            O => \N__29143\,
            I => \tok.n14_adj_658\
        );

    \I__7163\ : Odrv12
    port map (
            O => \N__29138\,
            I => \tok.n14_adj_658\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__29135\,
            I => \tok.n14_adj_658\
        );

    \I__7161\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29123\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__29123\,
            I => \N__29118\
        );

    \I__7159\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29113\
        );

    \I__7158\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29113\
        );

    \I__7157\ : Odrv4
    port map (
            O => \N__29118\,
            I => \tok.n11_adj_649\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__29113\,
            I => \tok.n11_adj_649\
        );

    \I__7155\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29096\
        );

    \I__7154\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29096\
        );

    \I__7153\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29085\
        );

    \I__7152\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29085\
        );

    \I__7151\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29085\
        );

    \I__7150\ : InMux
    port map (
            O => \N__29103\,
            I => \N__29085\
        );

    \I__7149\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29085\
        );

    \I__7148\ : SRMux
    port map (
            O => \N__29101\,
            I => \N__29082\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__29096\,
            I => \N__29072\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__29085\,
            I => \N__29072\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__29082\,
            I => \N__29069\
        );

    \I__7144\ : InMux
    port map (
            O => \N__29081\,
            I => \N__29064\
        );

    \I__7143\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29064\
        );

    \I__7142\ : InMux
    port map (
            O => \N__29079\,
            I => \N__29057\
        );

    \I__7141\ : InMux
    port map (
            O => \N__29078\,
            I => \N__29057\
        );

    \I__7140\ : InMux
    port map (
            O => \N__29077\,
            I => \N__29057\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__29072\,
            I => \N__29054\
        );

    \I__7138\ : Span4Mux_h
    port map (
            O => \N__29069\,
            I => \N__29051\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__29064\,
            I => \N__29046\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__29057\,
            I => \N__29046\
        );

    \I__7135\ : Span4Mux_h
    port map (
            O => \N__29054\,
            I => \N__29043\
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__29051\,
            I => \tok.write_flag\
        );

    \I__7133\ : Odrv12
    port map (
            O => \N__29046\,
            I => \tok.write_flag\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__29043\,
            I => \tok.write_flag\
        );

    \I__7131\ : InMux
    port map (
            O => \N__29036\,
            I => \N__29022\
        );

    \I__7130\ : InMux
    port map (
            O => \N__29035\,
            I => \N__29019\
        );

    \I__7129\ : InMux
    port map (
            O => \N__29034\,
            I => \N__29010\
        );

    \I__7128\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29010\
        );

    \I__7127\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29010\
        );

    \I__7126\ : InMux
    port map (
            O => \N__29031\,
            I => \N__29010\
        );

    \I__7125\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29000\
        );

    \I__7124\ : InMux
    port map (
            O => \N__29029\,
            I => \N__29000\
        );

    \I__7123\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29000\
        );

    \I__7122\ : InMux
    port map (
            O => \N__29027\,
            I => \N__28991\
        );

    \I__7121\ : InMux
    port map (
            O => \N__29026\,
            I => \N__28991\
        );

    \I__7120\ : InMux
    port map (
            O => \N__29025\,
            I => \N__28991\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__29022\,
            I => \N__28986\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__29019\,
            I => \N__28981\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__29010\,
            I => \N__28981\
        );

    \I__7116\ : InMux
    port map (
            O => \N__29009\,
            I => \N__28974\
        );

    \I__7115\ : InMux
    port map (
            O => \N__29008\,
            I => \N__28974\
        );

    \I__7114\ : InMux
    port map (
            O => \N__29007\,
            I => \N__28974\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__29000\,
            I => \N__28968\
        );

    \I__7112\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28963\
        );

    \I__7111\ : InMux
    port map (
            O => \N__28998\,
            I => \N__28963\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__28991\,
            I => \N__28959\
        );

    \I__7109\ : InMux
    port map (
            O => \N__28990\,
            I => \N__28956\
        );

    \I__7108\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28953\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__28986\,
            I => \N__28950\
        );

    \I__7106\ : Span4Mux_s2_v
    port map (
            O => \N__28981\,
            I => \N__28945\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__28974\,
            I => \N__28945\
        );

    \I__7104\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28942\
        );

    \I__7103\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28936\
        );

    \I__7102\ : InMux
    port map (
            O => \N__28971\,
            I => \N__28931\
        );

    \I__7101\ : Span4Mux_v
    port map (
            O => \N__28968\,
            I => \N__28926\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__28963\,
            I => \N__28926\
        );

    \I__7099\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28923\
        );

    \I__7098\ : Span4Mux_h
    port map (
            O => \N__28959\,
            I => \N__28920\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__28956\,
            I => \N__28917\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__28953\,
            I => \N__28914\
        );

    \I__7095\ : Span4Mux_h
    port map (
            O => \N__28950\,
            I => \N__28907\
        );

    \I__7094\ : Span4Mux_v
    port map (
            O => \N__28945\,
            I => \N__28907\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__28942\,
            I => \N__28907\
        );

    \I__7092\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28900\
        );

    \I__7091\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28895\
        );

    \I__7090\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28895\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__28936\,
            I => \N__28892\
        );

    \I__7088\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28887\
        );

    \I__7087\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28887\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__28931\,
            I => \N__28884\
        );

    \I__7085\ : Span4Mux_h
    port map (
            O => \N__28926\,
            I => \N__28881\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__28923\,
            I => \N__28876\
        );

    \I__7083\ : Span4Mux_h
    port map (
            O => \N__28920\,
            I => \N__28876\
        );

    \I__7082\ : Span4Mux_v
    port map (
            O => \N__28917\,
            I => \N__28869\
        );

    \I__7081\ : Span4Mux_v
    port map (
            O => \N__28914\,
            I => \N__28869\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__28907\,
            I => \N__28869\
        );

    \I__7079\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28866\
        );

    \I__7078\ : InMux
    port map (
            O => \N__28905\,
            I => \N__28859\
        );

    \I__7077\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28859\
        );

    \I__7076\ : InMux
    port map (
            O => \N__28903\,
            I => \N__28859\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__28900\,
            I => \N__28850\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__28895\,
            I => \N__28850\
        );

    \I__7073\ : Span12Mux_s6_v
    port map (
            O => \N__28892\,
            I => \N__28850\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__28887\,
            I => \N__28850\
        );

    \I__7071\ : Odrv4
    port map (
            O => \N__28884\,
            I => \tok.T_4\
        );

    \I__7070\ : Odrv4
    port map (
            O => \N__28881\,
            I => \tok.T_4\
        );

    \I__7069\ : Odrv4
    port map (
            O => \N__28876\,
            I => \tok.T_4\
        );

    \I__7068\ : Odrv4
    port map (
            O => \N__28869\,
            I => \tok.T_4\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__28866\,
            I => \tok.T_4\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__28859\,
            I => \tok.T_4\
        );

    \I__7065\ : Odrv12
    port map (
            O => \N__28850\,
            I => \tok.T_4\
        );

    \I__7064\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28823\
        );

    \I__7063\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28823\
        );

    \I__7062\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28816\
        );

    \I__7061\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28816\
        );

    \I__7060\ : CascadeMux
    port map (
            O => \N__28831\,
            I => \N__28813\
        );

    \I__7059\ : InMux
    port map (
            O => \N__28830\,
            I => \N__28809\
        );

    \I__7058\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28804\
        );

    \I__7057\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28801\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__28823\,
            I => \N__28798\
        );

    \I__7055\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28793\
        );

    \I__7054\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28793\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__28816\,
            I => \N__28790\
        );

    \I__7052\ : InMux
    port map (
            O => \N__28813\,
            I => \N__28785\
        );

    \I__7051\ : InMux
    port map (
            O => \N__28812\,
            I => \N__28785\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__28809\,
            I => \N__28782\
        );

    \I__7049\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28779\
        );

    \I__7048\ : CascadeMux
    port map (
            O => \N__28807\,
            I => \N__28776\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__28804\,
            I => \N__28770\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__28801\,
            I => \N__28767\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__28798\,
            I => \N__28764\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__28793\,
            I => \N__28757\
        );

    \I__7043\ : Span4Mux_v
    port map (
            O => \N__28790\,
            I => \N__28757\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__28785\,
            I => \N__28757\
        );

    \I__7041\ : Span4Mux_s3_h
    port map (
            O => \N__28782\,
            I => \N__28752\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__28779\,
            I => \N__28752\
        );

    \I__7039\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28747\
        );

    \I__7038\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28747\
        );

    \I__7037\ : CascadeMux
    port map (
            O => \N__28774\,
            I => \N__28743\
        );

    \I__7036\ : CascadeMux
    port map (
            O => \N__28773\,
            I => \N__28740\
        );

    \I__7035\ : Span4Mux_h
    port map (
            O => \N__28770\,
            I => \N__28736\
        );

    \I__7034\ : Span4Mux_h
    port map (
            O => \N__28767\,
            I => \N__28733\
        );

    \I__7033\ : Span4Mux_h
    port map (
            O => \N__28764\,
            I => \N__28728\
        );

    \I__7032\ : Span4Mux_h
    port map (
            O => \N__28757\,
            I => \N__28728\
        );

    \I__7031\ : Span4Mux_v
    port map (
            O => \N__28752\,
            I => \N__28723\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__28747\,
            I => \N__28723\
        );

    \I__7029\ : InMux
    port map (
            O => \N__28746\,
            I => \N__28720\
        );

    \I__7028\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28713\
        );

    \I__7027\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28713\
        );

    \I__7026\ : InMux
    port map (
            O => \N__28739\,
            I => \N__28713\
        );

    \I__7025\ : Odrv4
    port map (
            O => \N__28736\,
            I => \tok.T_7\
        );

    \I__7024\ : Odrv4
    port map (
            O => \N__28733\,
            I => \tok.T_7\
        );

    \I__7023\ : Odrv4
    port map (
            O => \N__28728\,
            I => \tok.T_7\
        );

    \I__7022\ : Odrv4
    port map (
            O => \N__28723\,
            I => \tok.T_7\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__28720\,
            I => \tok.T_7\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__28713\,
            I => \tok.T_7\
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__28700\,
            I => \N__28694\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__28699\,
            I => \N__28686\
        );

    \I__7017\ : InMux
    port map (
            O => \N__28698\,
            I => \N__28683\
        );

    \I__7016\ : InMux
    port map (
            O => \N__28697\,
            I => \N__28680\
        );

    \I__7015\ : InMux
    port map (
            O => \N__28694\,
            I => \N__28671\
        );

    \I__7014\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28671\
        );

    \I__7013\ : InMux
    port map (
            O => \N__28692\,
            I => \N__28671\
        );

    \I__7012\ : InMux
    port map (
            O => \N__28691\,
            I => \N__28668\
        );

    \I__7011\ : InMux
    port map (
            O => \N__28690\,
            I => \N__28663\
        );

    \I__7010\ : InMux
    port map (
            O => \N__28689\,
            I => \N__28663\
        );

    \I__7009\ : InMux
    port map (
            O => \N__28686\,
            I => \N__28659\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__28683\,
            I => \N__28655\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__28680\,
            I => \N__28652\
        );

    \I__7006\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28649\
        );

    \I__7005\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28646\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__28671\,
            I => \N__28643\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__28668\,
            I => \N__28638\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28638\
        );

    \I__7001\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28635\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__28659\,
            I => \N__28631\
        );

    \I__6999\ : InMux
    port map (
            O => \N__28658\,
            I => \N__28628\
        );

    \I__6998\ : Span4Mux_s3_v
    port map (
            O => \N__28655\,
            I => \N__28622\
        );

    \I__6997\ : Span4Mux_s2_v
    port map (
            O => \N__28652\,
            I => \N__28617\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__28649\,
            I => \N__28617\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__28646\,
            I => \N__28608\
        );

    \I__6994\ : Span4Mux_v
    port map (
            O => \N__28643\,
            I => \N__28608\
        );

    \I__6993\ : Span4Mux_v
    port map (
            O => \N__28638\,
            I => \N__28608\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__28635\,
            I => \N__28608\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__28634\,
            I => \N__28605\
        );

    \I__6990\ : Span4Mux_s3_h
    port map (
            O => \N__28631\,
            I => \N__28600\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__28628\,
            I => \N__28600\
        );

    \I__6988\ : InMux
    port map (
            O => \N__28627\,
            I => \N__28595\
        );

    \I__6987\ : InMux
    port map (
            O => \N__28626\,
            I => \N__28595\
        );

    \I__6986\ : CascadeMux
    port map (
            O => \N__28625\,
            I => \N__28591\
        );

    \I__6985\ : Span4Mux_v
    port map (
            O => \N__28622\,
            I => \N__28585\
        );

    \I__6984\ : Span4Mux_v
    port map (
            O => \N__28617\,
            I => \N__28585\
        );

    \I__6983\ : Span4Mux_h
    port map (
            O => \N__28608\,
            I => \N__28582\
        );

    \I__6982\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28579\
        );

    \I__6981\ : Span4Mux_v
    port map (
            O => \N__28600\,
            I => \N__28574\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__28595\,
            I => \N__28574\
        );

    \I__6979\ : InMux
    port map (
            O => \N__28594\,
            I => \N__28567\
        );

    \I__6978\ : InMux
    port map (
            O => \N__28591\,
            I => \N__28567\
        );

    \I__6977\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28567\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__28585\,
            I => \tok.T_5\
        );

    \I__6975\ : Odrv4
    port map (
            O => \N__28582\,
            I => \tok.T_5\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__28579\,
            I => \tok.T_5\
        );

    \I__6973\ : Odrv4
    port map (
            O => \N__28574\,
            I => \tok.T_5\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__28567\,
            I => \tok.T_5\
        );

    \I__6971\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28551\
        );

    \I__6970\ : CascadeMux
    port map (
            O => \N__28555\,
            I => \N__28545\
        );

    \I__6969\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28539\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__28551\,
            I => \N__28536\
        );

    \I__6967\ : InMux
    port map (
            O => \N__28550\,
            I => \N__28533\
        );

    \I__6966\ : InMux
    port map (
            O => \N__28549\,
            I => \N__28525\
        );

    \I__6965\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28518\
        );

    \I__6964\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28518\
        );

    \I__6963\ : CascadeMux
    port map (
            O => \N__28544\,
            I => \N__28514\
        );

    \I__6962\ : InMux
    port map (
            O => \N__28543\,
            I => \N__28509\
        );

    \I__6961\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28506\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28501\
        );

    \I__6959\ : Span4Mux_v
    port map (
            O => \N__28536\,
            I => \N__28498\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__28533\,
            I => \N__28495\
        );

    \I__6957\ : InMux
    port map (
            O => \N__28532\,
            I => \N__28492\
        );

    \I__6956\ : InMux
    port map (
            O => \N__28531\,
            I => \N__28489\
        );

    \I__6955\ : InMux
    port map (
            O => \N__28530\,
            I => \N__28486\
        );

    \I__6954\ : InMux
    port map (
            O => \N__28529\,
            I => \N__28481\
        );

    \I__6953\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28481\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__28525\,
            I => \N__28478\
        );

    \I__6951\ : InMux
    port map (
            O => \N__28524\,
            I => \N__28473\
        );

    \I__6950\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28473\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__28518\,
            I => \N__28470\
        );

    \I__6948\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28465\
        );

    \I__6947\ : InMux
    port map (
            O => \N__28514\,
            I => \N__28465\
        );

    \I__6946\ : InMux
    port map (
            O => \N__28513\,
            I => \N__28460\
        );

    \I__6945\ : InMux
    port map (
            O => \N__28512\,
            I => \N__28460\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__28509\,
            I => \N__28454\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__28506\,
            I => \N__28454\
        );

    \I__6942\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28451\
        );

    \I__6941\ : InMux
    port map (
            O => \N__28504\,
            I => \N__28446\
        );

    \I__6940\ : Span4Mux_v
    port map (
            O => \N__28501\,
            I => \N__28439\
        );

    \I__6939\ : Span4Mux_s0_h
    port map (
            O => \N__28498\,
            I => \N__28439\
        );

    \I__6938\ : Span4Mux_v
    port map (
            O => \N__28495\,
            I => \N__28439\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__28492\,
            I => \N__28436\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__28489\,
            I => \N__28431\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__28486\,
            I => \N__28431\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__28481\,
            I => \N__28428\
        );

    \I__6933\ : Span4Mux_h
    port map (
            O => \N__28478\,
            I => \N__28417\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__28473\,
            I => \N__28417\
        );

    \I__6931\ : Span4Mux_h
    port map (
            O => \N__28470\,
            I => \N__28417\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__28465\,
            I => \N__28417\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__28460\,
            I => \N__28417\
        );

    \I__6928\ : InMux
    port map (
            O => \N__28459\,
            I => \N__28413\
        );

    \I__6927\ : Span4Mux_s3_h
    port map (
            O => \N__28454\,
            I => \N__28408\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__28451\,
            I => \N__28408\
        );

    \I__6925\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28403\
        );

    \I__6924\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28403\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__28446\,
            I => \N__28397\
        );

    \I__6922\ : Sp12to4
    port map (
            O => \N__28439\,
            I => \N__28394\
        );

    \I__6921\ : Span4Mux_s2_h
    port map (
            O => \N__28436\,
            I => \N__28391\
        );

    \I__6920\ : Span4Mux_h
    port map (
            O => \N__28431\,
            I => \N__28388\
        );

    \I__6919\ : Span4Mux_v
    port map (
            O => \N__28428\,
            I => \N__28383\
        );

    \I__6918\ : Span4Mux_v
    port map (
            O => \N__28417\,
            I => \N__28383\
        );

    \I__6917\ : InMux
    port map (
            O => \N__28416\,
            I => \N__28380\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__28413\,
            I => \N__28373\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__28408\,
            I => \N__28373\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__28403\,
            I => \N__28373\
        );

    \I__6913\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28366\
        );

    \I__6912\ : InMux
    port map (
            O => \N__28401\,
            I => \N__28366\
        );

    \I__6911\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28366\
        );

    \I__6910\ : Odrv4
    port map (
            O => \N__28397\,
            I => \tok.T_6\
        );

    \I__6909\ : Odrv12
    port map (
            O => \N__28394\,
            I => \tok.T_6\
        );

    \I__6908\ : Odrv4
    port map (
            O => \N__28391\,
            I => \tok.T_6\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__28388\,
            I => \tok.T_6\
        );

    \I__6906\ : Odrv4
    port map (
            O => \N__28383\,
            I => \tok.T_6\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__28380\,
            I => \tok.T_6\
        );

    \I__6904\ : Odrv4
    port map (
            O => \N__28373\,
            I => \tok.T_6\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__28366\,
            I => \tok.T_6\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__28349\,
            I => \N__28345\
        );

    \I__6901\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28341\
        );

    \I__6900\ : InMux
    port map (
            O => \N__28345\,
            I => \N__28338\
        );

    \I__6899\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28334\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__28341\,
            I => \N__28329\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__28338\,
            I => \N__28329\
        );

    \I__6896\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28326\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__28334\,
            I => \N__28316\
        );

    \I__6894\ : Span4Mux_v
    port map (
            O => \N__28329\,
            I => \N__28316\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__28326\,
            I => \N__28316\
        );

    \I__6892\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28313\
        );

    \I__6891\ : InMux
    port map (
            O => \N__28324\,
            I => \N__28308\
        );

    \I__6890\ : InMux
    port map (
            O => \N__28323\,
            I => \N__28308\
        );

    \I__6889\ : Span4Mux_s3_v
    port map (
            O => \N__28316\,
            I => \N__28303\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__28313\,
            I => \N__28303\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__28308\,
            I => \N__28300\
        );

    \I__6886\ : Span4Mux_h
    port map (
            O => \N__28303\,
            I => \N__28294\
        );

    \I__6885\ : Span4Mux_s3_v
    port map (
            O => \N__28300\,
            I => \N__28294\
        );

    \I__6884\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28291\
        );

    \I__6883\ : Span4Mux_h
    port map (
            O => \N__28294\,
            I => \N__28288\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__28291\,
            I => \tok.n8\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__28288\,
            I => \tok.n8\
        );

    \I__6880\ : InMux
    port map (
            O => \N__28283\,
            I => \N__28280\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__28280\,
            I => \N__28277\
        );

    \I__6878\ : Span4Mux_h
    port map (
            O => \N__28277\,
            I => \N__28274\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__28274\,
            I => \tok.n18\
        );

    \I__6876\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28265\
        );

    \I__6875\ : CascadeMux
    port map (
            O => \N__28270\,
            I => \N__28261\
        );

    \I__6874\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28256\
        );

    \I__6873\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28248\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__28265\,
            I => \N__28245\
        );

    \I__6871\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28242\
        );

    \I__6870\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28239\
        );

    \I__6869\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28236\
        );

    \I__6868\ : InMux
    port map (
            O => \N__28259\,
            I => \N__28233\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__28256\,
            I => \N__28229\
        );

    \I__6866\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28226\
        );

    \I__6865\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28223\
        );

    \I__6864\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28220\
        );

    \I__6863\ : InMux
    port map (
            O => \N__28252\,
            I => \N__28213\
        );

    \I__6862\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28213\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__28248\,
            I => \N__28210\
        );

    \I__6860\ : Span4Mux_v
    port map (
            O => \N__28245\,
            I => \N__28207\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__28242\,
            I => \N__28202\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__28239\,
            I => \N__28202\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__28236\,
            I => \N__28199\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__28233\,
            I => \N__28196\
        );

    \I__6855\ : InMux
    port map (
            O => \N__28232\,
            I => \N__28193\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__28229\,
            I => \N__28184\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__28226\,
            I => \N__28184\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__28223\,
            I => \N__28184\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__28220\,
            I => \N__28184\
        );

    \I__6850\ : InMux
    port map (
            O => \N__28219\,
            I => \N__28179\
        );

    \I__6849\ : InMux
    port map (
            O => \N__28218\,
            I => \N__28179\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__28213\,
            I => \N__28176\
        );

    \I__6847\ : Span4Mux_v
    port map (
            O => \N__28210\,
            I => \N__28165\
        );

    \I__6846\ : Span4Mux_h
    port map (
            O => \N__28207\,
            I => \N__28165\
        );

    \I__6845\ : Span4Mux_v
    port map (
            O => \N__28202\,
            I => \N__28165\
        );

    \I__6844\ : Span4Mux_s3_h
    port map (
            O => \N__28199\,
            I => \N__28165\
        );

    \I__6843\ : Span4Mux_v
    port map (
            O => \N__28196\,
            I => \N__28165\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__28193\,
            I => \N__28162\
        );

    \I__6841\ : Span4Mux_h
    port map (
            O => \N__28184\,
            I => \N__28159\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__28179\,
            I => \tok.A_low_6\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__28176\,
            I => \tok.A_low_6\
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__28165\,
            I => \tok.A_low_6\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__28162\,
            I => \tok.A_low_6\
        );

    \I__6836\ : Odrv4
    port map (
            O => \N__28159\,
            I => \tok.A_low_6\
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__28148\,
            I => \N__28145\
        );

    \I__6834\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28142\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__28142\,
            I => \N__28139\
        );

    \I__6832\ : Span4Mux_v
    port map (
            O => \N__28139\,
            I => \N__28136\
        );

    \I__6831\ : Span4Mux_h
    port map (
            O => \N__28136\,
            I => \N__28133\
        );

    \I__6830\ : Odrv4
    port map (
            O => \N__28133\,
            I => \tok.n179\
        );

    \I__6829\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28127\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__28127\,
            I => \N__28124\
        );

    \I__6827\ : Span4Mux_h
    port map (
            O => \N__28124\,
            I => \N__28121\
        );

    \I__6826\ : Odrv4
    port map (
            O => \N__28121\,
            I => \tok.n10_adj_675\
        );

    \I__6825\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28111\
        );

    \I__6824\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28111\
        );

    \I__6823\ : InMux
    port map (
            O => \N__28116\,
            I => \N__28108\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__28111\,
            I => \N__28105\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__28108\,
            I => \N__28099\
        );

    \I__6820\ : Span4Mux_h
    port map (
            O => \N__28105\,
            I => \N__28096\
        );

    \I__6819\ : InMux
    port map (
            O => \N__28104\,
            I => \N__28093\
        );

    \I__6818\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28088\
        );

    \I__6817\ : InMux
    port map (
            O => \N__28102\,
            I => \N__28088\
        );

    \I__6816\ : Odrv4
    port map (
            O => \N__28099\,
            I => \tok.n9\
        );

    \I__6815\ : Odrv4
    port map (
            O => \N__28096\,
            I => \tok.n9\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__28093\,
            I => \tok.n9\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__28088\,
            I => \tok.n9\
        );

    \I__6812\ : CascadeMux
    port map (
            O => \N__28079\,
            I => \tok.n10_adj_675_cascade_\
        );

    \I__6811\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28068\
        );

    \I__6810\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28068\
        );

    \I__6809\ : InMux
    port map (
            O => \N__28074\,
            I => \N__28065\
        );

    \I__6808\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28062\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__28068\,
            I => \N__28059\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__28065\,
            I => \N__28051\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__28062\,
            I => \N__28048\
        );

    \I__6804\ : Span4Mux_h
    port map (
            O => \N__28059\,
            I => \N__28045\
        );

    \I__6803\ : InMux
    port map (
            O => \N__28058\,
            I => \N__28040\
        );

    \I__6802\ : InMux
    port map (
            O => \N__28057\,
            I => \N__28040\
        );

    \I__6801\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28037\
        );

    \I__6800\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28032\
        );

    \I__6799\ : InMux
    port map (
            O => \N__28054\,
            I => \N__28032\
        );

    \I__6798\ : Odrv12
    port map (
            O => \N__28051\,
            I => \tok.n2586\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__28048\,
            I => \tok.n2586\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__28045\,
            I => \tok.n2586\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__28040\,
            I => \tok.n2586\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__28037\,
            I => \tok.n2586\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__28032\,
            I => \tok.n2586\
        );

    \I__6792\ : InMux
    port map (
            O => \N__28019\,
            I => \N__28008\
        );

    \I__6791\ : InMux
    port map (
            O => \N__28018\,
            I => \N__28005\
        );

    \I__6790\ : InMux
    port map (
            O => \N__28017\,
            I => \N__28002\
        );

    \I__6789\ : InMux
    port map (
            O => \N__28016\,
            I => \N__27994\
        );

    \I__6788\ : InMux
    port map (
            O => \N__28015\,
            I => \N__27994\
        );

    \I__6787\ : InMux
    port map (
            O => \N__28014\,
            I => \N__27989\
        );

    \I__6786\ : CascadeMux
    port map (
            O => \N__28013\,
            I => \N__27983\
        );

    \I__6785\ : CascadeMux
    port map (
            O => \N__28012\,
            I => \N__27980\
        );

    \I__6784\ : CascadeMux
    port map (
            O => \N__28011\,
            I => \N__27976\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__28008\,
            I => \N__27969\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__28005\,
            I => \N__27969\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__28002\,
            I => \N__27969\
        );

    \I__6780\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27966\
        );

    \I__6779\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27963\
        );

    \I__6778\ : InMux
    port map (
            O => \N__27999\,
            I => \N__27960\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__27994\,
            I => \N__27957\
        );

    \I__6776\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27952\
        );

    \I__6775\ : InMux
    port map (
            O => \N__27992\,
            I => \N__27952\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__27989\,
            I => \N__27949\
        );

    \I__6773\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27946\
        );

    \I__6772\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27939\
        );

    \I__6771\ : InMux
    port map (
            O => \N__27986\,
            I => \N__27939\
        );

    \I__6770\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27939\
        );

    \I__6769\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27936\
        );

    \I__6768\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27931\
        );

    \I__6767\ : InMux
    port map (
            O => \N__27976\,
            I => \N__27931\
        );

    \I__6766\ : Span4Mux_s3_v
    port map (
            O => \N__27969\,
            I => \N__27920\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__27966\,
            I => \N__27915\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__27963\,
            I => \N__27915\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__27960\,
            I => \N__27908\
        );

    \I__6762\ : Span4Mux_v
    port map (
            O => \N__27957\,
            I => \N__27908\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__27952\,
            I => \N__27908\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__27949\,
            I => \N__27905\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__27946\,
            I => \N__27900\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__27939\,
            I => \N__27900\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__27936\,
            I => \N__27897\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27894\
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__27930\,
            I => \N__27891\
        );

    \I__6754\ : CascadeMux
    port map (
            O => \N__27929\,
            I => \N__27888\
        );

    \I__6753\ : CascadeMux
    port map (
            O => \N__27928\,
            I => \N__27885\
        );

    \I__6752\ : CascadeMux
    port map (
            O => \N__27927\,
            I => \N__27881\
        );

    \I__6751\ : CascadeMux
    port map (
            O => \N__27926\,
            I => \N__27876\
        );

    \I__6750\ : CascadeMux
    port map (
            O => \N__27925\,
            I => \N__27873\
        );

    \I__6749\ : CascadeMux
    port map (
            O => \N__27924\,
            I => \N__27870\
        );

    \I__6748\ : CascadeMux
    port map (
            O => \N__27923\,
            I => \N__27865\
        );

    \I__6747\ : Span4Mux_v
    port map (
            O => \N__27920\,
            I => \N__27860\
        );

    \I__6746\ : Span4Mux_v
    port map (
            O => \N__27915\,
            I => \N__27860\
        );

    \I__6745\ : Span4Mux_h
    port map (
            O => \N__27908\,
            I => \N__27857\
        );

    \I__6744\ : Span4Mux_h
    port map (
            O => \N__27905\,
            I => \N__27848\
        );

    \I__6743\ : Span4Mux_v
    port map (
            O => \N__27900\,
            I => \N__27848\
        );

    \I__6742\ : Span4Mux_v
    port map (
            O => \N__27897\,
            I => \N__27848\
        );

    \I__6741\ : Span4Mux_v
    port map (
            O => \N__27894\,
            I => \N__27848\
        );

    \I__6740\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27841\
        );

    \I__6739\ : InMux
    port map (
            O => \N__27888\,
            I => \N__27841\
        );

    \I__6738\ : InMux
    port map (
            O => \N__27885\,
            I => \N__27841\
        );

    \I__6737\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27834\
        );

    \I__6736\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27834\
        );

    \I__6735\ : InMux
    port map (
            O => \N__27880\,
            I => \N__27834\
        );

    \I__6734\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27819\
        );

    \I__6733\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27819\
        );

    \I__6732\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27819\
        );

    \I__6731\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27819\
        );

    \I__6730\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27819\
        );

    \I__6729\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27819\
        );

    \I__6728\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27819\
        );

    \I__6727\ : Odrv4
    port map (
            O => \N__27860\,
            I => \tok.T_3\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__27857\,
            I => \tok.T_3\
        );

    \I__6725\ : Odrv4
    port map (
            O => \N__27848\,
            I => \tok.T_3\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__27841\,
            I => \tok.T_3\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__27834\,
            I => \tok.T_3\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__27819\,
            I => \tok.T_3\
        );

    \I__6721\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27801\
        );

    \I__6720\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27796\
        );

    \I__6719\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27796\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__27801\,
            I => \N__27791\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__27796\,
            I => \N__27788\
        );

    \I__6716\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27785\
        );

    \I__6715\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27782\
        );

    \I__6714\ : Span4Mux_h
    port map (
            O => \N__27791\,
            I => \N__27777\
        );

    \I__6713\ : Span4Mux_h
    port map (
            O => \N__27788\,
            I => \N__27774\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__27785\,
            I => \N__27771\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__27782\,
            I => \N__27768\
        );

    \I__6710\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27763\
        );

    \I__6709\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27763\
        );

    \I__6708\ : Span4Mux_h
    port map (
            O => \N__27777\,
            I => \N__27759\
        );

    \I__6707\ : Span4Mux_h
    port map (
            O => \N__27774\,
            I => \N__27756\
        );

    \I__6706\ : Span4Mux_v
    port map (
            O => \N__27771\,
            I => \N__27749\
        );

    \I__6705\ : Span4Mux_v
    port map (
            O => \N__27768\,
            I => \N__27749\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__27763\,
            I => \N__27749\
        );

    \I__6703\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27746\
        );

    \I__6702\ : Odrv4
    port map (
            O => \N__27759\,
            I => \tok.n2178\
        );

    \I__6701\ : Odrv4
    port map (
            O => \N__27756\,
            I => \tok.n2178\
        );

    \I__6700\ : Odrv4
    port map (
            O => \N__27749\,
            I => \tok.n2178\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__27746\,
            I => \tok.n2178\
        );

    \I__6698\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27734\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__27734\,
            I => \N__27731\
        );

    \I__6696\ : Odrv12
    port map (
            O => \N__27731\,
            I => \tok.n41\
        );

    \I__6695\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27725\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__27725\,
            I => \tok.n4484\
        );

    \I__6693\ : CascadeMux
    port map (
            O => \N__27722\,
            I => \N__27719\
        );

    \I__6692\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27716\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__27716\,
            I => \tok.n40_adj_661\
        );

    \I__6690\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27710\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__27710\,
            I => \N__27707\
        );

    \I__6688\ : Odrv12
    port map (
            O => \N__27707\,
            I => \tok.n42\
        );

    \I__6687\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27701\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__27701\,
            I => \tok.n4688\
        );

    \I__6685\ : InMux
    port map (
            O => \N__27698\,
            I => \N__27695\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__27695\,
            I => \N__27692\
        );

    \I__6683\ : Span4Mux_s3_h
    port map (
            O => \N__27692\,
            I => \N__27687\
        );

    \I__6682\ : InMux
    port map (
            O => \N__27691\,
            I => \N__27684\
        );

    \I__6681\ : InMux
    port map (
            O => \N__27690\,
            I => \N__27681\
        );

    \I__6680\ : Span4Mux_v
    port map (
            O => \N__27687\,
            I => \N__27676\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27676\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__27681\,
            I => \tok.n10\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__27676\,
            I => \tok.n10\
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__27671\,
            I => \tok.n14_adj_658_cascade_\
        );

    \I__6675\ : InMux
    port map (
            O => \N__27668\,
            I => \N__27646\
        );

    \I__6674\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27646\
        );

    \I__6673\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27646\
        );

    \I__6672\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27637\
        );

    \I__6671\ : InMux
    port map (
            O => \N__27664\,
            I => \N__27637\
        );

    \I__6670\ : InMux
    port map (
            O => \N__27663\,
            I => \N__27637\
        );

    \I__6669\ : InMux
    port map (
            O => \N__27662\,
            I => \N__27637\
        );

    \I__6668\ : InMux
    port map (
            O => \N__27661\,
            I => \N__27626\
        );

    \I__6667\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27626\
        );

    \I__6666\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27626\
        );

    \I__6665\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27626\
        );

    \I__6664\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27626\
        );

    \I__6663\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27617\
        );

    \I__6662\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27617\
        );

    \I__6661\ : InMux
    port map (
            O => \N__27654\,
            I => \N__27617\
        );

    \I__6660\ : InMux
    port map (
            O => \N__27653\,
            I => \N__27617\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__27646\,
            I => \N__27614\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__27637\,
            I => \N__27607\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__27626\,
            I => \N__27607\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__27617\,
            I => \N__27607\
        );

    \I__6655\ : Span4Mux_v
    port map (
            O => \N__27614\,
            I => \N__27602\
        );

    \I__6654\ : Span4Mux_v
    port map (
            O => \N__27607\,
            I => \N__27602\
        );

    \I__6653\ : Span4Mux_h
    port map (
            O => \N__27602\,
            I => \N__27599\
        );

    \I__6652\ : Odrv4
    port map (
            O => \N__27599\,
            I => \tok.n399\
        );

    \I__6651\ : CascadeMux
    port map (
            O => \N__27596\,
            I => \N__27593\
        );

    \I__6650\ : InMux
    port map (
            O => \N__27593\,
            I => \N__27590\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__27590\,
            I => \N__27586\
        );

    \I__6648\ : InMux
    port map (
            O => \N__27589\,
            I => \N__27583\
        );

    \I__6647\ : Odrv12
    port map (
            O => \N__27586\,
            I => \tok.n14\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__27583\,
            I => \tok.n14\
        );

    \I__6645\ : CascadeMux
    port map (
            O => \N__27578\,
            I => \tok.n4422_cascade_\
        );

    \I__6644\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27572\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__27572\,
            I => \N__27567\
        );

    \I__6642\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27562\
        );

    \I__6641\ : InMux
    port map (
            O => \N__27570\,
            I => \N__27562\
        );

    \I__6640\ : Span4Mux_s3_v
    port map (
            O => \N__27567\,
            I => \N__27557\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__27562\,
            I => \N__27557\
        );

    \I__6638\ : Span4Mux_v
    port map (
            O => \N__27557\,
            I => \N__27552\
        );

    \I__6637\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27549\
        );

    \I__6636\ : InMux
    port map (
            O => \N__27555\,
            I => \N__27546\
        );

    \I__6635\ : Odrv4
    port map (
            O => \N__27552\,
            I => \tok.n11_adj_648\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__27549\,
            I => \tok.n11_adj_648\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__27546\,
            I => \tok.n11_adj_648\
        );

    \I__6632\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27533\
        );

    \I__6631\ : InMux
    port map (
            O => \N__27538\,
            I => \N__27533\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__27533\,
            I => \tok.n4558\
        );

    \I__6629\ : InMux
    port map (
            O => \N__27530\,
            I => \N__27525\
        );

    \I__6628\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27520\
        );

    \I__6627\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27520\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__27525\,
            I => \N__27517\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27514\
        );

    \I__6624\ : Odrv12
    port map (
            O => \N__27517\,
            I => \tok.n14_adj_650\
        );

    \I__6623\ : Odrv4
    port map (
            O => \N__27514\,
            I => \tok.n14_adj_650\
        );

    \I__6622\ : CascadeMux
    port map (
            O => \N__27509\,
            I => \tok.n51_cascade_\
        );

    \I__6621\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27503\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__27503\,
            I => \tok.n4424\
        );

    \I__6619\ : InMux
    port map (
            O => \N__27500\,
            I => \N__27497\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__27497\,
            I => \tok.n48\
        );

    \I__6617\ : InMux
    port map (
            O => \N__27494\,
            I => \N__27491\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__27491\,
            I => \N__27488\
        );

    \I__6615\ : Span4Mux_s3_h
    port map (
            O => \N__27488\,
            I => \N__27485\
        );

    \I__6614\ : Sp12to4
    port map (
            O => \N__27485\,
            I => \N__27482\
        );

    \I__6613\ : Odrv12
    port map (
            O => \N__27482\,
            I => \tok.table_rd_12\
        );

    \I__6612\ : InMux
    port map (
            O => \N__27479\,
            I => \N__27476\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__27476\,
            I => \N__27473\
        );

    \I__6610\ : Odrv12
    port map (
            O => \N__27473\,
            I => \tok.n5_adj_694\
        );

    \I__6609\ : InMux
    port map (
            O => \N__27470\,
            I => \N__27467\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__27467\,
            I => \N__27464\
        );

    \I__6607\ : Span4Mux_s2_h
    port map (
            O => \N__27464\,
            I => \N__27461\
        );

    \I__6606\ : Span4Mux_h
    port map (
            O => \N__27461\,
            I => \N__27458\
        );

    \I__6605\ : Odrv4
    port map (
            O => \N__27458\,
            I => \tok.n10_adj_697\
        );

    \I__6604\ : CascadeMux
    port map (
            O => \N__27455\,
            I => \tok.n14_adj_695_cascade_\
        );

    \I__6603\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27449\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__27449\,
            I => \N__27442\
        );

    \I__6601\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27439\
        );

    \I__6600\ : InMux
    port map (
            O => \N__27447\,
            I => \N__27436\
        );

    \I__6599\ : CascadeMux
    port map (
            O => \N__27446\,
            I => \N__27430\
        );

    \I__6598\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27424\
        );

    \I__6597\ : Span4Mux_h
    port map (
            O => \N__27442\,
            I => \N__27418\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__27439\,
            I => \N__27418\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__27436\,
            I => \N__27415\
        );

    \I__6594\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27412\
        );

    \I__6593\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27408\
        );

    \I__6592\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27403\
        );

    \I__6591\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27403\
        );

    \I__6590\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27400\
        );

    \I__6589\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27396\
        );

    \I__6588\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27393\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__27424\,
            I => \N__27389\
        );

    \I__6586\ : InMux
    port map (
            O => \N__27423\,
            I => \N__27386\
        );

    \I__6585\ : Span4Mux_v
    port map (
            O => \N__27418\,
            I => \N__27383\
        );

    \I__6584\ : Span4Mux_v
    port map (
            O => \N__27415\,
            I => \N__27378\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__27412\,
            I => \N__27378\
        );

    \I__6582\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27375\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__27408\,
            I => \N__27370\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__27403\,
            I => \N__27370\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__27400\,
            I => \N__27367\
        );

    \I__6578\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27364\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__27396\,
            I => \N__27359\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__27393\,
            I => \N__27359\
        );

    \I__6575\ : InMux
    port map (
            O => \N__27392\,
            I => \N__27356\
        );

    \I__6574\ : Span12Mux_s4_v
    port map (
            O => \N__27389\,
            I => \N__27353\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__27386\,
            I => \N__27346\
        );

    \I__6572\ : Span4Mux_h
    port map (
            O => \N__27383\,
            I => \N__27346\
        );

    \I__6571\ : Span4Mux_h
    port map (
            O => \N__27378\,
            I => \N__27346\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__27375\,
            I => \N__27341\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__27370\,
            I => \N__27341\
        );

    \I__6568\ : Sp12to4
    port map (
            O => \N__27367\,
            I => \N__27334\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__27364\,
            I => \N__27334\
        );

    \I__6566\ : Span12Mux_s8_h
    port map (
            O => \N__27359\,
            I => \N__27334\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__27356\,
            I => \tok.A_low_4\
        );

    \I__6564\ : Odrv12
    port map (
            O => \N__27353\,
            I => \tok.A_low_4\
        );

    \I__6563\ : Odrv4
    port map (
            O => \N__27346\,
            I => \tok.A_low_4\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__27341\,
            I => \tok.A_low_4\
        );

    \I__6561\ : Odrv12
    port map (
            O => \N__27334\,
            I => \tok.A_low_4\
        );

    \I__6560\ : InMux
    port map (
            O => \N__27323\,
            I => \N__27320\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__27320\,
            I => \N__27317\
        );

    \I__6558\ : Span4Mux_h
    port map (
            O => \N__27317\,
            I => \N__27314\
        );

    \I__6557\ : Odrv4
    port map (
            O => \N__27314\,
            I => \tok.n18_adj_698\
        );

    \I__6556\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27307\
        );

    \I__6555\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27304\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__27307\,
            I => \N__27299\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__27304\,
            I => \N__27299\
        );

    \I__6552\ : Span4Mux_v
    port map (
            O => \N__27299\,
            I => \N__27296\
        );

    \I__6551\ : Span4Mux_h
    port map (
            O => \N__27296\,
            I => \N__27293\
        );

    \I__6550\ : Odrv4
    port map (
            O => \N__27293\,
            I => \tok.n2177\
        );

    \I__6549\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27286\
        );

    \I__6548\ : InMux
    port map (
            O => \N__27289\,
            I => \N__27283\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__27286\,
            I => \tok.n14_adj_825\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__27283\,
            I => \tok.n14_adj_825\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__27278\,
            I => \tok.n2177_cascade_\
        );

    \I__6544\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27272\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__27272\,
            I => \N__27269\
        );

    \I__6542\ : Span4Mux_h
    port map (
            O => \N__27269\,
            I => \N__27263\
        );

    \I__6541\ : InMux
    port map (
            O => \N__27268\,
            I => \N__27260\
        );

    \I__6540\ : InMux
    port map (
            O => \N__27267\,
            I => \N__27257\
        );

    \I__6539\ : InMux
    port map (
            O => \N__27266\,
            I => \N__27254\
        );

    \I__6538\ : Odrv4
    port map (
            O => \N__27263\,
            I => \tok.n10_adj_646\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__27260\,
            I => \tok.n10_adj_646\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__27257\,
            I => \tok.n10_adj_646\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__27254\,
            I => \tok.n10_adj_646\
        );

    \I__6534\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27239\
        );

    \I__6533\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27236\
        );

    \I__6532\ : InMux
    port map (
            O => \N__27243\,
            I => \N__27233\
        );

    \I__6531\ : InMux
    port map (
            O => \N__27242\,
            I => \N__27229\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__27239\,
            I => \N__27225\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__27236\,
            I => \N__27222\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__27233\,
            I => \N__27219\
        );

    \I__6527\ : InMux
    port map (
            O => \N__27232\,
            I => \N__27212\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__27229\,
            I => \N__27205\
        );

    \I__6525\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27202\
        );

    \I__6524\ : Span4Mux_h
    port map (
            O => \N__27225\,
            I => \N__27199\
        );

    \I__6523\ : Span4Mux_h
    port map (
            O => \N__27222\,
            I => \N__27196\
        );

    \I__6522\ : Span4Mux_h
    port map (
            O => \N__27219\,
            I => \N__27193\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__27218\,
            I => \N__27189\
        );

    \I__6520\ : InMux
    port map (
            O => \N__27217\,
            I => \N__27181\
        );

    \I__6519\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27181\
        );

    \I__6518\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27181\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__27212\,
            I => \N__27178\
        );

    \I__6516\ : InMux
    port map (
            O => \N__27211\,
            I => \N__27169\
        );

    \I__6515\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27169\
        );

    \I__6514\ : InMux
    port map (
            O => \N__27209\,
            I => \N__27169\
        );

    \I__6513\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27169\
        );

    \I__6512\ : Span4Mux_h
    port map (
            O => \N__27205\,
            I => \N__27163\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__27202\,
            I => \N__27163\
        );

    \I__6510\ : Span4Mux_h
    port map (
            O => \N__27199\,
            I => \N__27160\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__27196\,
            I => \N__27155\
        );

    \I__6508\ : Span4Mux_h
    port map (
            O => \N__27193\,
            I => \N__27155\
        );

    \I__6507\ : InMux
    port map (
            O => \N__27192\,
            I => \N__27148\
        );

    \I__6506\ : InMux
    port map (
            O => \N__27189\,
            I => \N__27148\
        );

    \I__6505\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27148\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__27181\,
            I => \N__27141\
        );

    \I__6503\ : Span12Mux_s5_v
    port map (
            O => \N__27178\,
            I => \N__27141\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__27169\,
            I => \N__27141\
        );

    \I__6501\ : InMux
    port map (
            O => \N__27168\,
            I => \N__27138\
        );

    \I__6500\ : Span4Mux_h
    port map (
            O => \N__27163\,
            I => \N__27135\
        );

    \I__6499\ : Odrv4
    port map (
            O => \N__27160\,
            I => \tok.n132\
        );

    \I__6498\ : Odrv4
    port map (
            O => \N__27155\,
            I => \tok.n132\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__27148\,
            I => \tok.n132\
        );

    \I__6496\ : Odrv12
    port map (
            O => \N__27141\,
            I => \tok.n132\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__27138\,
            I => \tok.n132\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__27135\,
            I => \tok.n132\
        );

    \I__6493\ : InMux
    port map (
            O => \N__27122\,
            I => \N__27119\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__27119\,
            I => \N__27116\
        );

    \I__6491\ : Span12Mux_s1_h
    port map (
            O => \N__27116\,
            I => \N__27113\
        );

    \I__6490\ : Odrv12
    port map (
            O => \N__27113\,
            I => \tok.table_rd_8\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__27110\,
            I => \tok.n132_cascade_\
        );

    \I__6488\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27104\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__27104\,
            I => \N__27101\
        );

    \I__6486\ : Odrv4
    port map (
            O => \N__27101\,
            I => \tok.n5\
        );

    \I__6485\ : InMux
    port map (
            O => \N__27098\,
            I => \N__27095\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__27095\,
            I => \N__27092\
        );

    \I__6483\ : Span4Mux_h
    port map (
            O => \N__27092\,
            I => \N__27089\
        );

    \I__6482\ : Span4Mux_h
    port map (
            O => \N__27089\,
            I => \N__27086\
        );

    \I__6481\ : Odrv4
    port map (
            O => \N__27086\,
            I => \tok.n10_adj_652\
        );

    \I__6480\ : InMux
    port map (
            O => \N__27083\,
            I => \N__27080\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__27080\,
            I => \N__27077\
        );

    \I__6478\ : Odrv4
    port map (
            O => \N__27077\,
            I => \tok.n14_adj_651\
        );

    \I__6477\ : CascadeMux
    port map (
            O => \N__27074\,
            I => \N__27068\
        );

    \I__6476\ : CascadeMux
    port map (
            O => \N__27073\,
            I => \N__27064\
        );

    \I__6475\ : CascadeMux
    port map (
            O => \N__27072\,
            I => \N__27058\
        );

    \I__6474\ : CascadeMux
    port map (
            O => \N__27071\,
            I => \N__27054\
        );

    \I__6473\ : InMux
    port map (
            O => \N__27068\,
            I => \N__27051\
        );

    \I__6472\ : InMux
    port map (
            O => \N__27067\,
            I => \N__27047\
        );

    \I__6471\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27042\
        );

    \I__6470\ : InMux
    port map (
            O => \N__27063\,
            I => \N__27039\
        );

    \I__6469\ : InMux
    port map (
            O => \N__27062\,
            I => \N__27036\
        );

    \I__6468\ : CascadeMux
    port map (
            O => \N__27061\,
            I => \N__27033\
        );

    \I__6467\ : InMux
    port map (
            O => \N__27058\,
            I => \N__27030\
        );

    \I__6466\ : InMux
    port map (
            O => \N__27057\,
            I => \N__27027\
        );

    \I__6465\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27024\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__27051\,
            I => \N__27021\
        );

    \I__6463\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27018\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__27047\,
            I => \N__27015\
        );

    \I__6461\ : InMux
    port map (
            O => \N__27046\,
            I => \N__27012\
        );

    \I__6460\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27009\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__27042\,
            I => \N__27006\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__27039\,
            I => \N__27001\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__27036\,
            I => \N__27001\
        );

    \I__6456\ : InMux
    port map (
            O => \N__27033\,
            I => \N__26998\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__27030\,
            I => \N__26991\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__27027\,
            I => \N__26991\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__26991\
        );

    \I__6452\ : Span4Mux_v
    port map (
            O => \N__27021\,
            I => \N__26988\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__27018\,
            I => \N__26985\
        );

    \I__6450\ : Span4Mux_v
    port map (
            O => \N__27015\,
            I => \N__26980\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__27012\,
            I => \N__26980\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__27009\,
            I => \N__26977\
        );

    \I__6447\ : Span4Mux_v
    port map (
            O => \N__27006\,
            I => \N__26974\
        );

    \I__6446\ : Span4Mux_h
    port map (
            O => \N__27001\,
            I => \N__26971\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__26998\,
            I => \N__26968\
        );

    \I__6444\ : Span4Mux_v
    port map (
            O => \N__26991\,
            I => \N__26963\
        );

    \I__6443\ : Span4Mux_h
    port map (
            O => \N__26988\,
            I => \N__26963\
        );

    \I__6442\ : Span4Mux_v
    port map (
            O => \N__26985\,
            I => \N__26958\
        );

    \I__6441\ : Span4Mux_h
    port map (
            O => \N__26980\,
            I => \N__26958\
        );

    \I__6440\ : Span4Mux_s3_h
    port map (
            O => \N__26977\,
            I => \N__26955\
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__26974\,
            I => \tok.n109\
        );

    \I__6438\ : Odrv4
    port map (
            O => \N__26971\,
            I => \tok.n109\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__26968\,
            I => \tok.n109\
        );

    \I__6436\ : Odrv4
    port map (
            O => \N__26963\,
            I => \tok.n109\
        );

    \I__6435\ : Odrv4
    port map (
            O => \N__26958\,
            I => \tok.n109\
        );

    \I__6434\ : Odrv4
    port map (
            O => \N__26955\,
            I => \tok.n109\
        );

    \I__6433\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26938\
        );

    \I__6432\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26935\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__26938\,
            I => \N__26930\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__26935\,
            I => \N__26922\
        );

    \I__6429\ : InMux
    port map (
            O => \N__26934\,
            I => \N__26916\
        );

    \I__6428\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26913\
        );

    \I__6427\ : Span4Mux_v
    port map (
            O => \N__26930\,
            I => \N__26910\
        );

    \I__6426\ : InMux
    port map (
            O => \N__26929\,
            I => \N__26907\
        );

    \I__6425\ : InMux
    port map (
            O => \N__26928\,
            I => \N__26904\
        );

    \I__6424\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26901\
        );

    \I__6423\ : InMux
    port map (
            O => \N__26926\,
            I => \N__26894\
        );

    \I__6422\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26894\
        );

    \I__6421\ : Span4Mux_v
    port map (
            O => \N__26922\,
            I => \N__26891\
        );

    \I__6420\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26886\
        );

    \I__6419\ : InMux
    port map (
            O => \N__26920\,
            I => \N__26886\
        );

    \I__6418\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26883\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__26916\,
            I => \N__26879\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__26913\,
            I => \N__26876\
        );

    \I__6415\ : Span4Mux_h
    port map (
            O => \N__26910\,
            I => \N__26871\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26871\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__26904\,
            I => \N__26866\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__26901\,
            I => \N__26866\
        );

    \I__6411\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26863\
        );

    \I__6410\ : InMux
    port map (
            O => \N__26899\,
            I => \N__26860\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__26894\,
            I => \N__26857\
        );

    \I__6408\ : Span4Mux_h
    port map (
            O => \N__26891\,
            I => \N__26850\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__26886\,
            I => \N__26850\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__26883\,
            I => \N__26850\
        );

    \I__6405\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26847\
        );

    \I__6404\ : Span4Mux_v
    port map (
            O => \N__26879\,
            I => \N__26840\
        );

    \I__6403\ : Span4Mux_s3_h
    port map (
            O => \N__26876\,
            I => \N__26840\
        );

    \I__6402\ : Span4Mux_v
    port map (
            O => \N__26871\,
            I => \N__26840\
        );

    \I__6401\ : Span4Mux_h
    port map (
            O => \N__26866\,
            I => \N__26835\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__26863\,
            I => \N__26835\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__26860\,
            I => \N__26832\
        );

    \I__6398\ : Odrv4
    port map (
            O => \N__26857\,
            I => \tok.A_low_0\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__26850\,
            I => \tok.A_low_0\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__26847\,
            I => \tok.A_low_0\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__26840\,
            I => \tok.A_low_0\
        );

    \I__6394\ : Odrv4
    port map (
            O => \N__26835\,
            I => \tok.A_low_0\
        );

    \I__6393\ : Odrv4
    port map (
            O => \N__26832\,
            I => \tok.A_low_0\
        );

    \I__6392\ : CascadeMux
    port map (
            O => \N__26819\,
            I => \tok.ram.n14_adj_631_cascade_\
        );

    \I__6391\ : InMux
    port map (
            O => \N__26816\,
            I => \N__26805\
        );

    \I__6390\ : InMux
    port map (
            O => \N__26815\,
            I => \N__26805\
        );

    \I__6389\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26800\
        );

    \I__6388\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26797\
        );

    \I__6387\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26792\
        );

    \I__6386\ : InMux
    port map (
            O => \N__26811\,
            I => \N__26784\
        );

    \I__6385\ : InMux
    port map (
            O => \N__26810\,
            I => \N__26784\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__26805\,
            I => \N__26781\
        );

    \I__6383\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26776\
        );

    \I__6382\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26776\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__26800\,
            I => \N__26773\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__26797\,
            I => \N__26770\
        );

    \I__6379\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26765\
        );

    \I__6378\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26765\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__26792\,
            I => \N__26762\
        );

    \I__6376\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26759\
        );

    \I__6375\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26754\
        );

    \I__6374\ : InMux
    port map (
            O => \N__26789\,
            I => \N__26754\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__26784\,
            I => \N__26749\
        );

    \I__6372\ : Span4Mux_s3_v
    port map (
            O => \N__26781\,
            I => \N__26749\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__26776\,
            I => \N__26742\
        );

    \I__6370\ : Span4Mux_h
    port map (
            O => \N__26773\,
            I => \N__26742\
        );

    \I__6369\ : Span4Mux_s3_v
    port map (
            O => \N__26770\,
            I => \N__26742\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__26765\,
            I => \N__26739\
        );

    \I__6367\ : Span4Mux_h
    port map (
            O => \N__26762\,
            I => \N__26734\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__26759\,
            I => \N__26734\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26731\
        );

    \I__6364\ : Span4Mux_v
    port map (
            O => \N__26749\,
            I => \N__26727\
        );

    \I__6363\ : Span4Mux_v
    port map (
            O => \N__26742\,
            I => \N__26724\
        );

    \I__6362\ : Span4Mux_v
    port map (
            O => \N__26739\,
            I => \N__26717\
        );

    \I__6361\ : Span4Mux_v
    port map (
            O => \N__26734\,
            I => \N__26717\
        );

    \I__6360\ : Span4Mux_h
    port map (
            O => \N__26731\,
            I => \N__26717\
        );

    \I__6359\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26714\
        );

    \I__6358\ : Sp12to4
    port map (
            O => \N__26727\,
            I => \N__26709\
        );

    \I__6357\ : Sp12to4
    port map (
            O => \N__26724\,
            I => \N__26709\
        );

    \I__6356\ : Span4Mux_h
    port map (
            O => \N__26717\,
            I => \N__26706\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__26714\,
            I => \N__26703\
        );

    \I__6354\ : Odrv12
    port map (
            O => \N__26709\,
            I => \tok.n2635\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__26706\,
            I => \tok.n2635\
        );

    \I__6352\ : Odrv4
    port map (
            O => \N__26703\,
            I => \tok.n2635\
        );

    \I__6351\ : InMux
    port map (
            O => \N__26696\,
            I => \N__26691\
        );

    \I__6350\ : InMux
    port map (
            O => \N__26695\,
            I => \N__26688\
        );

    \I__6349\ : InMux
    port map (
            O => \N__26694\,
            I => \N__26685\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__26691\,
            I => \N__26679\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__26688\,
            I => \N__26674\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__26685\,
            I => \N__26674\
        );

    \I__6345\ : InMux
    port map (
            O => \N__26684\,
            I => \N__26670\
        );

    \I__6344\ : InMux
    port map (
            O => \N__26683\,
            I => \N__26667\
        );

    \I__6343\ : InMux
    port map (
            O => \N__26682\,
            I => \N__26664\
        );

    \I__6342\ : Span4Mux_h
    port map (
            O => \N__26679\,
            I => \N__26659\
        );

    \I__6341\ : Span4Mux_v
    port map (
            O => \N__26674\,
            I => \N__26659\
        );

    \I__6340\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26656\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__26670\,
            I => \N__26651\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__26667\,
            I => \N__26651\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__26664\,
            I => \N__26647\
        );

    \I__6336\ : Span4Mux_h
    port map (
            O => \N__26659\,
            I => \N__26644\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__26656\,
            I => \N__26639\
        );

    \I__6334\ : Span4Mux_h
    port map (
            O => \N__26651\,
            I => \N__26639\
        );

    \I__6333\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26636\
        );

    \I__6332\ : Odrv4
    port map (
            O => \N__26647\,
            I => \tok.n4_adj_795\
        );

    \I__6331\ : Odrv4
    port map (
            O => \N__26644\,
            I => \tok.n4_adj_795\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__26639\,
            I => \tok.n4_adj_795\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__26636\,
            I => \tok.n4_adj_795\
        );

    \I__6328\ : CascadeMux
    port map (
            O => \N__26627\,
            I => \tok.n41_cascade_\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__26624\,
            I => \N__26619\
        );

    \I__6326\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26610\
        );

    \I__6325\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26610\
        );

    \I__6324\ : InMux
    port map (
            O => \N__26619\,
            I => \N__26605\
        );

    \I__6323\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26605\
        );

    \I__6322\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26592\
        );

    \I__6321\ : InMux
    port map (
            O => \N__26616\,
            I => \N__26592\
        );

    \I__6320\ : InMux
    port map (
            O => \N__26615\,
            I => \N__26589\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__26610\,
            I => \N__26584\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__26605\,
            I => \N__26584\
        );

    \I__6317\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26581\
        );

    \I__6316\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26578\
        );

    \I__6315\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26573\
        );

    \I__6314\ : InMux
    port map (
            O => \N__26601\,
            I => \N__26573\
        );

    \I__6313\ : InMux
    port map (
            O => \N__26600\,
            I => \N__26570\
        );

    \I__6312\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26567\
        );

    \I__6311\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26564\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__26597\,
            I => \N__26559\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__26592\,
            I => \N__26554\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__26589\,
            I => \N__26554\
        );

    \I__6307\ : Span4Mux_h
    port map (
            O => \N__26584\,
            I => \N__26549\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__26581\,
            I => \N__26549\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__26578\,
            I => \N__26544\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__26573\,
            I => \N__26544\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__26570\,
            I => \N__26539\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__26567\,
            I => \N__26539\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__26564\,
            I => \N__26536\
        );

    \I__6300\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26529\
        );

    \I__6299\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26529\
        );

    \I__6298\ : InMux
    port map (
            O => \N__26559\,
            I => \N__26529\
        );

    \I__6297\ : Span4Mux_v
    port map (
            O => \N__26554\,
            I => \N__26526\
        );

    \I__6296\ : Span4Mux_v
    port map (
            O => \N__26549\,
            I => \N__26521\
        );

    \I__6295\ : Span4Mux_v
    port map (
            O => \N__26544\,
            I => \N__26521\
        );

    \I__6294\ : Span4Mux_s3_v
    port map (
            O => \N__26539\,
            I => \N__26514\
        );

    \I__6293\ : Span4Mux_h
    port map (
            O => \N__26536\,
            I => \N__26514\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__26529\,
            I => \N__26514\
        );

    \I__6291\ : Sp12to4
    port map (
            O => \N__26526\,
            I => \N__26511\
        );

    \I__6290\ : Span4Mux_h
    port map (
            O => \N__26521\,
            I => \N__26508\
        );

    \I__6289\ : Span4Mux_v
    port map (
            O => \N__26514\,
            I => \N__26505\
        );

    \I__6288\ : Odrv12
    port map (
            O => \N__26511\,
            I => \tok.n884\
        );

    \I__6287\ : Odrv4
    port map (
            O => \N__26508\,
            I => \tok.n884\
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__26505\,
            I => \tok.n884\
        );

    \I__6285\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26494\
        );

    \I__6284\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26491\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__26494\,
            I => \tok.n14_adj_702\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__26491\,
            I => \tok.n14_adj_702\
        );

    \I__6281\ : InMux
    port map (
            O => \N__26486\,
            I => \N__26482\
        );

    \I__6280\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26479\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__26482\,
            I => \N__26476\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__26479\,
            I => \N__26473\
        );

    \I__6277\ : Span4Mux_h
    port map (
            O => \N__26476\,
            I => \N__26470\
        );

    \I__6276\ : Span4Mux_v
    port map (
            O => \N__26473\,
            I => \N__26467\
        );

    \I__6275\ : Span4Mux_h
    port map (
            O => \N__26470\,
            I => \N__26464\
        );

    \I__6274\ : Span4Mux_h
    port map (
            O => \N__26467\,
            I => \N__26461\
        );

    \I__6273\ : Odrv4
    port map (
            O => \N__26464\,
            I => \tok.n15_adj_662\
        );

    \I__6272\ : Odrv4
    port map (
            O => \N__26461\,
            I => \tok.n15_adj_662\
        );

    \I__6271\ : CascadeMux
    port map (
            O => \N__26456\,
            I => \N__26452\
        );

    \I__6270\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26449\
        );

    \I__6269\ : InMux
    port map (
            O => \N__26452\,
            I => \N__26446\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__26449\,
            I => \tok.n4464\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__26446\,
            I => \tok.n4464\
        );

    \I__6266\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26438\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__26438\,
            I => \tok.n4573\
        );

    \I__6264\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26431\
        );

    \I__6263\ : CascadeMux
    port map (
            O => \N__26434\,
            I => \N__26428\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__26431\,
            I => \N__26425\
        );

    \I__6261\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26422\
        );

    \I__6260\ : Odrv12
    port map (
            O => \N__26425\,
            I => \tok.n9_adj_645\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__26422\,
            I => \tok.n9_adj_645\
        );

    \I__6258\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26411\
        );

    \I__6257\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26411\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__26411\,
            I => \N__26407\
        );

    \I__6255\ : InMux
    port map (
            O => \N__26410\,
            I => \N__26404\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__26407\,
            I => \N__26401\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__26404\,
            I => \N__26398\
        );

    \I__6252\ : Span4Mux_h
    port map (
            O => \N__26401\,
            I => \N__26394\
        );

    \I__6251\ : Span4Mux_v
    port map (
            O => \N__26398\,
            I => \N__26391\
        );

    \I__6250\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26388\
        );

    \I__6249\ : Odrv4
    port map (
            O => \N__26394\,
            I => \tok.n11\
        );

    \I__6248\ : Odrv4
    port map (
            O => \N__26391\,
            I => \tok.n11\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__26388\,
            I => \tok.n11\
        );

    \I__6246\ : CascadeMux
    port map (
            O => \N__26381\,
            I => \tok.n6_cascade_\
        );

    \I__6245\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26375\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__26375\,
            I => \N__26371\
        );

    \I__6243\ : InMux
    port map (
            O => \N__26374\,
            I => \N__26368\
        );

    \I__6242\ : Odrv12
    port map (
            O => \N__26371\,
            I => \tok.C_stk.tail_2\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__26368\,
            I => \tok.C_stk.tail_2\
        );

    \I__6240\ : CascadeMux
    port map (
            O => \N__26363\,
            I => \tok.C_stk.n4876_cascade_\
        );

    \I__6239\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26353\
        );

    \I__6238\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26353\
        );

    \I__6237\ : CascadeMux
    port map (
            O => \N__26358\,
            I => \N__26349\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__26353\,
            I => \N__26342\
        );

    \I__6235\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26337\
        );

    \I__6234\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26337\
        );

    \I__6233\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26332\
        );

    \I__6232\ : InMux
    port map (
            O => \N__26347\,
            I => \N__26332\
        );

    \I__6231\ : InMux
    port map (
            O => \N__26346\,
            I => \N__26325\
        );

    \I__6230\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26325\
        );

    \I__6229\ : Span4Mux_s3_v
    port map (
            O => \N__26342\,
            I => \N__26317\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__26337\,
            I => \N__26317\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__26332\,
            I => \N__26314\
        );

    \I__6226\ : InMux
    port map (
            O => \N__26331\,
            I => \N__26309\
        );

    \I__6225\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26309\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__26325\,
            I => \N__26306\
        );

    \I__6223\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26296\
        );

    \I__6222\ : InMux
    port map (
            O => \N__26323\,
            I => \N__26296\
        );

    \I__6221\ : InMux
    port map (
            O => \N__26322\,
            I => \N__26296\
        );

    \I__6220\ : Span4Mux_v
    port map (
            O => \N__26317\,
            I => \N__26291\
        );

    \I__6219\ : Span4Mux_s3_v
    port map (
            O => \N__26314\,
            I => \N__26291\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__26309\,
            I => \N__26286\
        );

    \I__6217\ : Span4Mux_h
    port map (
            O => \N__26306\,
            I => \N__26286\
        );

    \I__6216\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26279\
        );

    \I__6215\ : InMux
    port map (
            O => \N__26304\,
            I => \N__26279\
        );

    \I__6214\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26279\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__26296\,
            I => \tok.C_stk.n600\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__26291\,
            I => \tok.C_stk.n600\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__26286\,
            I => \tok.C_stk.n600\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__26279\,
            I => \tok.C_stk.n600\
        );

    \I__6209\ : ClkMux
    port map (
            O => \N__26270\,
            I => \N__26042\
        );

    \I__6208\ : ClkMux
    port map (
            O => \N__26269\,
            I => \N__26042\
        );

    \I__6207\ : ClkMux
    port map (
            O => \N__26268\,
            I => \N__26042\
        );

    \I__6206\ : ClkMux
    port map (
            O => \N__26267\,
            I => \N__26042\
        );

    \I__6205\ : ClkMux
    port map (
            O => \N__26266\,
            I => \N__26042\
        );

    \I__6204\ : ClkMux
    port map (
            O => \N__26265\,
            I => \N__26042\
        );

    \I__6203\ : ClkMux
    port map (
            O => \N__26264\,
            I => \N__26042\
        );

    \I__6202\ : ClkMux
    port map (
            O => \N__26263\,
            I => \N__26042\
        );

    \I__6201\ : ClkMux
    port map (
            O => \N__26262\,
            I => \N__26042\
        );

    \I__6200\ : ClkMux
    port map (
            O => \N__26261\,
            I => \N__26042\
        );

    \I__6199\ : ClkMux
    port map (
            O => \N__26260\,
            I => \N__26042\
        );

    \I__6198\ : ClkMux
    port map (
            O => \N__26259\,
            I => \N__26042\
        );

    \I__6197\ : ClkMux
    port map (
            O => \N__26258\,
            I => \N__26042\
        );

    \I__6196\ : ClkMux
    port map (
            O => \N__26257\,
            I => \N__26042\
        );

    \I__6195\ : ClkMux
    port map (
            O => \N__26256\,
            I => \N__26042\
        );

    \I__6194\ : ClkMux
    port map (
            O => \N__26255\,
            I => \N__26042\
        );

    \I__6193\ : ClkMux
    port map (
            O => \N__26254\,
            I => \N__26042\
        );

    \I__6192\ : ClkMux
    port map (
            O => \N__26253\,
            I => \N__26042\
        );

    \I__6191\ : ClkMux
    port map (
            O => \N__26252\,
            I => \N__26042\
        );

    \I__6190\ : ClkMux
    port map (
            O => \N__26251\,
            I => \N__26042\
        );

    \I__6189\ : ClkMux
    port map (
            O => \N__26250\,
            I => \N__26042\
        );

    \I__6188\ : ClkMux
    port map (
            O => \N__26249\,
            I => \N__26042\
        );

    \I__6187\ : ClkMux
    port map (
            O => \N__26248\,
            I => \N__26042\
        );

    \I__6186\ : ClkMux
    port map (
            O => \N__26247\,
            I => \N__26042\
        );

    \I__6185\ : ClkMux
    port map (
            O => \N__26246\,
            I => \N__26042\
        );

    \I__6184\ : ClkMux
    port map (
            O => \N__26245\,
            I => \N__26042\
        );

    \I__6183\ : ClkMux
    port map (
            O => \N__26244\,
            I => \N__26042\
        );

    \I__6182\ : ClkMux
    port map (
            O => \N__26243\,
            I => \N__26042\
        );

    \I__6181\ : ClkMux
    port map (
            O => \N__26242\,
            I => \N__26042\
        );

    \I__6180\ : ClkMux
    port map (
            O => \N__26241\,
            I => \N__26042\
        );

    \I__6179\ : ClkMux
    port map (
            O => \N__26240\,
            I => \N__26042\
        );

    \I__6178\ : ClkMux
    port map (
            O => \N__26239\,
            I => \N__26042\
        );

    \I__6177\ : ClkMux
    port map (
            O => \N__26238\,
            I => \N__26042\
        );

    \I__6176\ : ClkMux
    port map (
            O => \N__26237\,
            I => \N__26042\
        );

    \I__6175\ : ClkMux
    port map (
            O => \N__26236\,
            I => \N__26042\
        );

    \I__6174\ : ClkMux
    port map (
            O => \N__26235\,
            I => \N__26042\
        );

    \I__6173\ : ClkMux
    port map (
            O => \N__26234\,
            I => \N__26042\
        );

    \I__6172\ : ClkMux
    port map (
            O => \N__26233\,
            I => \N__26042\
        );

    \I__6171\ : ClkMux
    port map (
            O => \N__26232\,
            I => \N__26042\
        );

    \I__6170\ : ClkMux
    port map (
            O => \N__26231\,
            I => \N__26042\
        );

    \I__6169\ : ClkMux
    port map (
            O => \N__26230\,
            I => \N__26042\
        );

    \I__6168\ : ClkMux
    port map (
            O => \N__26229\,
            I => \N__26042\
        );

    \I__6167\ : ClkMux
    port map (
            O => \N__26228\,
            I => \N__26042\
        );

    \I__6166\ : ClkMux
    port map (
            O => \N__26227\,
            I => \N__26042\
        );

    \I__6165\ : ClkMux
    port map (
            O => \N__26226\,
            I => \N__26042\
        );

    \I__6164\ : ClkMux
    port map (
            O => \N__26225\,
            I => \N__26042\
        );

    \I__6163\ : ClkMux
    port map (
            O => \N__26224\,
            I => \N__26042\
        );

    \I__6162\ : ClkMux
    port map (
            O => \N__26223\,
            I => \N__26042\
        );

    \I__6161\ : ClkMux
    port map (
            O => \N__26222\,
            I => \N__26042\
        );

    \I__6160\ : ClkMux
    port map (
            O => \N__26221\,
            I => \N__26042\
        );

    \I__6159\ : ClkMux
    port map (
            O => \N__26220\,
            I => \N__26042\
        );

    \I__6158\ : ClkMux
    port map (
            O => \N__26219\,
            I => \N__26042\
        );

    \I__6157\ : ClkMux
    port map (
            O => \N__26218\,
            I => \N__26042\
        );

    \I__6156\ : ClkMux
    port map (
            O => \N__26217\,
            I => \N__26042\
        );

    \I__6155\ : ClkMux
    port map (
            O => \N__26216\,
            I => \N__26042\
        );

    \I__6154\ : ClkMux
    port map (
            O => \N__26215\,
            I => \N__26042\
        );

    \I__6153\ : ClkMux
    port map (
            O => \N__26214\,
            I => \N__26042\
        );

    \I__6152\ : ClkMux
    port map (
            O => \N__26213\,
            I => \N__26042\
        );

    \I__6151\ : ClkMux
    port map (
            O => \N__26212\,
            I => \N__26042\
        );

    \I__6150\ : ClkMux
    port map (
            O => \N__26211\,
            I => \N__26042\
        );

    \I__6149\ : ClkMux
    port map (
            O => \N__26210\,
            I => \N__26042\
        );

    \I__6148\ : ClkMux
    port map (
            O => \N__26209\,
            I => \N__26042\
        );

    \I__6147\ : ClkMux
    port map (
            O => \N__26208\,
            I => \N__26042\
        );

    \I__6146\ : ClkMux
    port map (
            O => \N__26207\,
            I => \N__26042\
        );

    \I__6145\ : ClkMux
    port map (
            O => \N__26206\,
            I => \N__26042\
        );

    \I__6144\ : ClkMux
    port map (
            O => \N__26205\,
            I => \N__26042\
        );

    \I__6143\ : ClkMux
    port map (
            O => \N__26204\,
            I => \N__26042\
        );

    \I__6142\ : ClkMux
    port map (
            O => \N__26203\,
            I => \N__26042\
        );

    \I__6141\ : ClkMux
    port map (
            O => \N__26202\,
            I => \N__26042\
        );

    \I__6140\ : ClkMux
    port map (
            O => \N__26201\,
            I => \N__26042\
        );

    \I__6139\ : ClkMux
    port map (
            O => \N__26200\,
            I => \N__26042\
        );

    \I__6138\ : ClkMux
    port map (
            O => \N__26199\,
            I => \N__26042\
        );

    \I__6137\ : ClkMux
    port map (
            O => \N__26198\,
            I => \N__26042\
        );

    \I__6136\ : ClkMux
    port map (
            O => \N__26197\,
            I => \N__26042\
        );

    \I__6135\ : ClkMux
    port map (
            O => \N__26196\,
            I => \N__26042\
        );

    \I__6134\ : ClkMux
    port map (
            O => \N__26195\,
            I => \N__26042\
        );

    \I__6133\ : GlobalMux
    port map (
            O => \N__26042\,
            I => \N__26039\
        );

    \I__6132\ : DummyBuf
    port map (
            O => \N__26039\,
            I => clk
        );

    \I__6131\ : CascadeMux
    port map (
            O => \N__26036\,
            I => \N__26033\
        );

    \I__6130\ : InMux
    port map (
            O => \N__26033\,
            I => \N__26027\
        );

    \I__6129\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26024\
        );

    \I__6128\ : InMux
    port map (
            O => \N__26031\,
            I => \N__26019\
        );

    \I__6127\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26019\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__26027\,
            I => \N__26016\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__26024\,
            I => \N__26011\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__26019\,
            I => \N__26011\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__26016\,
            I => \N__26008\
        );

    \I__6122\ : Span4Mux_s3_h
    port map (
            O => \N__26011\,
            I => \N__26005\
        );

    \I__6121\ : Odrv4
    port map (
            O => \N__26008\,
            I => \tok.tc_plus_1_2\
        );

    \I__6120\ : Odrv4
    port map (
            O => \N__26005\,
            I => \tok.tc_plus_1_2\
        );

    \I__6119\ : InMux
    port map (
            O => \N__26000\,
            I => \N__25997\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__25997\,
            I => \N__25991\
        );

    \I__6117\ : InMux
    port map (
            O => \N__25996\,
            I => \N__25987\
        );

    \I__6116\ : InMux
    port map (
            O => \N__25995\,
            I => \N__25984\
        );

    \I__6115\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25980\
        );

    \I__6114\ : Span4Mux_v
    port map (
            O => \N__25991\,
            I => \N__25975\
        );

    \I__6113\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25972\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__25987\,
            I => \N__25969\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__25984\,
            I => \N__25966\
        );

    \I__6110\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25963\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__25980\,
            I => \N__25960\
        );

    \I__6108\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25957\
        );

    \I__6107\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25954\
        );

    \I__6106\ : Span4Mux_h
    port map (
            O => \N__25975\,
            I => \N__25949\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__25972\,
            I => \N__25949\
        );

    \I__6104\ : Span4Mux_h
    port map (
            O => \N__25969\,
            I => \N__25946\
        );

    \I__6103\ : Span4Mux_h
    port map (
            O => \N__25966\,
            I => \N__25943\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__25963\,
            I => \N__25938\
        );

    \I__6101\ : Span4Mux_v
    port map (
            O => \N__25960\,
            I => \N__25938\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__25957\,
            I => \N__25933\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__25954\,
            I => \N__25933\
        );

    \I__6098\ : Odrv4
    port map (
            O => \N__25949\,
            I => \tok.tc__7__N_134\
        );

    \I__6097\ : Odrv4
    port map (
            O => \N__25946\,
            I => \tok.tc__7__N_134\
        );

    \I__6096\ : Odrv4
    port map (
            O => \N__25943\,
            I => \tok.tc__7__N_134\
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__25938\,
            I => \tok.tc__7__N_134\
        );

    \I__6094\ : Odrv12
    port map (
            O => \N__25933\,
            I => \tok.tc__7__N_134\
        );

    \I__6093\ : CascadeMux
    port map (
            O => \N__25922\,
            I => \tok.ram.n4711_cascade_\
        );

    \I__6092\ : CascadeMux
    port map (
            O => \N__25919\,
            I => \tok.n1_adj_724_cascade_\
        );

    \I__6091\ : InMux
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__25913\,
            I => \tok.n13_adj_725\
        );

    \I__6089\ : InMux
    port map (
            O => \N__25910\,
            I => \N__25905\
        );

    \I__6088\ : InMux
    port map (
            O => \N__25909\,
            I => \N__25900\
        );

    \I__6087\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25900\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__25905\,
            I => \N__25894\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__25900\,
            I => \N__25891\
        );

    \I__6084\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25888\
        );

    \I__6083\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25885\
        );

    \I__6082\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25881\
        );

    \I__6081\ : Span4Mux_s1_h
    port map (
            O => \N__25894\,
            I => \N__25874\
        );

    \I__6080\ : Span4Mux_v
    port map (
            O => \N__25891\,
            I => \N__25874\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__25888\,
            I => \N__25874\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__25885\,
            I => \N__25869\
        );

    \I__6077\ : InMux
    port map (
            O => \N__25884\,
            I => \N__25866\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__25881\,
            I => \N__25861\
        );

    \I__6075\ : Span4Mux_h
    port map (
            O => \N__25874\,
            I => \N__25861\
        );

    \I__6074\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25858\
        );

    \I__6073\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25855\
        );

    \I__6072\ : Odrv4
    port map (
            O => \N__25869\,
            I => \tok.n101_adj_776\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__25866\,
            I => \tok.n101_adj_776\
        );

    \I__6070\ : Odrv4
    port map (
            O => \N__25861\,
            I => \tok.n101_adj_776\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__25858\,
            I => \tok.n101_adj_776\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__25855\,
            I => \tok.n101_adj_776\
        );

    \I__6067\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25841\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__25841\,
            I => \tok.ram.n4708\
        );

    \I__6065\ : InMux
    port map (
            O => \N__25838\,
            I => \N__25835\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__25835\,
            I => \tok.n1_adj_736\
        );

    \I__6063\ : InMux
    port map (
            O => \N__25832\,
            I => \N__25829\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__25829\,
            I => \tok.n5_adj_737\
        );

    \I__6061\ : InMux
    port map (
            O => \N__25826\,
            I => \N__25822\
        );

    \I__6060\ : CascadeMux
    port map (
            O => \N__25825\,
            I => \N__25817\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__25822\,
            I => \N__25813\
        );

    \I__6058\ : InMux
    port map (
            O => \N__25821\,
            I => \N__25806\
        );

    \I__6057\ : InMux
    port map (
            O => \N__25820\,
            I => \N__25806\
        );

    \I__6056\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25806\
        );

    \I__6055\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25803\
        );

    \I__6054\ : Odrv4
    port map (
            O => \N__25813\,
            I => \tok.c_stk_r_2\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__25806\,
            I => \tok.c_stk_r_2\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__25803\,
            I => \tok.c_stk_r_2\
        );

    \I__6051\ : CascadeMux
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__6050\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25789\
        );

    \I__6049\ : InMux
    port map (
            O => \N__25792\,
            I => \N__25786\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__25789\,
            I => \N__25783\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__25786\,
            I => \N__25780\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__25783\,
            I => \N__25777\
        );

    \I__6045\ : Span4Mux_v
    port map (
            O => \N__25780\,
            I => \N__25774\
        );

    \I__6044\ : Span4Mux_h
    port map (
            O => \N__25777\,
            I => \N__25771\
        );

    \I__6043\ : Span4Mux_h
    port map (
            O => \N__25774\,
            I => \N__25768\
        );

    \I__6042\ : Span4Mux_h
    port map (
            O => \N__25771\,
            I => \N__25765\
        );

    \I__6041\ : Odrv4
    port map (
            O => \N__25768\,
            I => \tok.table_rd_2\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__25765\,
            I => \tok.table_rd_2\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__25760\,
            I => \tok.n83_adj_721_cascade_\
        );

    \I__6038\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__25754\,
            I => \tok.n4692\
        );

    \I__6036\ : InMux
    port map (
            O => \N__25751\,
            I => \N__25748\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__25748\,
            I => \N__25744\
        );

    \I__6034\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25741\
        );

    \I__6033\ : Span4Mux_s2_v
    port map (
            O => \N__25744\,
            I => \N__25738\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__25741\,
            I => \tok.tail_10\
        );

    \I__6031\ : Odrv4
    port map (
            O => \N__25738\,
            I => \tok.tail_10\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__25733\,
            I => \N__25701\
        );

    \I__6029\ : CascadeMux
    port map (
            O => \N__25732\,
            I => \N__25698\
        );

    \I__6028\ : InMux
    port map (
            O => \N__25731\,
            I => \N__25678\
        );

    \I__6027\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25678\
        );

    \I__6026\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25678\
        );

    \I__6025\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25678\
        );

    \I__6024\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25678\
        );

    \I__6023\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25678\
        );

    \I__6022\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25678\
        );

    \I__6021\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25678\
        );

    \I__6020\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25661\
        );

    \I__6019\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25661\
        );

    \I__6018\ : InMux
    port map (
            O => \N__25721\,
            I => \N__25661\
        );

    \I__6017\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25661\
        );

    \I__6016\ : InMux
    port map (
            O => \N__25719\,
            I => \N__25661\
        );

    \I__6015\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25661\
        );

    \I__6014\ : InMux
    port map (
            O => \N__25717\,
            I => \N__25661\
        );

    \I__6013\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25661\
        );

    \I__6012\ : InMux
    port map (
            O => \N__25715\,
            I => \N__25643\
        );

    \I__6011\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25643\
        );

    \I__6010\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25643\
        );

    \I__6009\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25643\
        );

    \I__6008\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25643\
        );

    \I__6007\ : InMux
    port map (
            O => \N__25710\,
            I => \N__25643\
        );

    \I__6006\ : InMux
    port map (
            O => \N__25709\,
            I => \N__25643\
        );

    \I__6005\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25643\
        );

    \I__6004\ : CascadeMux
    port map (
            O => \N__25707\,
            I => \N__25632\
        );

    \I__6003\ : CascadeMux
    port map (
            O => \N__25706\,
            I => \N__25629\
        );

    \I__6002\ : CascadeMux
    port map (
            O => \N__25705\,
            I => \N__25626\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__25704\,
            I => \N__25623\
        );

    \I__6000\ : InMux
    port map (
            O => \N__25701\,
            I => \N__25608\
        );

    \I__5999\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25608\
        );

    \I__5998\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25608\
        );

    \I__5997\ : InMux
    port map (
            O => \N__25696\,
            I => \N__25608\
        );

    \I__5996\ : InMux
    port map (
            O => \N__25695\,
            I => \N__25608\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__25678\,
            I => \N__25605\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__25661\,
            I => \N__25602\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__25660\,
            I => \N__25599\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__25643\,
            I => \N__25578\
        );

    \I__5991\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25561\
        );

    \I__5990\ : InMux
    port map (
            O => \N__25641\,
            I => \N__25561\
        );

    \I__5989\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25561\
        );

    \I__5988\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25561\
        );

    \I__5987\ : InMux
    port map (
            O => \N__25638\,
            I => \N__25561\
        );

    \I__5986\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25561\
        );

    \I__5985\ : InMux
    port map (
            O => \N__25636\,
            I => \N__25561\
        );

    \I__5984\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25561\
        );

    \I__5983\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25544\
        );

    \I__5982\ : InMux
    port map (
            O => \N__25629\,
            I => \N__25544\
        );

    \I__5981\ : InMux
    port map (
            O => \N__25626\,
            I => \N__25544\
        );

    \I__5980\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25544\
        );

    \I__5979\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25544\
        );

    \I__5978\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25544\
        );

    \I__5977\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25544\
        );

    \I__5976\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25544\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__25608\,
            I => \N__25537\
        );

    \I__5974\ : Span4Mux_s3_v
    port map (
            O => \N__25605\,
            I => \N__25537\
        );

    \I__5973\ : Span4Mux_s1_h
    port map (
            O => \N__25602\,
            I => \N__25537\
        );

    \I__5972\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25530\
        );

    \I__5971\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25530\
        );

    \I__5970\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25530\
        );

    \I__5969\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25513\
        );

    \I__5968\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25513\
        );

    \I__5967\ : InMux
    port map (
            O => \N__25594\,
            I => \N__25513\
        );

    \I__5966\ : InMux
    port map (
            O => \N__25593\,
            I => \N__25513\
        );

    \I__5965\ : InMux
    port map (
            O => \N__25592\,
            I => \N__25513\
        );

    \I__5964\ : InMux
    port map (
            O => \N__25591\,
            I => \N__25513\
        );

    \I__5963\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25513\
        );

    \I__5962\ : InMux
    port map (
            O => \N__25589\,
            I => \N__25513\
        );

    \I__5961\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25496\
        );

    \I__5960\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25496\
        );

    \I__5959\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25496\
        );

    \I__5958\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25496\
        );

    \I__5957\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25496\
        );

    \I__5956\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25496\
        );

    \I__5955\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25496\
        );

    \I__5954\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25496\
        );

    \I__5953\ : Span4Mux_s2_v
    port map (
            O => \N__25578\,
            I => \N__25493\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__25561\,
            I => \N__25488\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__25544\,
            I => \N__25488\
        );

    \I__5950\ : Span4Mux_h
    port map (
            O => \N__25537\,
            I => \N__25485\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__25530\,
            I => \tok.C_stk_delta_1\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__25513\,
            I => \tok.C_stk_delta_1\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__25496\,
            I => \tok.C_stk_delta_1\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__25493\,
            I => \tok.C_stk_delta_1\
        );

    \I__5945\ : Odrv12
    port map (
            O => \N__25488\,
            I => \tok.C_stk_delta_1\
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__25485\,
            I => \tok.C_stk_delta_1\
        );

    \I__5943\ : CEMux
    port map (
            O => \N__25472\,
            I => \N__25468\
        );

    \I__5942\ : CEMux
    port map (
            O => \N__25471\,
            I => \N__25455\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__25468\,
            I => \N__25452\
        );

    \I__5940\ : CEMux
    port map (
            O => \N__25467\,
            I => \N__25449\
        );

    \I__5939\ : CEMux
    port map (
            O => \N__25466\,
            I => \N__25446\
        );

    \I__5938\ : CEMux
    port map (
            O => \N__25465\,
            I => \N__25443\
        );

    \I__5937\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25428\
        );

    \I__5936\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25428\
        );

    \I__5935\ : InMux
    port map (
            O => \N__25462\,
            I => \N__25428\
        );

    \I__5934\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25428\
        );

    \I__5933\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25428\
        );

    \I__5932\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25428\
        );

    \I__5931\ : InMux
    port map (
            O => \N__25458\,
            I => \N__25428\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__25455\,
            I => \N__25423\
        );

    \I__5929\ : Span4Mux_s2_h
    port map (
            O => \N__25452\,
            I => \N__25417\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__25449\,
            I => \N__25414\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__25446\,
            I => \N__25411\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__25443\,
            I => \N__25408\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__25428\,
            I => \N__25405\
        );

    \I__5924\ : CEMux
    port map (
            O => \N__25427\,
            I => \N__25402\
        );

    \I__5923\ : CEMux
    port map (
            O => \N__25426\,
            I => \N__25399\
        );

    \I__5922\ : Span4Mux_h
    port map (
            O => \N__25423\,
            I => \N__25396\
        );

    \I__5921\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25389\
        );

    \I__5920\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25389\
        );

    \I__5919\ : InMux
    port map (
            O => \N__25420\,
            I => \N__25389\
        );

    \I__5918\ : Span4Mux_h
    port map (
            O => \N__25417\,
            I => \N__25386\
        );

    \I__5917\ : Span4Mux_s2_h
    port map (
            O => \N__25414\,
            I => \N__25377\
        );

    \I__5916\ : Span4Mux_s2_h
    port map (
            O => \N__25411\,
            I => \N__25377\
        );

    \I__5915\ : Span4Mux_s2_v
    port map (
            O => \N__25408\,
            I => \N__25377\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__25405\,
            I => \N__25377\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__25402\,
            I => \tok.rd_7__N_374\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__25399\,
            I => \tok.rd_7__N_374\
        );

    \I__5911\ : Odrv4
    port map (
            O => \N__25396\,
            I => \tok.rd_7__N_374\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__25389\,
            I => \tok.rd_7__N_374\
        );

    \I__5909\ : Odrv4
    port map (
            O => \N__25386\,
            I => \tok.rd_7__N_374\
        );

    \I__5908\ : Odrv4
    port map (
            O => \N__25377\,
            I => \tok.rd_7__N_374\
        );

    \I__5907\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25360\
        );

    \I__5906\ : InMux
    port map (
            O => \N__25363\,
            I => \N__25356\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__25360\,
            I => \N__25353\
        );

    \I__5904\ : InMux
    port map (
            O => \N__25359\,
            I => \N__25349\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__25356\,
            I => \N__25344\
        );

    \I__5902\ : Span4Mux_v
    port map (
            O => \N__25353\,
            I => \N__25344\
        );

    \I__5901\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25341\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__25349\,
            I => \c_stk_w_7_N_18_4\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__25344\,
            I => \c_stk_w_7_N_18_4\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__25341\,
            I => \c_stk_w_7_N_18_4\
        );

    \I__5897\ : InMux
    port map (
            O => \N__25334\,
            I => \N__25331\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__5895\ : Span12Mux_v
    port map (
            O => \N__25328\,
            I => \N__25324\
        );

    \I__5894\ : InMux
    port map (
            O => \N__25327\,
            I => \N__25321\
        );

    \I__5893\ : Odrv12
    port map (
            O => \N__25324\,
            I => \tok.C_stk.tail_4\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__25321\,
            I => \tok.C_stk.tail_4\
        );

    \I__5891\ : CascadeMux
    port map (
            O => \N__25316\,
            I => \tok.C_stk.n4888_cascade_\
        );

    \I__5890\ : CascadeMux
    port map (
            O => \N__25313\,
            I => \tok.ram.n4705_cascade_\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__25310\,
            I => \tok.n1_adj_745_cascade_\
        );

    \I__5888\ : CascadeMux
    port map (
            O => \N__25307\,
            I => \N__25304\
        );

    \I__5887\ : InMux
    port map (
            O => \N__25304\,
            I => \N__25301\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__5885\ : Span4Mux_v
    port map (
            O => \N__25298\,
            I => \N__25292\
        );

    \I__5884\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25285\
        );

    \I__5883\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25285\
        );

    \I__5882\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25285\
        );

    \I__5881\ : Span4Mux_h
    port map (
            O => \N__25292\,
            I => \N__25280\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__25285\,
            I => \N__25280\
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__25280\,
            I => \tok.tc_plus_1_4\
        );

    \I__5878\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25272\
        );

    \I__5877\ : CascadeMux
    port map (
            O => \N__25276\,
            I => \N__25269\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__25275\,
            I => \N__25266\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__25272\,
            I => \N__25262\
        );

    \I__5874\ : InMux
    port map (
            O => \N__25269\,
            I => \N__25252\
        );

    \I__5873\ : InMux
    port map (
            O => \N__25266\,
            I => \N__25252\
        );

    \I__5872\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25252\
        );

    \I__5871\ : Span4Mux_s2_h
    port map (
            O => \N__25262\,
            I => \N__25248\
        );

    \I__5870\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25245\
        );

    \I__5869\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25242\
        );

    \I__5868\ : CascadeMux
    port map (
            O => \N__25259\,
            I => \N__25239\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__25252\,
            I => \N__25236\
        );

    \I__5866\ : InMux
    port map (
            O => \N__25251\,
            I => \N__25233\
        );

    \I__5865\ : Span4Mux_h
    port map (
            O => \N__25248\,
            I => \N__25230\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__25245\,
            I => \N__25225\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__25242\,
            I => \N__25225\
        );

    \I__5862\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25222\
        );

    \I__5861\ : Span4Mux_v
    port map (
            O => \N__25236\,
            I => \N__25217\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__25233\,
            I => \N__25217\
        );

    \I__5859\ : Odrv4
    port map (
            O => \N__25230\,
            I => \tok.n802\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__25225\,
            I => \tok.n802\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__25222\,
            I => \tok.n802\
        );

    \I__5856\ : Odrv4
    port map (
            O => \N__25217\,
            I => \tok.n802\
        );

    \I__5855\ : CascadeMux
    port map (
            O => \N__25208\,
            I => \tok.n13_adj_746_cascade_\
        );

    \I__5854\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25195\
        );

    \I__5853\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25195\
        );

    \I__5852\ : InMux
    port map (
            O => \N__25203\,
            I => \N__25195\
        );

    \I__5851\ : InMux
    port map (
            O => \N__25202\,
            I => \N__25192\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__25195\,
            I => \N__25184\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__25192\,
            I => \N__25184\
        );

    \I__5848\ : InMux
    port map (
            O => \N__25191\,
            I => \N__25180\
        );

    \I__5847\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25177\
        );

    \I__5846\ : InMux
    port map (
            O => \N__25189\,
            I => \N__25174\
        );

    \I__5845\ : Span4Mux_v
    port map (
            O => \N__25184\,
            I => \N__25171\
        );

    \I__5844\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25168\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__25180\,
            I => \N__25165\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25160\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__25174\,
            I => \N__25160\
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__25171\,
            I => \tok.n86\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__25168\,
            I => \tok.n86\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__25165\,
            I => \tok.n86\
        );

    \I__5837\ : Odrv12
    port map (
            O => \N__25160\,
            I => \tok.n86\
        );

    \I__5836\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25148\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__25148\,
            I => \N__25145\
        );

    \I__5834\ : Span4Mux_v
    port map (
            O => \N__25145\,
            I => \N__25141\
        );

    \I__5833\ : InMux
    port map (
            O => \N__25144\,
            I => \N__25138\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__25141\,
            I => n10
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__25138\,
            I => n10
        );

    \I__5830\ : InMux
    port map (
            O => \N__25133\,
            I => \N__25129\
        );

    \I__5829\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25126\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__25129\,
            I => \tok.C_stk.tail_3\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__25126\,
            I => \tok.C_stk.tail_3\
        );

    \I__5826\ : CascadeMux
    port map (
            O => \N__25121\,
            I => \N__25118\
        );

    \I__5825\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25115\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__25115\,
            I => \tok.C_stk.n4882\
        );

    \I__5823\ : CascadeMux
    port map (
            O => \N__25112\,
            I => \N__25108\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__25111\,
            I => \N__25102\
        );

    \I__5821\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25098\
        );

    \I__5820\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25095\
        );

    \I__5819\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25092\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__25105\,
            I => \N__25089\
        );

    \I__5817\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25086\
        );

    \I__5816\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25083\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__25098\,
            I => \N__25078\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__25095\,
            I => \N__25078\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__25092\,
            I => \N__25075\
        );

    \I__5812\ : InMux
    port map (
            O => \N__25089\,
            I => \N__25070\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__25086\,
            I => \N__25067\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__25083\,
            I => \N__25062\
        );

    \I__5809\ : Span4Mux_v
    port map (
            O => \N__25078\,
            I => \N__25062\
        );

    \I__5808\ : Span4Mux_s3_v
    port map (
            O => \N__25075\,
            I => \N__25059\
        );

    \I__5807\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25054\
        );

    \I__5806\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25054\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__25070\,
            I => \tok.n602\
        );

    \I__5804\ : Odrv4
    port map (
            O => \N__25067\,
            I => \tok.n602\
        );

    \I__5803\ : Odrv4
    port map (
            O => \N__25062\,
            I => \tok.n602\
        );

    \I__5802\ : Odrv4
    port map (
            O => \N__25059\,
            I => \tok.n602\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__25054\,
            I => \tok.n602\
        );

    \I__5800\ : InMux
    port map (
            O => \N__25043\,
            I => \N__25038\
        );

    \I__5799\ : InMux
    port map (
            O => \N__25042\,
            I => \N__25035\
        );

    \I__5798\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25031\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__25038\,
            I => \N__25026\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__25035\,
            I => \N__25026\
        );

    \I__5795\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25023\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__25031\,
            I => \c_stk_w_7_N_18_2\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__25026\,
            I => \c_stk_w_7_N_18_2\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__25023\,
            I => \c_stk_w_7_N_18_2\
        );

    \I__5791\ : InMux
    port map (
            O => \N__25016\,
            I => \N__25012\
        );

    \I__5790\ : InMux
    port map (
            O => \N__25015\,
            I => \N__25009\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__25012\,
            I => \tok.tail_61\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__25009\,
            I => \tok.tail_61\
        );

    \I__5787\ : InMux
    port map (
            O => \N__25004\,
            I => \N__24998\
        );

    \I__5786\ : InMux
    port map (
            O => \N__25003\,
            I => \N__24998\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__24998\,
            I => \tok.tail_45\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__24995\,
            I => \N__24992\
        );

    \I__5783\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__24989\,
            I => \N__24986\
        );

    \I__5781\ : Span4Mux_h
    port map (
            O => \N__24986\,
            I => \N__24982\
        );

    \I__5780\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24979\
        );

    \I__5779\ : Odrv4
    port map (
            O => \N__24982\,
            I => \tok.tail_53\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__24979\,
            I => \tok.tail_53\
        );

    \I__5777\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24970\
        );

    \I__5776\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24967\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__24970\,
            I => \tok.C_stk.tail_22\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__24967\,
            I => \tok.C_stk.tail_22\
        );

    \I__5773\ : InMux
    port map (
            O => \N__24962\,
            I => \N__24959\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__24959\,
            I => \N__24956\
        );

    \I__5771\ : Span4Mux_h
    port map (
            O => \N__24956\,
            I => \N__24953\
        );

    \I__5770\ : Span4Mux_s2_h
    port map (
            O => \N__24953\,
            I => \N__24949\
        );

    \I__5769\ : InMux
    port map (
            O => \N__24952\,
            I => \N__24946\
        );

    \I__5768\ : Odrv4
    port map (
            O => \N__24949\,
            I => \tok.C_stk.tail_6\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__24946\,
            I => \tok.C_stk.tail_6\
        );

    \I__5766\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24935\
        );

    \I__5765\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24935\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__24935\,
            I => \tok.tail_14\
        );

    \I__5763\ : InMux
    port map (
            O => \N__24932\,
            I => \N__24926\
        );

    \I__5762\ : InMux
    port map (
            O => \N__24931\,
            I => \N__24926\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__24926\,
            I => \tok.tail_11\
        );

    \I__5760\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24917\
        );

    \I__5759\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24917\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__24917\,
            I => \tok.C_stk.tail_19\
        );

    \I__5757\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24908\
        );

    \I__5756\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24908\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__24908\,
            I => \tok.tail_27\
        );

    \I__5754\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24899\
        );

    \I__5753\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24899\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__24899\,
            I => \tok.C_stk.tail_35\
        );

    \I__5751\ : InMux
    port map (
            O => \N__24896\,
            I => \N__24892\
        );

    \I__5750\ : InMux
    port map (
            O => \N__24895\,
            I => \N__24889\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__24892\,
            I => \tok.tail_59\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__24889\,
            I => \tok.tail_59\
        );

    \I__5747\ : InMux
    port map (
            O => \N__24884\,
            I => \N__24878\
        );

    \I__5746\ : InMux
    port map (
            O => \N__24883\,
            I => \N__24878\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__24878\,
            I => \tok.tail_43\
        );

    \I__5744\ : CascadeMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__5743\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24869\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__24869\,
            I => \N__24865\
        );

    \I__5741\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24862\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__24865\,
            I => \tok.tail_51\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__24862\,
            I => \tok.tail_51\
        );

    \I__5738\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24851\
        );

    \I__5737\ : CascadeMux
    port map (
            O => \N__24856\,
            I => \N__24848\
        );

    \I__5736\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24840\
        );

    \I__5735\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24836\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__24851\,
            I => \N__24832\
        );

    \I__5733\ : InMux
    port map (
            O => \N__24848\,
            I => \N__24829\
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__24847\,
            I => \N__24826\
        );

    \I__5731\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24823\
        );

    \I__5730\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24820\
        );

    \I__5729\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24815\
        );

    \I__5728\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24815\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__24840\,
            I => \N__24812\
        );

    \I__5726\ : InMux
    port map (
            O => \N__24839\,
            I => \N__24809\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__24836\,
            I => \N__24806\
        );

    \I__5724\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24803\
        );

    \I__5723\ : Span4Mux_s3_h
    port map (
            O => \N__24832\,
            I => \N__24798\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24798\
        );

    \I__5721\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24795\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__24823\,
            I => \N__24791\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__24820\,
            I => \N__24786\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24786\
        );

    \I__5717\ : Span4Mux_s3_h
    port map (
            O => \N__24812\,
            I => \N__24782\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24775\
        );

    \I__5715\ : Span4Mux_v
    port map (
            O => \N__24806\,
            I => \N__24775\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__24803\,
            I => \N__24775\
        );

    \I__5713\ : Span4Mux_v
    port map (
            O => \N__24798\,
            I => \N__24770\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__24795\,
            I => \N__24770\
        );

    \I__5711\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24767\
        );

    \I__5710\ : Span4Mux_h
    port map (
            O => \N__24791\,
            I => \N__24762\
        );

    \I__5709\ : Span4Mux_h
    port map (
            O => \N__24786\,
            I => \N__24762\
        );

    \I__5708\ : InMux
    port map (
            O => \N__24785\,
            I => \N__24759\
        );

    \I__5707\ : Span4Mux_h
    port map (
            O => \N__24782\,
            I => \N__24754\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__24775\,
            I => \N__24754\
        );

    \I__5705\ : Span4Mux_h
    port map (
            O => \N__24770\,
            I => \N__24751\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__24767\,
            I => \N__24748\
        );

    \I__5703\ : Odrv4
    port map (
            O => \N__24762\,
            I => \tok.n60\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__24759\,
            I => \tok.n60\
        );

    \I__5701\ : Odrv4
    port map (
            O => \N__24754\,
            I => \tok.n60\
        );

    \I__5700\ : Odrv4
    port map (
            O => \N__24751\,
            I => \tok.n60\
        );

    \I__5699\ : Odrv12
    port map (
            O => \N__24748\,
            I => \tok.n60\
        );

    \I__5698\ : InMux
    port map (
            O => \N__24737\,
            I => \N__24730\
        );

    \I__5697\ : InMux
    port map (
            O => \N__24736\,
            I => \N__24730\
        );

    \I__5696\ : InMux
    port map (
            O => \N__24735\,
            I => \N__24721\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__24730\,
            I => \N__24718\
        );

    \I__5694\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24713\
        );

    \I__5693\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24713\
        );

    \I__5692\ : InMux
    port map (
            O => \N__24727\,
            I => \N__24709\
        );

    \I__5691\ : InMux
    port map (
            O => \N__24726\,
            I => \N__24706\
        );

    \I__5690\ : InMux
    port map (
            O => \N__24725\,
            I => \N__24698\
        );

    \I__5689\ : InMux
    port map (
            O => \N__24724\,
            I => \N__24698\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__24721\,
            I => \N__24695\
        );

    \I__5687\ : Span4Mux_v
    port map (
            O => \N__24718\,
            I => \N__24692\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__24713\,
            I => \N__24689\
        );

    \I__5685\ : InMux
    port map (
            O => \N__24712\,
            I => \N__24686\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__24709\,
            I => \N__24683\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__24706\,
            I => \N__24680\
        );

    \I__5682\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24677\
        );

    \I__5681\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24672\
        );

    \I__5680\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24672\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__24698\,
            I => \N__24667\
        );

    \I__5678\ : Span4Mux_s2_v
    port map (
            O => \N__24695\,
            I => \N__24667\
        );

    \I__5677\ : Span4Mux_h
    port map (
            O => \N__24692\,
            I => \N__24660\
        );

    \I__5676\ : Span4Mux_v
    port map (
            O => \N__24689\,
            I => \N__24660\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__24686\,
            I => \N__24660\
        );

    \I__5674\ : Span12Mux_s5_v
    port map (
            O => \N__24683\,
            I => \N__24652\
        );

    \I__5673\ : Span12Mux_s5_h
    port map (
            O => \N__24680\,
            I => \N__24652\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__24677\,
            I => \N__24652\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__24672\,
            I => \N__24645\
        );

    \I__5670\ : Span4Mux_h
    port map (
            O => \N__24667\,
            I => \N__24645\
        );

    \I__5669\ : Span4Mux_h
    port map (
            O => \N__24660\,
            I => \N__24645\
        );

    \I__5668\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24642\
        );

    \I__5667\ : Odrv12
    port map (
            O => \N__24652\,
            I => \tok.n83\
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__24645\,
            I => \tok.n83\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__24642\,
            I => \tok.n83\
        );

    \I__5664\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24632\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__24632\,
            I => \N__24629\
        );

    \I__5662\ : Span4Mux_s3_v
    port map (
            O => \N__24629\,
            I => \N__24626\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__24626\,
            I => \tok.n3\
        );

    \I__5660\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24618\
        );

    \I__5659\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24615\
        );

    \I__5658\ : CascadeMux
    port map (
            O => \N__24621\,
            I => \N__24612\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__24618\,
            I => \N__24609\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__24615\,
            I => \N__24606\
        );

    \I__5655\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24603\
        );

    \I__5654\ : Span12Mux_s5_v
    port map (
            O => \N__24609\,
            I => \N__24600\
        );

    \I__5653\ : Span4Mux_v
    port map (
            O => \N__24606\,
            I => \N__24595\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__24603\,
            I => \N__24595\
        );

    \I__5651\ : Odrv12
    port map (
            O => \N__24600\,
            I => \tok.n4478\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__24595\,
            I => \tok.n4478\
        );

    \I__5649\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24586\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__24589\,
            I => \N__24580\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__24586\,
            I => \N__24577\
        );

    \I__5646\ : InMux
    port map (
            O => \N__24585\,
            I => \N__24574\
        );

    \I__5645\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24567\
        );

    \I__5644\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24567\
        );

    \I__5643\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24567\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__24577\,
            I => \tok.c_stk_r_5\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__24574\,
            I => \tok.c_stk_r_5\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__24567\,
            I => \tok.c_stk_r_5\
        );

    \I__5639\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__24557\,
            I => \N__24554\
        );

    \I__5637\ : Span4Mux_h
    port map (
            O => \N__24554\,
            I => \N__24550\
        );

    \I__5636\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24547\
        );

    \I__5635\ : Odrv4
    port map (
            O => \N__24550\,
            I => \tok.C_stk.tail_5\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__24547\,
            I => \tok.C_stk.tail_5\
        );

    \I__5633\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24536\
        );

    \I__5632\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24536\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__24536\,
            I => \tok.tail_13\
        );

    \I__5630\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24527\
        );

    \I__5629\ : InMux
    port map (
            O => \N__24532\,
            I => \N__24527\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__24527\,
            I => \tok.C_stk.tail_21\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__24524\,
            I => \N__24521\
        );

    \I__5626\ : InMux
    port map (
            O => \N__24521\,
            I => \N__24515\
        );

    \I__5625\ : InMux
    port map (
            O => \N__24520\,
            I => \N__24515\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__24515\,
            I => \N__24512\
        );

    \I__5623\ : Odrv4
    port map (
            O => \N__24512\,
            I => \tok.tail_29\
        );

    \I__5622\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24503\
        );

    \I__5621\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24503\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__24503\,
            I => \tok.C_stk.tail_37\
        );

    \I__5619\ : CascadeMux
    port map (
            O => \N__24500\,
            I => \tok.n4460_cascade_\
        );

    \I__5618\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24486\
        );

    \I__5617\ : InMux
    port map (
            O => \N__24496\,
            I => \N__24486\
        );

    \I__5616\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24482\
        );

    \I__5615\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24479\
        );

    \I__5614\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24474\
        );

    \I__5613\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24474\
        );

    \I__5612\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24466\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__24486\,
            I => \N__24463\
        );

    \I__5610\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24460\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__24482\,
            I => \N__24457\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__24479\,
            I => \N__24451\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__24474\,
            I => \N__24451\
        );

    \I__5606\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24448\
        );

    \I__5605\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24443\
        );

    \I__5604\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24443\
        );

    \I__5603\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24438\
        );

    \I__5602\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24438\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__24466\,
            I => \N__24435\
        );

    \I__5600\ : Span4Mux_s3_v
    port map (
            O => \N__24463\,
            I => \N__24428\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__24460\,
            I => \N__24428\
        );

    \I__5598\ : Span4Mux_v
    port map (
            O => \N__24457\,
            I => \N__24428\
        );

    \I__5597\ : InMux
    port map (
            O => \N__24456\,
            I => \N__24425\
        );

    \I__5596\ : Span4Mux_v
    port map (
            O => \N__24451\,
            I => \N__24420\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__24448\,
            I => \N__24420\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__24443\,
            I => \N__24415\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__24438\,
            I => \N__24415\
        );

    \I__5592\ : Span4Mux_s3_v
    port map (
            O => \N__24435\,
            I => \N__24408\
        );

    \I__5591\ : Span4Mux_h
    port map (
            O => \N__24428\,
            I => \N__24408\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__24425\,
            I => \N__24408\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__24420\,
            I => \N__24403\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__24415\,
            I => \N__24403\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__24408\,
            I => \N__24400\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__24403\,
            I => \tok.n2726\
        );

    \I__5585\ : Odrv4
    port map (
            O => \N__24400\,
            I => \tok.n2726\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__24395\,
            I => \N__24390\
        );

    \I__5583\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24386\
        );

    \I__5582\ : CascadeMux
    port map (
            O => \N__24393\,
            I => \N__24383\
        );

    \I__5581\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24380\
        );

    \I__5580\ : CascadeMux
    port map (
            O => \N__24389\,
            I => \N__24377\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__24386\,
            I => \N__24372\
        );

    \I__5578\ : InMux
    port map (
            O => \N__24383\,
            I => \N__24369\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__24380\,
            I => \N__24363\
        );

    \I__5576\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24360\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__24376\,
            I => \N__24357\
        );

    \I__5574\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24354\
        );

    \I__5573\ : Span4Mux_h
    port map (
            O => \N__24372\,
            I => \N__24349\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__24369\,
            I => \N__24349\
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__24368\,
            I => \N__24346\
        );

    \I__5570\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24343\
        );

    \I__5569\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24340\
        );

    \I__5568\ : Span4Mux_s3_h
    port map (
            O => \N__24363\,
            I => \N__24335\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__24360\,
            I => \N__24335\
        );

    \I__5566\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24332\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__24354\,
            I => \N__24329\
        );

    \I__5564\ : Span4Mux_v
    port map (
            O => \N__24349\,
            I => \N__24326\
        );

    \I__5563\ : InMux
    port map (
            O => \N__24346\,
            I => \N__24323\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__24343\,
            I => \N__24320\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__24340\,
            I => \N__24315\
        );

    \I__5560\ : Span4Mux_h
    port map (
            O => \N__24335\,
            I => \N__24315\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__24332\,
            I => \N__24306\
        );

    \I__5558\ : Span4Mux_v
    port map (
            O => \N__24329\,
            I => \N__24306\
        );

    \I__5557\ : Span4Mux_h
    port map (
            O => \N__24326\,
            I => \N__24306\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__24323\,
            I => \N__24306\
        );

    \I__5555\ : Span4Mux_v
    port map (
            O => \N__24320\,
            I => \N__24303\
        );

    \I__5554\ : Span4Mux_h
    port map (
            O => \N__24315\,
            I => \N__24300\
        );

    \I__5553\ : Odrv4
    port map (
            O => \N__24306\,
            I => \tok.S_4\
        );

    \I__5552\ : Odrv4
    port map (
            O => \N__24303\,
            I => \tok.S_4\
        );

    \I__5551\ : Odrv4
    port map (
            O => \N__24300\,
            I => \tok.S_4\
        );

    \I__5550\ : InMux
    port map (
            O => \N__24293\,
            I => \N__24290\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__5548\ : Span4Mux_s3_h
    port map (
            O => \N__24287\,
            I => \N__24284\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__24284\,
            I => \tok.n13_adj_787\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__24281\,
            I => \tok.n10_adj_829_cascade_\
        );

    \I__5545\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24275\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__24275\,
            I => \N__24272\
        );

    \I__5543\ : Odrv12
    port map (
            O => \N__24272\,
            I => \tok.n13_adj_833\
        );

    \I__5542\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24265\
        );

    \I__5541\ : InMux
    port map (
            O => \N__24268\,
            I => \N__24262\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__24265\,
            I => \N__24258\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__24262\,
            I => \N__24255\
        );

    \I__5538\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24252\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__24258\,
            I => \N__24247\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__24255\,
            I => \N__24247\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__24252\,
            I => \tok.n2746\
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__24247\,
            I => \tok.n2746\
        );

    \I__5533\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24239\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__24239\,
            I => \N__24236\
        );

    \I__5531\ : Odrv12
    port map (
            O => \N__24236\,
            I => \tok.n8_adj_839\
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__24233\,
            I => \N__24230\
        );

    \I__5529\ : InMux
    port map (
            O => \N__24230\,
            I => \N__24227\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__24227\,
            I => \N__24223\
        );

    \I__5527\ : CascadeMux
    port map (
            O => \N__24226\,
            I => \N__24220\
        );

    \I__5526\ : Span4Mux_s3_v
    port map (
            O => \N__24223\,
            I => \N__24217\
        );

    \I__5525\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24214\
        );

    \I__5524\ : Span4Mux_h
    port map (
            O => \N__24217\,
            I => \N__24211\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24208\
        );

    \I__5522\ : Span4Mux_v
    port map (
            O => \N__24211\,
            I => \N__24205\
        );

    \I__5521\ : Odrv12
    port map (
            O => \N__24208\,
            I => \tok.table_rd_0\
        );

    \I__5520\ : Odrv4
    port map (
            O => \N__24205\,
            I => \tok.table_rd_0\
        );

    \I__5519\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24197\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__5517\ : Span4Mux_v
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__5516\ : Odrv4
    port map (
            O => \N__24191\,
            I => \tok.n18_adj_681\
        );

    \I__5515\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24182\
        );

    \I__5514\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24177\
        );

    \I__5513\ : InMux
    port map (
            O => \N__24186\,
            I => \N__24174\
        );

    \I__5512\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24170\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__24182\,
            I => \N__24165\
        );

    \I__5510\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24162\
        );

    \I__5509\ : InMux
    port map (
            O => \N__24180\,
            I => \N__24159\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__24177\,
            I => \N__24156\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__24174\,
            I => \N__24153\
        );

    \I__5506\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24150\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__24170\,
            I => \N__24146\
        );

    \I__5504\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24141\
        );

    \I__5503\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24141\
        );

    \I__5502\ : Span4Mux_s2_v
    port map (
            O => \N__24165\,
            I => \N__24137\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__24162\,
            I => \N__24132\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__24159\,
            I => \N__24132\
        );

    \I__5499\ : Span4Mux_h
    port map (
            O => \N__24156\,
            I => \N__24122\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__24153\,
            I => \N__24122\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__24150\,
            I => \N__24122\
        );

    \I__5496\ : CascadeMux
    port map (
            O => \N__24149\,
            I => \N__24119\
        );

    \I__5495\ : Span4Mux_v
    port map (
            O => \N__24146\,
            I => \N__24113\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__24141\,
            I => \N__24113\
        );

    \I__5493\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24110\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__24137\,
            I => \N__24105\
        );

    \I__5491\ : Span4Mux_v
    port map (
            O => \N__24132\,
            I => \N__24105\
        );

    \I__5490\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24102\
        );

    \I__5489\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24097\
        );

    \I__5488\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24097\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__24122\,
            I => \N__24094\
        );

    \I__5486\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24089\
        );

    \I__5485\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24089\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__24113\,
            I => \tok.A_low_1\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__24110\,
            I => \tok.A_low_1\
        );

    \I__5482\ : Odrv4
    port map (
            O => \N__24105\,
            I => \tok.A_low_1\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__24102\,
            I => \tok.A_low_1\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__24097\,
            I => \tok.A_low_1\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__24094\,
            I => \tok.A_low_1\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__24089\,
            I => \tok.A_low_1\
        );

    \I__5477\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24070\
        );

    \I__5476\ : InMux
    port map (
            O => \N__24073\,
            I => \N__24063\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__24070\,
            I => \N__24060\
        );

    \I__5474\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24057\
        );

    \I__5473\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24054\
        );

    \I__5472\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24051\
        );

    \I__5471\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24048\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__24063\,
            I => \N__24045\
        );

    \I__5469\ : Span4Mux_v
    port map (
            O => \N__24060\,
            I => \N__24042\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__24057\,
            I => \N__24039\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__24054\,
            I => \N__24036\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__24051\,
            I => \N__24031\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24031\
        );

    \I__5464\ : Span4Mux_v
    port map (
            O => \N__24045\,
            I => \N__24022\
        );

    \I__5463\ : Span4Mux_h
    port map (
            O => \N__24042\,
            I => \N__24022\
        );

    \I__5462\ : Span4Mux_v
    port map (
            O => \N__24039\,
            I => \N__24022\
        );

    \I__5461\ : Span4Mux_s2_h
    port map (
            O => \N__24036\,
            I => \N__24022\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__24031\,
            I => \N__24019\
        );

    \I__5459\ : Odrv4
    port map (
            O => \N__24022\,
            I => \tok.n101\
        );

    \I__5458\ : Odrv4
    port map (
            O => \N__24019\,
            I => \tok.n101\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__24014\,
            I => \N__24010\
        );

    \I__5456\ : InMux
    port map (
            O => \N__24013\,
            I => \N__24005\
        );

    \I__5455\ : InMux
    port map (
            O => \N__24010\,
            I => \N__24000\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__24009\,
            I => \N__23997\
        );

    \I__5453\ : InMux
    port map (
            O => \N__24008\,
            I => \N__23994\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__24005\,
            I => \N__23991\
        );

    \I__5451\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23988\
        );

    \I__5450\ : InMux
    port map (
            O => \N__24003\,
            I => \N__23985\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__24000\,
            I => \N__23979\
        );

    \I__5448\ : InMux
    port map (
            O => \N__23997\,
            I => \N__23976\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__23994\,
            I => \N__23971\
        );

    \I__5446\ : Span4Mux_v
    port map (
            O => \N__23991\,
            I => \N__23971\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__23988\,
            I => \N__23968\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__23985\,
            I => \N__23965\
        );

    \I__5443\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23962\
        );

    \I__5442\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23959\
        );

    \I__5441\ : CascadeMux
    port map (
            O => \N__23982\,
            I => \N__23956\
        );

    \I__5440\ : Span4Mux_h
    port map (
            O => \N__23979\,
            I => \N__23953\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__23976\,
            I => \N__23947\
        );

    \I__5438\ : Span4Mux_h
    port map (
            O => \N__23971\,
            I => \N__23947\
        );

    \I__5437\ : Span4Mux_h
    port map (
            O => \N__23968\,
            I => \N__23942\
        );

    \I__5436\ : Span4Mux_v
    port map (
            O => \N__23965\,
            I => \N__23942\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__23962\,
            I => \N__23937\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__23959\,
            I => \N__23937\
        );

    \I__5433\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23934\
        );

    \I__5432\ : Span4Mux_h
    port map (
            O => \N__23953\,
            I => \N__23931\
        );

    \I__5431\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23928\
        );

    \I__5430\ : Span4Mux_v
    port map (
            O => \N__23947\,
            I => \N__23925\
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__23942\,
            I => \tok.n54\
        );

    \I__5428\ : Odrv12
    port map (
            O => \N__23937\,
            I => \tok.n54\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__23934\,
            I => \tok.n54\
        );

    \I__5426\ : Odrv4
    port map (
            O => \N__23931\,
            I => \tok.n54\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__23928\,
            I => \tok.n54\
        );

    \I__5424\ : Odrv4
    port map (
            O => \N__23925\,
            I => \tok.n54\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__23912\,
            I => \tok.n244_cascade_\
        );

    \I__5422\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23906\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__23906\,
            I => \N__23903\
        );

    \I__5420\ : Odrv12
    port map (
            O => \N__23903\,
            I => \tok.n17_adj_785\
        );

    \I__5419\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23890\
        );

    \I__5418\ : InMux
    port map (
            O => \N__23899\,
            I => \N__23879\
        );

    \I__5417\ : InMux
    port map (
            O => \N__23898\,
            I => \N__23879\
        );

    \I__5416\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23879\
        );

    \I__5415\ : InMux
    port map (
            O => \N__23896\,
            I => \N__23879\
        );

    \I__5414\ : InMux
    port map (
            O => \N__23895\,
            I => \N__23879\
        );

    \I__5413\ : CascadeMux
    port map (
            O => \N__23894\,
            I => \N__23872\
        );

    \I__5412\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23862\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__23890\,
            I => \N__23859\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23856\
        );

    \I__5409\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23847\
        );

    \I__5408\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23847\
        );

    \I__5407\ : InMux
    port map (
            O => \N__23876\,
            I => \N__23847\
        );

    \I__5406\ : InMux
    port map (
            O => \N__23875\,
            I => \N__23847\
        );

    \I__5405\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23838\
        );

    \I__5404\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23838\
        );

    \I__5403\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23838\
        );

    \I__5402\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23838\
        );

    \I__5401\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23833\
        );

    \I__5400\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23833\
        );

    \I__5399\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23828\
        );

    \I__5398\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23828\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__23862\,
            I => \N__23825\
        );

    \I__5396\ : Span4Mux_v
    port map (
            O => \N__23859\,
            I => \N__23818\
        );

    \I__5395\ : Span4Mux_v
    port map (
            O => \N__23856\,
            I => \N__23818\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__23847\,
            I => \N__23818\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__23838\,
            I => \N__23815\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__23833\,
            I => \N__23812\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__23828\,
            I => \N__23809\
        );

    \I__5390\ : Span4Mux_v
    port map (
            O => \N__23825\,
            I => \N__23802\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__23818\,
            I => \N__23802\
        );

    \I__5388\ : Span4Mux_v
    port map (
            O => \N__23815\,
            I => \N__23802\
        );

    \I__5387\ : Span4Mux_v
    port map (
            O => \N__23812\,
            I => \N__23798\
        );

    \I__5386\ : Span4Mux_h
    port map (
            O => \N__23809\,
            I => \N__23795\
        );

    \I__5385\ : Span4Mux_h
    port map (
            O => \N__23802\,
            I => \N__23792\
        );

    \I__5384\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23789\
        );

    \I__5383\ : Odrv4
    port map (
            O => \N__23798\,
            I => \tok.n11_adj_647\
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__23795\,
            I => \tok.n11_adj_647\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__23792\,
            I => \tok.n11_adj_647\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__23789\,
            I => \tok.n11_adj_647\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__23780\,
            I => \tok.n4575_cascade_\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__23777\,
            I => \tok.n83_cascade_\
        );

    \I__5377\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23768\
        );

    \I__5376\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23768\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__23768\,
            I => \N__23765\
        );

    \I__5374\ : Span4Mux_s3_h
    port map (
            O => \N__23765\,
            I => \N__23762\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__23762\,
            I => \tok.n40\
        );

    \I__5372\ : CascadeMux
    port map (
            O => \N__23759\,
            I => \tok.n4571_cascade_\
        );

    \I__5371\ : InMux
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__23753\,
            I => \tok.n4393\
        );

    \I__5369\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23747\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__23747\,
            I => \N__23741\
        );

    \I__5367\ : InMux
    port map (
            O => \N__23746\,
            I => \N__23736\
        );

    \I__5366\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23736\
        );

    \I__5365\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23733\
        );

    \I__5364\ : Span4Mux_v
    port map (
            O => \N__23741\,
            I => \N__23728\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23728\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__23733\,
            I => \N__23725\
        );

    \I__5361\ : Span4Mux_h
    port map (
            O => \N__23728\,
            I => \N__23720\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__23725\,
            I => \N__23720\
        );

    \I__5359\ : Odrv4
    port map (
            O => \N__23720\,
            I => \tok.n9_adj_797\
        );

    \I__5358\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__23714\,
            I => \tok.n13_adj_758\
        );

    \I__5356\ : InMux
    port map (
            O => \N__23711\,
            I => \N__23708\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__23708\,
            I => \N__23705\
        );

    \I__5354\ : Odrv12
    port map (
            O => \N__23705\,
            I => n10_adj_873
        );

    \I__5353\ : CascadeMux
    port map (
            O => \N__23702\,
            I => \n10_adj_873_cascade_\
        );

    \I__5352\ : CascadeMux
    port map (
            O => \N__23699\,
            I => \N__23696\
        );

    \I__5351\ : InMux
    port map (
            O => \N__23696\,
            I => \N__23693\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__23693\,
            I => \N__23688\
        );

    \I__5349\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23685\
        );

    \I__5348\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23681\
        );

    \I__5347\ : Span4Mux_s3_h
    port map (
            O => \N__23688\,
            I => \N__23678\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__23685\,
            I => \N__23675\
        );

    \I__5345\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23672\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__23681\,
            I => \c_stk_w_7_N_18_5\
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__23678\,
            I => \c_stk_w_7_N_18_5\
        );

    \I__5342\ : Odrv12
    port map (
            O => \N__23675\,
            I => \c_stk_w_7_N_18_5\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__23672\,
            I => \c_stk_w_7_N_18_5\
        );

    \I__5340\ : CascadeMux
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__5339\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23657\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__23657\,
            I => \tok.tc_5\
        );

    \I__5337\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__23651\,
            I => \N__23648\
        );

    \I__5335\ : Span4Mux_h
    port map (
            O => \N__23648\,
            I => \N__23645\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__23645\,
            I => n10_adj_874
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__23642\,
            I => \n10_adj_874_cascade_\
        );

    \I__5332\ : CascadeMux
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__5331\ : InMux
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__5329\ : Odrv4
    port map (
            O => \N__23630\,
            I => \tok.tc_2\
        );

    \I__5328\ : CascadeMux
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__5327\ : InMux
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__23621\,
            I => \N__23616\
        );

    \I__5325\ : InMux
    port map (
            O => \N__23620\,
            I => \N__23610\
        );

    \I__5324\ : InMux
    port map (
            O => \N__23619\,
            I => \N__23610\
        );

    \I__5323\ : Span4Mux_v
    port map (
            O => \N__23616\,
            I => \N__23607\
        );

    \I__5322\ : InMux
    port map (
            O => \N__23615\,
            I => \N__23604\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__23610\,
            I => \N__23601\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__23607\,
            I => \N__23598\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__23604\,
            I => \N__23595\
        );

    \I__5318\ : Span4Mux_s3_h
    port map (
            O => \N__23601\,
            I => \N__23592\
        );

    \I__5317\ : Odrv4
    port map (
            O => \N__23598\,
            I => \tok.tc_plus_1_3\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__23595\,
            I => \tok.tc_plus_1_3\
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__23592\,
            I => \tok.tc_plus_1_3\
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__5313\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23579\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__5311\ : Odrv4
    port map (
            O => \N__23576\,
            I => n92_adj_870
        );

    \I__5310\ : CascadeMux
    port map (
            O => \N__23573\,
            I => \n92_adj_870_cascade_\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__5308\ : InMux
    port map (
            O => \N__23567\,
            I => \N__23564\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__23564\,
            I => \N__23559\
        );

    \I__5306\ : InMux
    port map (
            O => \N__23563\,
            I => \N__23556\
        );

    \I__5305\ : InMux
    port map (
            O => \N__23562\,
            I => \N__23552\
        );

    \I__5304\ : Span4Mux_v
    port map (
            O => \N__23559\,
            I => \N__23549\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__23556\,
            I => \N__23546\
        );

    \I__5302\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23543\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__23552\,
            I => \c_stk_w_7_N_18_3\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__23549\,
            I => \c_stk_w_7_N_18_3\
        );

    \I__5299\ : Odrv12
    port map (
            O => \N__23546\,
            I => \c_stk_w_7_N_18_3\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__23543\,
            I => \c_stk_w_7_N_18_3\
        );

    \I__5297\ : CascadeMux
    port map (
            O => \N__23534\,
            I => \N__23531\
        );

    \I__5296\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23528\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__23528\,
            I => \N__23525\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__23525\,
            I => \tok.tc_3\
        );

    \I__5293\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23507\
        );

    \I__5292\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23507\
        );

    \I__5291\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23507\
        );

    \I__5290\ : InMux
    port map (
            O => \N__23519\,
            I => \N__23507\
        );

    \I__5289\ : InMux
    port map (
            O => \N__23518\,
            I => \N__23493\
        );

    \I__5288\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23493\
        );

    \I__5287\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23490\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__23507\,
            I => \N__23487\
        );

    \I__5285\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23470\
        );

    \I__5284\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23470\
        );

    \I__5283\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23470\
        );

    \I__5282\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23470\
        );

    \I__5281\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23470\
        );

    \I__5280\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23470\
        );

    \I__5279\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23470\
        );

    \I__5278\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23470\
        );

    \I__5277\ : InMux
    port map (
            O => \N__23498\,
            I => \N__23467\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__23493\,
            I => \N__23464\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__23490\,
            I => \N__23461\
        );

    \I__5274\ : Span4Mux_v
    port map (
            O => \N__23487\,
            I => \N__23458\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__23470\,
            I => \stall_\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__23467\,
            I => \stall_\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__23464\,
            I => \stall_\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__23461\,
            I => \stall_\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__23458\,
            I => \stall_\
        );

    \I__5268\ : CascadeMux
    port map (
            O => \N__23447\,
            I => \N__23444\
        );

    \I__5267\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23441\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__23441\,
            I => \tok.tc_4\
        );

    \I__5265\ : CascadeMux
    port map (
            O => \N__23438\,
            I => \tok.C_stk.n4900_cascade_\
        );

    \I__5264\ : CascadeMux
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__5263\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23429\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__23429\,
            I => \N__23425\
        );

    \I__5261\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23422\
        );

    \I__5260\ : Span4Mux_v
    port map (
            O => \N__23425\,
            I => \N__23419\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__23422\,
            I => \N__23416\
        );

    \I__5258\ : Span4Mux_h
    port map (
            O => \N__23419\,
            I => \N__23413\
        );

    \I__5257\ : Span4Mux_v
    port map (
            O => \N__23416\,
            I => \N__23410\
        );

    \I__5256\ : Span4Mux_h
    port map (
            O => \N__23413\,
            I => \N__23407\
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__23410\,
            I => \tok.table_rd_5\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__23407\,
            I => \tok.table_rd_5\
        );

    \I__5253\ : CascadeMux
    port map (
            O => \N__23402\,
            I => \tok.n83_adj_742_cascade_\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__23399\,
            I => \tok.n4651_cascade_\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__23396\,
            I => \tok.ram.n4702_cascade_\
        );

    \I__5250\ : InMux
    port map (
            O => \N__23393\,
            I => \N__23390\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__23390\,
            I => \tok.n1_adj_757\
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__23387\,
            I => \N__23384\
        );

    \I__5247\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23380\
        );

    \I__5246\ : InMux
    port map (
            O => \N__23383\,
            I => \N__23377\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__23380\,
            I => \N__23374\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__23377\,
            I => \N__23369\
        );

    \I__5243\ : Span4Mux_v
    port map (
            O => \N__23374\,
            I => \N__23366\
        );

    \I__5242\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23361\
        );

    \I__5241\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23361\
        );

    \I__5240\ : Span4Mux_v
    port map (
            O => \N__23369\,
            I => \N__23356\
        );

    \I__5239\ : Span4Mux_s2_h
    port map (
            O => \N__23366\,
            I => \N__23356\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__23361\,
            I => \N__23353\
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__23356\,
            I => \tok.tc_plus_1_5\
        );

    \I__5236\ : Odrv4
    port map (
            O => \N__23353\,
            I => \tok.tc_plus_1_5\
        );

    \I__5235\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__23345\,
            I => \N__23341\
        );

    \I__5233\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23338\
        );

    \I__5232\ : Span4Mux_v
    port map (
            O => \N__23341\,
            I => \N__23335\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__23338\,
            I => \tok.tail_44\
        );

    \I__5230\ : Odrv4
    port map (
            O => \N__23335\,
            I => \tok.tail_44\
        );

    \I__5229\ : InMux
    port map (
            O => \N__23330\,
            I => \N__23327\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__5227\ : Span4Mux_s3_h
    port map (
            O => \N__23324\,
            I => \N__23320\
        );

    \I__5226\ : InMux
    port map (
            O => \N__23323\,
            I => \N__23317\
        );

    \I__5225\ : Odrv4
    port map (
            O => \N__23320\,
            I => \tok.C_stk.tail_18\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__23317\,
            I => \tok.C_stk.tail_18\
        );

    \I__5223\ : CascadeMux
    port map (
            O => \N__23312\,
            I => \N__23308\
        );

    \I__5222\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23303\
        );

    \I__5221\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23303\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__5219\ : Span4Mux_s2_h
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__23297\,
            I => \N__23294\
        );

    \I__5217\ : Odrv4
    port map (
            O => \N__23294\,
            I => \tok.n240\
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__23291\,
            I => \N__23287\
        );

    \I__5215\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23284\
        );

    \I__5214\ : InMux
    port map (
            O => \N__23287\,
            I => \N__23281\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__23284\,
            I => \N__23278\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__23281\,
            I => \N__23275\
        );

    \I__5211\ : Odrv4
    port map (
            O => \N__23278\,
            I => \tok.tail_55\
        );

    \I__5210\ : Odrv12
    port map (
            O => \N__23275\,
            I => \tok.tail_55\
        );

    \I__5209\ : InMux
    port map (
            O => \N__23270\,
            I => \N__23267\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__23267\,
            I => \N__23263\
        );

    \I__5207\ : InMux
    port map (
            O => \N__23266\,
            I => \N__23260\
        );

    \I__5206\ : Odrv4
    port map (
            O => \N__23263\,
            I => \tok.tail_63\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__23260\,
            I => \tok.tail_63\
        );

    \I__5204\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23251\
        );

    \I__5203\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23248\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__23251\,
            I => \tok.tail_54\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__23248\,
            I => \tok.tail_54\
        );

    \I__5200\ : InMux
    port map (
            O => \N__23243\,
            I => \N__23239\
        );

    \I__5199\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23236\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__23239\,
            I => \tok.tail_62\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__23236\,
            I => \tok.tail_62\
        );

    \I__5196\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23227\
        );

    \I__5195\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23224\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__23227\,
            I => \N__23221\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__23224\,
            I => \N__23218\
        );

    \I__5192\ : Span4Mux_h
    port map (
            O => \N__23221\,
            I => \N__23215\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__23218\,
            I => \tok.tail_52\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__23215\,
            I => \tok.tail_52\
        );

    \I__5189\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23206\
        );

    \I__5188\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23203\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__23206\,
            I => \tok.tail_60\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__23203\,
            I => \tok.tail_60\
        );

    \I__5185\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23192\
        );

    \I__5184\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23192\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__23192\,
            I => \tok.C_stk.tail_39\
        );

    \I__5182\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23183\
        );

    \I__5181\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23183\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__23183\,
            I => \tok.tail_47\
        );

    \I__5179\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23174\
        );

    \I__5178\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23174\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__23174\,
            I => \tok.C_stk.tail_16\
        );

    \I__5176\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23168\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23164\
        );

    \I__5174\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23161\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__23164\,
            I => \tok.C_stk.tail_32\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__23161\,
            I => \tok.C_stk.tail_32\
        );

    \I__5171\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23152\
        );

    \I__5170\ : InMux
    port map (
            O => \N__23155\,
            I => \N__23149\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__23152\,
            I => \N__23146\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__23149\,
            I => \tok.tail_24\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__23146\,
            I => \tok.tail_24\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__23141\,
            I => \N__23138\
        );

    \I__5165\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23132\
        );

    \I__5164\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23132\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__23132\,
            I => \tok.tail_30\
        );

    \I__5162\ : InMux
    port map (
            O => \N__23129\,
            I => \N__23123\
        );

    \I__5161\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23123\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__23123\,
            I => \tok.C_stk.tail_38\
        );

    \I__5159\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23114\
        );

    \I__5158\ : InMux
    port map (
            O => \N__23119\,
            I => \N__23114\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__23114\,
            I => \tok.tail_46\
        );

    \I__5156\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23107\
        );

    \I__5155\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23103\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__23107\,
            I => \N__23100\
        );

    \I__5153\ : CascadeMux
    port map (
            O => \N__23106\,
            I => \N__23095\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__23103\,
            I => \N__23092\
        );

    \I__5151\ : Span4Mux_h
    port map (
            O => \N__23100\,
            I => \N__23089\
        );

    \I__5150\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23086\
        );

    \I__5149\ : InMux
    port map (
            O => \N__23098\,
            I => \N__23081\
        );

    \I__5148\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23081\
        );

    \I__5147\ : Span4Mux_v
    port map (
            O => \N__23092\,
            I => \N__23078\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__23089\,
            I => \tok.c_stk_r_6\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__23086\,
            I => \tok.c_stk_r_6\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__23081\,
            I => \tok.c_stk_r_6\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__23078\,
            I => \tok.c_stk_r_6\
        );

    \I__5142\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__23066\,
            I => \N__23063\
        );

    \I__5140\ : Span12Mux_s6_v
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__5139\ : Odrv12
    port map (
            O => \N__23060\,
            I => \tok.n9_adj_807\
        );

    \I__5138\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23051\
        );

    \I__5137\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23051\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__23051\,
            I => uart_rx_data_4
        );

    \I__5135\ : InMux
    port map (
            O => \N__23048\,
            I => \N__23045\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__23045\,
            I => \N__23042\
        );

    \I__5133\ : Span4Mux_h
    port map (
            O => \N__23042\,
            I => \N__23039\
        );

    \I__5132\ : Span4Mux_h
    port map (
            O => \N__23039\,
            I => \N__23036\
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__23036\,
            I => \tok.n3_adj_826\
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__23033\,
            I => \tok.n6_adj_827_cascade_\
        );

    \I__5129\ : InMux
    port map (
            O => \N__23030\,
            I => \N__23027\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__23027\,
            I => \N__23024\
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__23024\,
            I => \tok.n36\
        );

    \I__5126\ : CascadeMux
    port map (
            O => \N__23021\,
            I => \tok.n33_adj_828_cascade_\
        );

    \I__5125\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23015\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__23015\,
            I => \N__23012\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__23012\,
            I => \N__23009\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__23009\,
            I => \tok.n11_adj_831\
        );

    \I__5121\ : InMux
    port map (
            O => \N__23006\,
            I => \N__23000\
        );

    \I__5120\ : InMux
    port map (
            O => \N__23005\,
            I => \N__22997\
        );

    \I__5119\ : InMux
    port map (
            O => \N__23004\,
            I => \N__22989\
        );

    \I__5118\ : InMux
    port map (
            O => \N__23003\,
            I => \N__22989\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22986\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__22997\,
            I => \N__22983\
        );

    \I__5115\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22980\
        );

    \I__5114\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22976\
        );

    \I__5113\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22973\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__22989\,
            I => \N__22970\
        );

    \I__5111\ : Span4Mux_s1_v
    port map (
            O => \N__22986\,
            I => \N__22966\
        );

    \I__5110\ : Span4Mux_v
    port map (
            O => \N__22983\,
            I => \N__22961\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__22980\,
            I => \N__22961\
        );

    \I__5108\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22958\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__22976\,
            I => \N__22955\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__22973\,
            I => \N__22952\
        );

    \I__5105\ : Span4Mux_v
    port map (
            O => \N__22970\,
            I => \N__22949\
        );

    \I__5104\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22946\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__22966\,
            I => \N__22939\
        );

    \I__5102\ : Span4Mux_h
    port map (
            O => \N__22961\,
            I => \N__22939\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__22958\,
            I => \N__22939\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__22955\,
            I => \N__22936\
        );

    \I__5099\ : Span4Mux_s3_v
    port map (
            O => \N__22952\,
            I => \N__22933\
        );

    \I__5098\ : Span4Mux_h
    port map (
            O => \N__22949\,
            I => \N__22925\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__22946\,
            I => \N__22925\
        );

    \I__5096\ : Span4Mux_v
    port map (
            O => \N__22939\,
            I => \N__22925\
        );

    \I__5095\ : Span4Mux_v
    port map (
            O => \N__22936\,
            I => \N__22920\
        );

    \I__5094\ : Span4Mux_h
    port map (
            O => \N__22933\,
            I => \N__22920\
        );

    \I__5093\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22917\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__22925\,
            I => \N__22914\
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__22920\,
            I => \tok.n56\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__22917\,
            I => \tok.n56\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__22914\,
            I => \tok.n56\
        );

    \I__5088\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22904\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__22904\,
            I => \N__22901\
        );

    \I__5086\ : Span4Mux_h
    port map (
            O => \N__22901\,
            I => \N__22898\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__22898\,
            I => \N__22895\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__22895\,
            I => \tok.n2514\
        );

    \I__5083\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22889\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__22889\,
            I => \N__22885\
        );

    \I__5081\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22882\
        );

    \I__5080\ : Span4Mux_s3_h
    port map (
            O => \N__22885\,
            I => \N__22879\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__22882\,
            I => \tok.C_stk.tail_0\
        );

    \I__5078\ : Odrv4
    port map (
            O => \N__22879\,
            I => \tok.C_stk.tail_0\
        );

    \I__5077\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22871\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__5075\ : Span4Mux_s1_v
    port map (
            O => \N__22868\,
            I => \N__22864\
        );

    \I__5074\ : InMux
    port map (
            O => \N__22867\,
            I => \N__22861\
        );

    \I__5073\ : Odrv4
    port map (
            O => \N__22864\,
            I => \tok.tail_8\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__22861\,
            I => \tok.tail_8\
        );

    \I__5071\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22852\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__22855\,
            I => \N__22849\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__22852\,
            I => \N__22846\
        );

    \I__5068\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22843\
        );

    \I__5067\ : Odrv4
    port map (
            O => \N__22846\,
            I => \tok.tail_15\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__22843\,
            I => \tok.tail_15\
        );

    \I__5065\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22835\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__22835\,
            I => \N__22832\
        );

    \I__5063\ : Span4Mux_s1_v
    port map (
            O => \N__22832\,
            I => \N__22828\
        );

    \I__5062\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22825\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__22828\,
            I => \tok.C_stk.tail_23\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__22825\,
            I => \tok.C_stk.tail_23\
        );

    \I__5059\ : InMux
    port map (
            O => \N__22820\,
            I => \N__22814\
        );

    \I__5058\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22814\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__22814\,
            I => \tok.tail_31\
        );

    \I__5056\ : InMux
    port map (
            O => \N__22811\,
            I => \N__22808\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__22808\,
            I => \tok.n211\
        );

    \I__5054\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22799\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__22799\,
            I => \tok.n2_adj_810\
        );

    \I__5051\ : InMux
    port map (
            O => \N__22796\,
            I => \N__22793\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__22793\,
            I => \N__22790\
        );

    \I__5049\ : Odrv4
    port map (
            O => \N__22790\,
            I => \tok.n5_adj_710\
        );

    \I__5048\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22784\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__22784\,
            I => \N__22781\
        );

    \I__5046\ : Span4Mux_h
    port map (
            O => \N__22781\,
            I => \N__22778\
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__22778\,
            I => \tok.n6_adj_711\
        );

    \I__5044\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__5042\ : Span12Mux_s7_h
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__5041\ : Odrv12
    port map (
            O => \N__22766\,
            I => \tok.n4664\
        );

    \I__5040\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__5038\ : Odrv4
    port map (
            O => \N__22757\,
            I => \tok.n4663\
        );

    \I__5037\ : InMux
    port map (
            O => \N__22754\,
            I => \N__22751\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__22751\,
            I => \tok.n33\
        );

    \I__5035\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22745\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__22745\,
            I => \N__22742\
        );

    \I__5033\ : Odrv12
    port map (
            O => \N__22742\,
            I => \tok.n27\
        );

    \I__5032\ : CascadeMux
    port map (
            O => \N__22739\,
            I => \N__22736\
        );

    \I__5031\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__5029\ : Span4Mux_h
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__5028\ : Span4Mux_h
    port map (
            O => \N__22727\,
            I => \N__22724\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__22724\,
            I => \tok.n296\
        );

    \I__5026\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22713\
        );

    \I__5025\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22710\
        );

    \I__5024\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22705\
        );

    \I__5023\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22705\
        );

    \I__5022\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22702\
        );

    \I__5021\ : CascadeMux
    port map (
            O => \N__22716\,
            I => \N__22698\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__22713\,
            I => \N__22694\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__22710\,
            I => \N__22691\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__22705\,
            I => \N__22688\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__22702\,
            I => \N__22685\
        );

    \I__5016\ : InMux
    port map (
            O => \N__22701\,
            I => \N__22680\
        );

    \I__5015\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22680\
        );

    \I__5014\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22677\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__22694\,
            I => \N__22672\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__22691\,
            I => \N__22672\
        );

    \I__5011\ : Span12Mux_s5_h
    port map (
            O => \N__22688\,
            I => \N__22665\
        );

    \I__5010\ : Span12Mux_s11_v
    port map (
            O => \N__22685\,
            I => \N__22665\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__22680\,
            I => \N__22665\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__22677\,
            I => \tok.n191\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__22672\,
            I => \tok.n191\
        );

    \I__5006\ : Odrv12
    port map (
            O => \N__22665\,
            I => \tok.n191\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__22658\,
            I => \N__22652\
        );

    \I__5004\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22647\
        );

    \I__5003\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22644\
        );

    \I__5002\ : InMux
    port map (
            O => \N__22655\,
            I => \N__22641\
        );

    \I__5001\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22637\
        );

    \I__5000\ : InMux
    port map (
            O => \N__22651\,
            I => \N__22633\
        );

    \I__4999\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22628\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__22647\,
            I => \N__22625\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__22644\,
            I => \N__22622\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__22641\,
            I => \N__22619\
        );

    \I__4995\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22616\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__22637\,
            I => \N__22613\
        );

    \I__4993\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22610\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__22633\,
            I => \N__22607\
        );

    \I__4991\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22604\
        );

    \I__4990\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22601\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__22628\,
            I => \N__22598\
        );

    \I__4988\ : Span4Mux_v
    port map (
            O => \N__22625\,
            I => \N__22593\
        );

    \I__4987\ : Span4Mux_v
    port map (
            O => \N__22622\,
            I => \N__22593\
        );

    \I__4986\ : Span4Mux_h
    port map (
            O => \N__22619\,
            I => \N__22590\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__22616\,
            I => \N__22583\
        );

    \I__4984\ : Span4Mux_h
    port map (
            O => \N__22613\,
            I => \N__22583\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__22610\,
            I => \N__22580\
        );

    \I__4982\ : Span4Mux_s2_h
    port map (
            O => \N__22607\,
            I => \N__22577\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__22604\,
            I => \N__22566\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22566\
        );

    \I__4979\ : Span4Mux_v
    port map (
            O => \N__22598\,
            I => \N__22566\
        );

    \I__4978\ : Span4Mux_h
    port map (
            O => \N__22593\,
            I => \N__22566\
        );

    \I__4977\ : Span4Mux_v
    port map (
            O => \N__22590\,
            I => \N__22566\
        );

    \I__4976\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22561\
        );

    \I__4975\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22561\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__22583\,
            I => \N__22558\
        );

    \I__4973\ : Span4Mux_h
    port map (
            O => \N__22580\,
            I => \N__22555\
        );

    \I__4972\ : Span4Mux_v
    port map (
            O => \N__22577\,
            I => \N__22550\
        );

    \I__4971\ : Span4Mux_h
    port map (
            O => \N__22566\,
            I => \N__22550\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__22561\,
            I => \tok.n59\
        );

    \I__4969\ : Odrv4
    port map (
            O => \N__22558\,
            I => \tok.n59\
        );

    \I__4968\ : Odrv4
    port map (
            O => \N__22555\,
            I => \tok.n59\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__22550\,
            I => \tok.n59\
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__4965\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__22532\,
            I => \tok.n2_adj_703\
        );

    \I__4962\ : CascadeMux
    port map (
            O => \N__22529\,
            I => \N__22523\
        );

    \I__4961\ : InMux
    port map (
            O => \N__22528\,
            I => \N__22516\
        );

    \I__4960\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22513\
        );

    \I__4959\ : InMux
    port map (
            O => \N__22526\,
            I => \N__22508\
        );

    \I__4958\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22508\
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__22522\,
            I => \N__22504\
        );

    \I__4956\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22500\
        );

    \I__4955\ : InMux
    port map (
            O => \N__22520\,
            I => \N__22497\
        );

    \I__4954\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22494\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__22516\,
            I => \N__22486\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__22513\,
            I => \N__22481\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__22508\,
            I => \N__22481\
        );

    \I__4950\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22474\
        );

    \I__4949\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22474\
        );

    \I__4948\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22474\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__22500\,
            I => \N__22469\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__22497\,
            I => \N__22469\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__22494\,
            I => \N__22466\
        );

    \I__4944\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22461\
        );

    \I__4943\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22461\
        );

    \I__4942\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22458\
        );

    \I__4941\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22455\
        );

    \I__4940\ : CascadeMux
    port map (
            O => \N__22489\,
            I => \N__22452\
        );

    \I__4939\ : Span4Mux_s3_v
    port map (
            O => \N__22486\,
            I => \N__22443\
        );

    \I__4938\ : Span4Mux_s3_v
    port map (
            O => \N__22481\,
            I => \N__22443\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__22474\,
            I => \N__22443\
        );

    \I__4936\ : Span4Mux_s2_v
    port map (
            O => \N__22469\,
            I => \N__22440\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__22466\,
            I => \N__22435\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__22461\,
            I => \N__22435\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22430\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__22455\,
            I => \N__22430\
        );

    \I__4931\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22427\
        );

    \I__4930\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22422\
        );

    \I__4929\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22422\
        );

    \I__4928\ : Span4Mux_v
    port map (
            O => \N__22443\,
            I => \N__22417\
        );

    \I__4927\ : Span4Mux_v
    port map (
            O => \N__22440\,
            I => \N__22417\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__22435\,
            I => \N__22414\
        );

    \I__4925\ : Odrv12
    port map (
            O => \N__22430\,
            I => \tok.stall\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__22427\,
            I => \tok.stall\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__22422\,
            I => \tok.stall\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__22417\,
            I => \tok.stall\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__22414\,
            I => \tok.stall\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__22403\,
            I => \N__22397\
        );

    \I__4919\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22394\
        );

    \I__4918\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22390\
        );

    \I__4917\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22386\
        );

    \I__4916\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22383\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__22394\,
            I => \N__22380\
        );

    \I__4914\ : InMux
    port map (
            O => \N__22393\,
            I => \N__22377\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__22390\,
            I => \N__22370\
        );

    \I__4912\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22367\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__22386\,
            I => \N__22361\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22361\
        );

    \I__4909\ : Span4Mux_v
    port map (
            O => \N__22380\,
            I => \N__22358\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__22377\,
            I => \N__22355\
        );

    \I__4907\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22350\
        );

    \I__4906\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22350\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__22374\,
            I => \N__22346\
        );

    \I__4904\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22343\
        );

    \I__4903\ : Span4Mux_v
    port map (
            O => \N__22370\,
            I => \N__22338\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__22367\,
            I => \N__22338\
        );

    \I__4901\ : InMux
    port map (
            O => \N__22366\,
            I => \N__22335\
        );

    \I__4900\ : Span4Mux_v
    port map (
            O => \N__22361\,
            I => \N__22329\
        );

    \I__4899\ : Span4Mux_v
    port map (
            O => \N__22358\,
            I => \N__22322\
        );

    \I__4898\ : Span4Mux_s2_v
    port map (
            O => \N__22355\,
            I => \N__22322\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__22350\,
            I => \N__22322\
        );

    \I__4896\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22317\
        );

    \I__4895\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22317\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__22343\,
            I => \N__22312\
        );

    \I__4893\ : Span4Mux_h
    port map (
            O => \N__22338\,
            I => \N__22312\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__22335\,
            I => \N__22309\
        );

    \I__4891\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22304\
        );

    \I__4890\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22304\
        );

    \I__4889\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22301\
        );

    \I__4888\ : Span4Mux_h
    port map (
            O => \N__22329\,
            I => \N__22298\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__22322\,
            I => \tok.A_low_5\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__22317\,
            I => \tok.A_low_5\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__22312\,
            I => \tok.A_low_5\
        );

    \I__4884\ : Odrv12
    port map (
            O => \N__22309\,
            I => \tok.A_low_5\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__22304\,
            I => \tok.A_low_5\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__22301\,
            I => \tok.A_low_5\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__22298\,
            I => \tok.A_low_5\
        );

    \I__4880\ : CascadeMux
    port map (
            O => \N__22283\,
            I => \N__22278\
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__22282\,
            I => \N__22274\
        );

    \I__4878\ : CascadeMux
    port map (
            O => \N__22281\,
            I => \N__22269\
        );

    \I__4877\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22266\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__22277\,
            I => \N__22263\
        );

    \I__4875\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22254\
        );

    \I__4874\ : InMux
    port map (
            O => \N__22273\,
            I => \N__22254\
        );

    \I__4873\ : InMux
    port map (
            O => \N__22272\,
            I => \N__22254\
        );

    \I__4872\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22251\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__22266\,
            I => \N__22248\
        );

    \I__4870\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22245\
        );

    \I__4869\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22240\
        );

    \I__4868\ : InMux
    port map (
            O => \N__22261\,
            I => \N__22240\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__22254\,
            I => \N__22232\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__22251\,
            I => \N__22232\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__22248\,
            I => \N__22229\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__22245\,
            I => \N__22226\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__22240\,
            I => \N__22223\
        );

    \I__4862\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22216\
        );

    \I__4861\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22216\
        );

    \I__4860\ : InMux
    port map (
            O => \N__22237\,
            I => \N__22216\
        );

    \I__4859\ : Span12Mux_s6_h
    port map (
            O => \N__22232\,
            I => \N__22213\
        );

    \I__4858\ : Span4Mux_v
    port map (
            O => \N__22229\,
            I => \N__22210\
        );

    \I__4857\ : Span4Mux_s3_v
    port map (
            O => \N__22226\,
            I => \N__22205\
        );

    \I__4856\ : Span4Mux_h
    port map (
            O => \N__22223\,
            I => \N__22205\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__22216\,
            I => \tok.search_clk\
        );

    \I__4854\ : Odrv12
    port map (
            O => \N__22213\,
            I => \tok.search_clk\
        );

    \I__4853\ : Odrv4
    port map (
            O => \N__22210\,
            I => \tok.search_clk\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__22205\,
            I => \tok.search_clk\
        );

    \I__4851\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__22193\,
            I => \tok.n33_adj_817\
        );

    \I__4849\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__4847\ : Odrv12
    port map (
            O => \N__22184\,
            I => \tok.n27_adj_868\
        );

    \I__4846\ : InMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__22178\,
            I => \N__22172\
        );

    \I__4844\ : InMux
    port map (
            O => \N__22177\,
            I => \N__22169\
        );

    \I__4843\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22164\
        );

    \I__4842\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22164\
        );

    \I__4841\ : Span4Mux_h
    port map (
            O => \N__22172\,
            I => \N__22161\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22158\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__22164\,
            I => \N__22155\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__22161\,
            I => \tok.n82\
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__22158\,
            I => \tok.n82\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__22155\,
            I => \tok.n82\
        );

    \I__4835\ : InMux
    port map (
            O => \N__22148\,
            I => \N__22145\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__4833\ : Span4Mux_h
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__4832\ : Span4Mux_h
    port map (
            O => \N__22139\,
            I => \N__22134\
        );

    \I__4831\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22129\
        );

    \I__4830\ : InMux
    port map (
            O => \N__22137\,
            I => \N__22129\
        );

    \I__4829\ : Odrv4
    port map (
            O => \N__22134\,
            I => capture_5
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__22129\,
            I => capture_5
        );

    \I__4827\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22118\
        );

    \I__4826\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22115\
        );

    \I__4825\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22109\
        );

    \I__4824\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22106\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__22118\,
            I => \N__22103\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__22115\,
            I => \N__22098\
        );

    \I__4821\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22095\
        );

    \I__4820\ : InMux
    port map (
            O => \N__22113\,
            I => \N__22092\
        );

    \I__4819\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22089\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__22109\,
            I => \N__22086\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__22106\,
            I => \N__22083\
        );

    \I__4816\ : Span4Mux_h
    port map (
            O => \N__22103\,
            I => \N__22080\
        );

    \I__4815\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22075\
        );

    \I__4814\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22075\
        );

    \I__4813\ : Span4Mux_v
    port map (
            O => \N__22098\,
            I => \N__22072\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__22095\,
            I => \N__22069\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__22092\,
            I => \N__22064\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22064\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__22086\,
            I => \N__22061\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__22083\,
            I => \N__22058\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__22080\,
            I => \N__22053\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__22075\,
            I => \N__22053\
        );

    \I__4805\ : Span4Mux_h
    port map (
            O => \N__22072\,
            I => \N__22046\
        );

    \I__4804\ : Span4Mux_v
    port map (
            O => \N__22069\,
            I => \N__22046\
        );

    \I__4803\ : Span4Mux_h
    port map (
            O => \N__22064\,
            I => \N__22046\
        );

    \I__4802\ : Span4Mux_h
    port map (
            O => \N__22061\,
            I => \N__22043\
        );

    \I__4801\ : Span4Mux_v
    port map (
            O => \N__22058\,
            I => \N__22038\
        );

    \I__4800\ : Span4Mux_v
    port map (
            O => \N__22053\,
            I => \N__22038\
        );

    \I__4799\ : Span4Mux_h
    port map (
            O => \N__22046\,
            I => \N__22035\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__22043\,
            I => \rx_data_7__N_511\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__22038\,
            I => \rx_data_7__N_511\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__22035\,
            I => \rx_data_7__N_511\
        );

    \I__4795\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__4793\ : Odrv4
    port map (
            O => \N__22022\,
            I => \tok.n13_adj_816\
        );

    \I__4792\ : InMux
    port map (
            O => \N__22019\,
            I => \tok.n3902\
        );

    \I__4791\ : InMux
    port map (
            O => \N__22016\,
            I => \N__22013\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__22013\,
            I => \N__22010\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__22010\,
            I => \tok.n2_adj_811\
        );

    \I__4788\ : InMux
    port map (
            O => \N__22007\,
            I => \tok.n3903\
        );

    \I__4787\ : InMux
    port map (
            O => \N__22004\,
            I => \N__22001\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__22001\,
            I => \tok.n26_adj_808\
        );

    \I__4785\ : InMux
    port map (
            O => \N__21998\,
            I => \tok.n3904\
        );

    \I__4784\ : InMux
    port map (
            O => \N__21995\,
            I => \tok.n3905\
        );

    \I__4783\ : InMux
    port map (
            O => \N__21992\,
            I => \tok.n3906\
        );

    \I__4782\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21982\
        );

    \I__4781\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21978\
        );

    \I__4780\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21973\
        );

    \I__4779\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21968\
        );

    \I__4778\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21964\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__21982\,
            I => \N__21961\
        );

    \I__4776\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21958\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__21978\,
            I => \N__21954\
        );

    \I__4774\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21949\
        );

    \I__4773\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21949\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__21973\,
            I => \N__21946\
        );

    \I__4771\ : InMux
    port map (
            O => \N__21972\,
            I => \N__21943\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__21971\,
            I => \N__21939\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__21968\,
            I => \N__21934\
        );

    \I__4768\ : InMux
    port map (
            O => \N__21967\,
            I => \N__21931\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__21964\,
            I => \N__21924\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__21961\,
            I => \N__21924\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__21958\,
            I => \N__21924\
        );

    \I__4764\ : InMux
    port map (
            O => \N__21957\,
            I => \N__21921\
        );

    \I__4763\ : Span4Mux_v
    port map (
            O => \N__21954\,
            I => \N__21916\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__21949\,
            I => \N__21916\
        );

    \I__4761\ : Span4Mux_h
    port map (
            O => \N__21946\,
            I => \N__21913\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__21943\,
            I => \N__21910\
        );

    \I__4759\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21907\
        );

    \I__4758\ : InMux
    port map (
            O => \N__21939\,
            I => \N__21904\
        );

    \I__4757\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21901\
        );

    \I__4756\ : InMux
    port map (
            O => \N__21937\,
            I => \N__21898\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__21934\,
            I => \N__21893\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__21931\,
            I => \N__21893\
        );

    \I__4753\ : Span4Mux_h
    port map (
            O => \N__21924\,
            I => \N__21890\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__21921\,
            I => \N__21885\
        );

    \I__4751\ : Span4Mux_h
    port map (
            O => \N__21916\,
            I => \N__21885\
        );

    \I__4750\ : Odrv4
    port map (
            O => \N__21913\,
            I => \tok.A_low_2\
        );

    \I__4749\ : Odrv12
    port map (
            O => \N__21910\,
            I => \tok.A_low_2\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__21907\,
            I => \tok.A_low_2\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__21904\,
            I => \tok.A_low_2\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__21901\,
            I => \tok.A_low_2\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__21898\,
            I => \tok.A_low_2\
        );

    \I__4744\ : Odrv4
    port map (
            O => \N__21893\,
            I => \tok.A_low_2\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__21890\,
            I => \tok.A_low_2\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__21885\,
            I => \tok.A_low_2\
        );

    \I__4741\ : InMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__21863\,
            I => \N__21860\
        );

    \I__4739\ : Span4Mux_h
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__21857\,
            I => \tok.n210\
        );

    \I__4737\ : InMux
    port map (
            O => \N__21854\,
            I => \tok.n3907\
        );

    \I__4736\ : InMux
    port map (
            O => \N__21851\,
            I => \N__21847\
        );

    \I__4735\ : InMux
    port map (
            O => \N__21850\,
            I => \N__21842\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21836\
        );

    \I__4733\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21833\
        );

    \I__4732\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21828\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__21842\,
            I => \N__21825\
        );

    \I__4730\ : InMux
    port map (
            O => \N__21841\,
            I => \N__21820\
        );

    \I__4729\ : InMux
    port map (
            O => \N__21840\,
            I => \N__21817\
        );

    \I__4728\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21814\
        );

    \I__4727\ : Span4Mux_v
    port map (
            O => \N__21836\,
            I => \N__21808\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__21833\,
            I => \N__21808\
        );

    \I__4725\ : InMux
    port map (
            O => \N__21832\,
            I => \N__21803\
        );

    \I__4724\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21803\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__21828\,
            I => \N__21800\
        );

    \I__4722\ : Span4Mux_v
    port map (
            O => \N__21825\,
            I => \N__21797\
        );

    \I__4721\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21791\
        );

    \I__4720\ : InMux
    port map (
            O => \N__21823\,
            I => \N__21788\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__21820\,
            I => \N__21785\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__21817\,
            I => \N__21782\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__21814\,
            I => \N__21779\
        );

    \I__4716\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21776\
        );

    \I__4715\ : Span4Mux_h
    port map (
            O => \N__21808\,
            I => \N__21773\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__21803\,
            I => \N__21770\
        );

    \I__4713\ : Span4Mux_h
    port map (
            O => \N__21800\,
            I => \N__21767\
        );

    \I__4712\ : Sp12to4
    port map (
            O => \N__21797\,
            I => \N__21764\
        );

    \I__4711\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21761\
        );

    \I__4710\ : InMux
    port map (
            O => \N__21795\,
            I => \N__21758\
        );

    \I__4709\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21755\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__21791\,
            I => \N__21752\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__21788\,
            I => \N__21743\
        );

    \I__4706\ : Span4Mux_h
    port map (
            O => \N__21785\,
            I => \N__21743\
        );

    \I__4705\ : Span4Mux_h
    port map (
            O => \N__21782\,
            I => \N__21743\
        );

    \I__4704\ : Span4Mux_v
    port map (
            O => \N__21779\,
            I => \N__21743\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__21776\,
            I => \N__21736\
        );

    \I__4702\ : Span4Mux_v
    port map (
            O => \N__21773\,
            I => \N__21736\
        );

    \I__4701\ : Span4Mux_h
    port map (
            O => \N__21770\,
            I => \N__21736\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__21767\,
            I => \tok.A_low_3\
        );

    \I__4699\ : Odrv12
    port map (
            O => \N__21764\,
            I => \tok.A_low_3\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__21761\,
            I => \tok.A_low_3\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__21758\,
            I => \tok.A_low_3\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__21755\,
            I => \tok.A_low_3\
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__21752\,
            I => \tok.A_low_3\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__21743\,
            I => \tok.A_low_3\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__21736\,
            I => \tok.A_low_3\
        );

    \I__4692\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21713\
        );

    \I__4690\ : Span4Mux_h
    port map (
            O => \N__21713\,
            I => \N__21710\
        );

    \I__4689\ : Span4Mux_h
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__21707\,
            I => \tok.n209\
        );

    \I__4687\ : InMux
    port map (
            O => \N__21704\,
            I => \tok.n3908\
        );

    \I__4686\ : DummyBuf
    port map (
            O => \N__21701\,
            I => \N__21695\
        );

    \I__4685\ : DummyBuf
    port map (
            O => \N__21700\,
            I => \N__21692\
        );

    \I__4684\ : SRMux
    port map (
            O => \N__21699\,
            I => \N__21686\
        );

    \I__4683\ : SRMux
    port map (
            O => \N__21698\,
            I => \N__21682\
        );

    \I__4682\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21678\
        );

    \I__4681\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21675\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__21691\,
            I => \N__21672\
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__21690\,
            I => \N__21669\
        );

    \I__4678\ : CascadeMux
    port map (
            O => \N__21689\,
            I => \N__21666\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__21686\,
            I => \N__21662\
        );

    \I__4676\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21659\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__21682\,
            I => \N__21656\
        );

    \I__4674\ : SRMux
    port map (
            O => \N__21681\,
            I => \N__21653\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__21678\,
            I => \N__21650\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__21675\,
            I => \N__21647\
        );

    \I__4671\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21644\
        );

    \I__4670\ : InMux
    port map (
            O => \N__21669\,
            I => \N__21639\
        );

    \I__4669\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21639\
        );

    \I__4668\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21636\
        );

    \I__4667\ : Span4Mux_v
    port map (
            O => \N__21662\,
            I => \N__21633\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__21659\,
            I => \N__21630\
        );

    \I__4665\ : Span4Mux_v
    port map (
            O => \N__21656\,
            I => \N__21625\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__21653\,
            I => \N__21625\
        );

    \I__4663\ : Span4Mux_s3_v
    port map (
            O => \N__21650\,
            I => \N__21620\
        );

    \I__4662\ : Span4Mux_s3_v
    port map (
            O => \N__21647\,
            I => \N__21620\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__21644\,
            I => \N__21617\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__21639\,
            I => \N__21614\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__21636\,
            I => \N__21611\
        );

    \I__4658\ : Span4Mux_h
    port map (
            O => \N__21633\,
            I => \N__21607\
        );

    \I__4657\ : Span4Mux_v
    port map (
            O => \N__21630\,
            I => \N__21604\
        );

    \I__4656\ : Span4Mux_v
    port map (
            O => \N__21625\,
            I => \N__21601\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__21620\,
            I => \N__21598\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__21617\,
            I => \N__21591\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__21614\,
            I => \N__21591\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__21611\,
            I => \N__21591\
        );

    \I__4651\ : InMux
    port map (
            O => \N__21610\,
            I => \N__21588\
        );

    \I__4650\ : Span4Mux_h
    port map (
            O => \N__21607\,
            I => \N__21585\
        );

    \I__4649\ : Span4Mux_h
    port map (
            O => \N__21604\,
            I => \N__21582\
        );

    \I__4648\ : Span4Mux_s2_v
    port map (
            O => \N__21601\,
            I => \N__21579\
        );

    \I__4647\ : Span4Mux_v
    port map (
            O => \N__21598\,
            I => \N__21572\
        );

    \I__4646\ : Span4Mux_h
    port map (
            O => \N__21591\,
            I => \N__21572\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__21588\,
            I => \N__21572\
        );

    \I__4644\ : Odrv4
    port map (
            O => \N__21585\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4643\ : Odrv4
    port map (
            O => \N__21582\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__21579\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__21572\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4640\ : InMux
    port map (
            O => \N__21563\,
            I => \bfn_9_12_0_\
        );

    \I__4639\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21557\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__21557\,
            I => \tok.n2598\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__21554\,
            I => \tok.n5_adj_837_cascade_\
        );

    \I__4636\ : CascadeMux
    port map (
            O => \N__21551\,
            I => \N__21547\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__21550\,
            I => \N__21541\
        );

    \I__4634\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21535\
        );

    \I__4633\ : InMux
    port map (
            O => \N__21546\,
            I => \N__21532\
        );

    \I__4632\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21529\
        );

    \I__4631\ : CascadeMux
    port map (
            O => \N__21544\,
            I => \N__21526\
        );

    \I__4630\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21523\
        );

    \I__4629\ : CascadeMux
    port map (
            O => \N__21540\,
            I => \N__21520\
        );

    \I__4628\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21517\
        );

    \I__4627\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21514\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__21535\,
            I => \N__21511\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__21532\,
            I => \N__21506\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__21529\,
            I => \N__21506\
        );

    \I__4623\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21503\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__21523\,
            I => \N__21500\
        );

    \I__4621\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21497\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__21517\,
            I => \N__21492\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__21514\,
            I => \N__21492\
        );

    \I__4618\ : Span4Mux_h
    port map (
            O => \N__21511\,
            I => \N__21484\
        );

    \I__4617\ : Span4Mux_v
    port map (
            O => \N__21506\,
            I => \N__21484\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__21503\,
            I => \N__21484\
        );

    \I__4615\ : Span4Mux_h
    port map (
            O => \N__21500\,
            I => \N__21477\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__21497\,
            I => \N__21477\
        );

    \I__4613\ : Span4Mux_s3_v
    port map (
            O => \N__21492\,
            I => \N__21477\
        );

    \I__4612\ : InMux
    port map (
            O => \N__21491\,
            I => \N__21474\
        );

    \I__4611\ : Span4Mux_v
    port map (
            O => \N__21484\,
            I => \N__21471\
        );

    \I__4610\ : Span4Mux_v
    port map (
            O => \N__21477\,
            I => \N__21468\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__21474\,
            I => \tok.S_3\
        );

    \I__4608\ : Odrv4
    port map (
            O => \N__21471\,
            I => \tok.S_3\
        );

    \I__4607\ : Odrv4
    port map (
            O => \N__21468\,
            I => \tok.S_3\
        );

    \I__4606\ : InMux
    port map (
            O => \N__21461\,
            I => \N__21458\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__21458\,
            I => \N__21455\
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__21455\,
            I => \tok.n23_adj_788\
        );

    \I__4603\ : CascadeMux
    port map (
            O => \N__21452\,
            I => \tok.n10_adj_838_cascade_\
        );

    \I__4602\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21446\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__21446\,
            I => \N__21443\
        );

    \I__4600\ : Odrv4
    port map (
            O => \N__21443\,
            I => \tok.n12_adj_840\
        );

    \I__4599\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__21437\,
            I => \N__21431\
        );

    \I__4597\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21425\
        );

    \I__4596\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21422\
        );

    \I__4595\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21419\
        );

    \I__4594\ : Span4Mux_v
    port map (
            O => \N__21431\,
            I => \N__21416\
        );

    \I__4593\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21411\
        );

    \I__4592\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21411\
        );

    \I__4591\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21407\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__21425\,
            I => \N__21404\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__21422\,
            I => \N__21397\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__21419\,
            I => \N__21394\
        );

    \I__4587\ : Span4Mux_h
    port map (
            O => \N__21416\,
            I => \N__21389\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__21411\,
            I => \N__21389\
        );

    \I__4585\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21386\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__21407\,
            I => \N__21383\
        );

    \I__4583\ : Span4Mux_h
    port map (
            O => \N__21404\,
            I => \N__21380\
        );

    \I__4582\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21375\
        );

    \I__4581\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21375\
        );

    \I__4580\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21370\
        );

    \I__4579\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21370\
        );

    \I__4578\ : Span4Mux_h
    port map (
            O => \N__21397\,
            I => \N__21363\
        );

    \I__4577\ : Span4Mux_v
    port map (
            O => \N__21394\,
            I => \N__21363\
        );

    \I__4576\ : Span4Mux_v
    port map (
            O => \N__21389\,
            I => \N__21363\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__21386\,
            I => \N__21358\
        );

    \I__4574\ : Span4Mux_h
    port map (
            O => \N__21383\,
            I => \N__21358\
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__21380\,
            I => \tok.n57\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__21375\,
            I => \tok.n57\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__21370\,
            I => \tok.n57\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__21363\,
            I => \tok.n57\
        );

    \I__4569\ : Odrv4
    port map (
            O => \N__21358\,
            I => \tok.n57\
        );

    \I__4568\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__21344\,
            I => \tok.n6_adj_835\
        );

    \I__4566\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21337\
        );

    \I__4565\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21334\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__21337\,
            I => \N__21331\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__21334\,
            I => uart_rx_data_6
        );

    \I__4562\ : Odrv12
    port map (
            O => \N__21331\,
            I => uart_rx_data_6
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__21326\,
            I => \tok.n109_cascade_\
        );

    \I__4560\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21316\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__21322\,
            I => \N__21313\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__21321\,
            I => \N__21310\
        );

    \I__4557\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21307\
        );

    \I__4556\ : InMux
    port map (
            O => \N__21319\,
            I => \N__21304\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21300\
        );

    \I__4554\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21295\
        );

    \I__4553\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21292\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21287\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__21304\,
            I => \N__21287\
        );

    \I__4550\ : CascadeMux
    port map (
            O => \N__21303\,
            I => \N__21284\
        );

    \I__4549\ : Span4Mux_v
    port map (
            O => \N__21300\,
            I => \N__21281\
        );

    \I__4548\ : InMux
    port map (
            O => \N__21299\,
            I => \N__21278\
        );

    \I__4547\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21275\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__21295\,
            I => \N__21270\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__21292\,
            I => \N__21270\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__21287\,
            I => \N__21266\
        );

    \I__4543\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21263\
        );

    \I__4542\ : Span4Mux_h
    port map (
            O => \N__21281\,
            I => \N__21258\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__21278\,
            I => \N__21258\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__21275\,
            I => \N__21253\
        );

    \I__4539\ : Span4Mux_h
    port map (
            O => \N__21270\,
            I => \N__21253\
        );

    \I__4538\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21250\
        );

    \I__4537\ : Sp12to4
    port map (
            O => \N__21266\,
            I => \N__21245\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__21263\,
            I => \N__21245\
        );

    \I__4535\ : Span4Mux_v
    port map (
            O => \N__21258\,
            I => \N__21240\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__21253\,
            I => \N__21240\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__21250\,
            I => \tok.S_6\
        );

    \I__4532\ : Odrv12
    port map (
            O => \N__21245\,
            I => \tok.S_6\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__21240\,
            I => \tok.S_6\
        );

    \I__4530\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21230\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__21230\,
            I => \N__21227\
        );

    \I__4528\ : Span4Mux_v
    port map (
            O => \N__21227\,
            I => \N__21224\
        );

    \I__4527\ : Odrv4
    port map (
            O => \N__21224\,
            I => \tok.n18_adj_782\
        );

    \I__4526\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__4524\ : Span4Mux_h
    port map (
            O => \N__21215\,
            I => \N__21211\
        );

    \I__4523\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21208\
        );

    \I__4522\ : Span4Mux_h
    port map (
            O => \N__21211\,
            I => \N__21202\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__21208\,
            I => \N__21202\
        );

    \I__4520\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21199\
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__21202\,
            I => capture_4
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__21199\,
            I => capture_4
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__21194\,
            I => \N__21190\
        );

    \I__4516\ : InMux
    port map (
            O => \N__21193\,
            I => \N__21185\
        );

    \I__4515\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21185\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__21185\,
            I => uart_rx_data_3
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__21182\,
            I => \N__21177\
        );

    \I__4512\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21174\
        );

    \I__4511\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21170\
        );

    \I__4510\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21165\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__21174\,
            I => \N__21162\
        );

    \I__4508\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21159\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__21170\,
            I => \N__21155\
        );

    \I__4506\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21152\
        );

    \I__4505\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21149\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__21165\,
            I => \N__21146\
        );

    \I__4503\ : Span4Mux_h
    port map (
            O => \N__21162\,
            I => \N__21142\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__21159\,
            I => \N__21139\
        );

    \I__4501\ : InMux
    port map (
            O => \N__21158\,
            I => \N__21136\
        );

    \I__4500\ : Span4Mux_v
    port map (
            O => \N__21155\,
            I => \N__21129\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__21152\,
            I => \N__21129\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__21149\,
            I => \N__21129\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__21146\,
            I => \N__21126\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__21145\,
            I => \N__21123\
        );

    \I__4495\ : Span4Mux_s0_h
    port map (
            O => \N__21142\,
            I => \N__21118\
        );

    \I__4494\ : Span4Mux_h
    port map (
            O => \N__21139\,
            I => \N__21118\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__21136\,
            I => \N__21115\
        );

    \I__4492\ : Span4Mux_v
    port map (
            O => \N__21129\,
            I => \N__21112\
        );

    \I__4491\ : Span4Mux_h
    port map (
            O => \N__21126\,
            I => \N__21109\
        );

    \I__4490\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21106\
        );

    \I__4489\ : Span4Mux_v
    port map (
            O => \N__21118\,
            I => \N__21103\
        );

    \I__4488\ : Span4Mux_v
    port map (
            O => \N__21115\,
            I => \N__21096\
        );

    \I__4487\ : Span4Mux_h
    port map (
            O => \N__21112\,
            I => \N__21096\
        );

    \I__4486\ : Span4Mux_h
    port map (
            O => \N__21109\,
            I => \N__21096\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__21106\,
            I => \tok.S_9\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__21103\,
            I => \tok.S_9\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__21096\,
            I => \tok.S_9\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__21089\,
            I => \N__21086\
        );

    \I__4481\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21083\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__4479\ : Span4Mux_v
    port map (
            O => \N__21080\,
            I => \N__21077\
        );

    \I__4478\ : Span4Mux_h
    port map (
            O => \N__21077\,
            I => \N__21074\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__21074\,
            I => \tok.n21\
        );

    \I__4476\ : InMux
    port map (
            O => \N__21071\,
            I => \tok.n3933\
        );

    \I__4475\ : InMux
    port map (
            O => \N__21068\,
            I => \N__21064\
        );

    \I__4474\ : InMux
    port map (
            O => \N__21067\,
            I => \N__21061\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__21064\,
            I => \N__21056\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__21061\,
            I => \N__21051\
        );

    \I__4471\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21048\
        );

    \I__4470\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21044\
        );

    \I__4469\ : Span4Mux_v
    port map (
            O => \N__21056\,
            I => \N__21041\
        );

    \I__4468\ : InMux
    port map (
            O => \N__21055\,
            I => \N__21038\
        );

    \I__4467\ : InMux
    port map (
            O => \N__21054\,
            I => \N__21035\
        );

    \I__4466\ : Span4Mux_v
    port map (
            O => \N__21051\,
            I => \N__21026\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__21048\,
            I => \N__21023\
        );

    \I__4464\ : InMux
    port map (
            O => \N__21047\,
            I => \N__21020\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__21044\,
            I => \N__21017\
        );

    \I__4462\ : Span4Mux_h
    port map (
            O => \N__21041\,
            I => \N__21012\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__21038\,
            I => \N__21012\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__21035\,
            I => \N__21009\
        );

    \I__4459\ : InMux
    port map (
            O => \N__21034\,
            I => \N__21006\
        );

    \I__4458\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21001\
        );

    \I__4457\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21001\
        );

    \I__4456\ : InMux
    port map (
            O => \N__21031\,
            I => \N__20994\
        );

    \I__4455\ : InMux
    port map (
            O => \N__21030\,
            I => \N__20994\
        );

    \I__4454\ : InMux
    port map (
            O => \N__21029\,
            I => \N__20994\
        );

    \I__4453\ : Span4Mux_h
    port map (
            O => \N__21026\,
            I => \N__20987\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__21023\,
            I => \N__20987\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__21020\,
            I => \N__20987\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__21017\,
            I => \N__20982\
        );

    \I__4449\ : Span4Mux_h
    port map (
            O => \N__21012\,
            I => \N__20982\
        );

    \I__4448\ : Span4Mux_h
    port map (
            O => \N__21009\,
            I => \N__20977\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__21006\,
            I => \N__20977\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__21001\,
            I => \tok.n58\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__20994\,
            I => \tok.n58\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__20987\,
            I => \tok.n58\
        );

    \I__4443\ : Odrv4
    port map (
            O => \N__20982\,
            I => \tok.n58\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__20977\,
            I => \tok.n58\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__20966\,
            I => \N__20962\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__20965\,
            I => \N__20959\
        );

    \I__4439\ : InMux
    port map (
            O => \N__20962\,
            I => \N__20955\
        );

    \I__4438\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20949\
        );

    \I__4437\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20944\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__20955\,
            I => \N__20941\
        );

    \I__4435\ : InMux
    port map (
            O => \N__20954\,
            I => \N__20938\
        );

    \I__4434\ : InMux
    port map (
            O => \N__20953\,
            I => \N__20935\
        );

    \I__4433\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20932\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20929\
        );

    \I__4431\ : CascadeMux
    port map (
            O => \N__20948\,
            I => \N__20926\
        );

    \I__4430\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20923\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__20944\,
            I => \N__20918\
        );

    \I__4428\ : Span4Mux_h
    port map (
            O => \N__20941\,
            I => \N__20918\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__20938\,
            I => \N__20913\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__20935\,
            I => \N__20913\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__20932\,
            I => \N__20908\
        );

    \I__4424\ : Span4Mux_h
    port map (
            O => \N__20929\,
            I => \N__20908\
        );

    \I__4423\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20905\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__20923\,
            I => \N__20902\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__20918\,
            I => \N__20899\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__20913\,
            I => \N__20896\
        );

    \I__4419\ : Span4Mux_h
    port map (
            O => \N__20908\,
            I => \N__20893\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__20905\,
            I => \tok.S_10\
        );

    \I__4417\ : Odrv12
    port map (
            O => \N__20902\,
            I => \tok.S_10\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__20899\,
            I => \tok.S_10\
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__20896\,
            I => \tok.S_10\
        );

    \I__4414\ : Odrv4
    port map (
            O => \N__20893\,
            I => \tok.S_10\
        );

    \I__4413\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__20876\,
            I => \tok.n5_adj_668\
        );

    \I__4410\ : InMux
    port map (
            O => \N__20873\,
            I => \tok.n3934\
        );

    \I__4409\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20864\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__20869\,
            I => \N__20861\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__20868\,
            I => \N__20858\
        );

    \I__4406\ : InMux
    port map (
            O => \N__20867\,
            I => \N__20854\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__20864\,
            I => \N__20850\
        );

    \I__4404\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20847\
        );

    \I__4403\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20844\
        );

    \I__4402\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20839\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__20854\,
            I => \N__20836\
        );

    \I__4400\ : InMux
    port map (
            O => \N__20853\,
            I => \N__20833\
        );

    \I__4399\ : Span4Mux_s3_v
    port map (
            O => \N__20850\,
            I => \N__20828\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__20847\,
            I => \N__20828\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__20844\,
            I => \N__20825\
        );

    \I__4396\ : CascadeMux
    port map (
            O => \N__20843\,
            I => \N__20822\
        );

    \I__4395\ : InMux
    port map (
            O => \N__20842\,
            I => \N__20819\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__20839\,
            I => \N__20816\
        );

    \I__4393\ : Span4Mux_s3_v
    port map (
            O => \N__20836\,
            I => \N__20811\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20811\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__20828\,
            I => \N__20808\
        );

    \I__4390\ : Span4Mux_v
    port map (
            O => \N__20825\,
            I => \N__20805\
        );

    \I__4389\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20802\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__20819\,
            I => \N__20799\
        );

    \I__4387\ : Span4Mux_h
    port map (
            O => \N__20816\,
            I => \N__20792\
        );

    \I__4386\ : Span4Mux_v
    port map (
            O => \N__20811\,
            I => \N__20792\
        );

    \I__4385\ : Span4Mux_h
    port map (
            O => \N__20808\,
            I => \N__20792\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__20805\,
            I => \N__20789\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__20802\,
            I => \N__20784\
        );

    \I__4382\ : Span4Mux_v
    port map (
            O => \N__20799\,
            I => \N__20784\
        );

    \I__4381\ : Span4Mux_h
    port map (
            O => \N__20792\,
            I => \N__20781\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__20789\,
            I => \tok.S_11\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__20784\,
            I => \tok.S_11\
        );

    \I__4378\ : Odrv4
    port map (
            O => \N__20781\,
            I => \tok.S_11\
        );

    \I__4377\ : InMux
    port map (
            O => \N__20774\,
            I => \N__20771\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__20771\,
            I => \N__20768\
        );

    \I__4375\ : Odrv12
    port map (
            O => \N__20768\,
            I => \tok.n5_adj_690\
        );

    \I__4374\ : InMux
    port map (
            O => \N__20765\,
            I => \tok.n3935\
        );

    \I__4373\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20757\
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__20761\,
            I => \N__20754\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__20760\,
            I => \N__20748\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__20757\,
            I => \N__20745\
        );

    \I__4369\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20742\
        );

    \I__4368\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20739\
        );

    \I__4367\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20736\
        );

    \I__4366\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20733\
        );

    \I__4365\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20729\
        );

    \I__4364\ : Span4Mux_v
    port map (
            O => \N__20745\,
            I => \N__20724\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__20742\,
            I => \N__20724\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__20739\,
            I => \N__20716\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__20736\,
            I => \N__20716\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__20733\,
            I => \N__20716\
        );

    \I__4359\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20713\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__20729\,
            I => \N__20710\
        );

    \I__4357\ : Span4Mux_v
    port map (
            O => \N__20724\,
            I => \N__20707\
        );

    \I__4356\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20704\
        );

    \I__4355\ : Span12Mux_v
    port map (
            O => \N__20716\,
            I => \N__20701\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__20713\,
            I => \N__20696\
        );

    \I__4353\ : Span12Mux_s8_h
    port map (
            O => \N__20710\,
            I => \N__20696\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__20707\,
            I => \N__20693\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__20704\,
            I => \tok.S_12\
        );

    \I__4350\ : Odrv12
    port map (
            O => \N__20701\,
            I => \tok.S_12\
        );

    \I__4349\ : Odrv12
    port map (
            O => \N__20696\,
            I => \tok.S_12\
        );

    \I__4348\ : Odrv4
    port map (
            O => \N__20693\,
            I => \tok.S_12\
        );

    \I__4347\ : InMux
    port map (
            O => \N__20684\,
            I => \tok.n3936\
        );

    \I__4346\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20673\
        );

    \I__4345\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20670\
        );

    \I__4344\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20667\
        );

    \I__4343\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20664\
        );

    \I__4342\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20661\
        );

    \I__4341\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20658\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__20673\,
            I => \N__20653\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__20670\,
            I => \N__20653\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__20667\,
            I => \N__20647\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__20664\,
            I => \N__20647\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__20661\,
            I => \N__20644\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20638\
        );

    \I__4334\ : Span4Mux_v
    port map (
            O => \N__20653\,
            I => \N__20635\
        );

    \I__4333\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20632\
        );

    \I__4332\ : Span4Mux_v
    port map (
            O => \N__20647\,
            I => \N__20627\
        );

    \I__4331\ : Span4Mux_h
    port map (
            O => \N__20644\,
            I => \N__20627\
        );

    \I__4330\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20622\
        );

    \I__4329\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20622\
        );

    \I__4328\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20619\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__20638\,
            I => \N__20616\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__20635\,
            I => \N__20611\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__20632\,
            I => \N__20611\
        );

    \I__4324\ : Span4Mux_v
    port map (
            O => \N__20627\,
            I => \N__20608\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__20622\,
            I => \tok.n55\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__20619\,
            I => \tok.n55\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__20616\,
            I => \tok.n55\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__20611\,
            I => \tok.n55\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__20608\,
            I => \tok.n55\
        );

    \I__4318\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20592\
        );

    \I__4317\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20589\
        );

    \I__4316\ : CascadeMux
    port map (
            O => \N__20595\,
            I => \N__20584\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__20592\,
            I => \N__20580\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__20589\,
            I => \N__20577\
        );

    \I__4313\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20574\
        );

    \I__4312\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20571\
        );

    \I__4311\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20568\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__20583\,
            I => \N__20565\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__20580\,
            I => \N__20554\
        );

    \I__4308\ : Span4Mux_s3_h
    port map (
            O => \N__20577\,
            I => \N__20554\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20554\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__20571\,
            I => \N__20554\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__20568\,
            I => \N__20551\
        );

    \I__4304\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20548\
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__20564\,
            I => \N__20545\
        );

    \I__4302\ : InMux
    port map (
            O => \N__20563\,
            I => \N__20542\
        );

    \I__4301\ : Span4Mux_h
    port map (
            O => \N__20554\,
            I => \N__20537\
        );

    \I__4300\ : Span4Mux_h
    port map (
            O => \N__20551\,
            I => \N__20537\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__20548\,
            I => \N__20534\
        );

    \I__4298\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20531\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20528\
        );

    \I__4296\ : Span4Mux_v
    port map (
            O => \N__20537\,
            I => \N__20525\
        );

    \I__4295\ : Span4Mux_h
    port map (
            O => \N__20534\,
            I => \N__20522\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__20531\,
            I => \tok.S_13\
        );

    \I__4293\ : Odrv12
    port map (
            O => \N__20528\,
            I => \tok.S_13\
        );

    \I__4292\ : Odrv4
    port map (
            O => \N__20525\,
            I => \tok.S_13\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__20522\,
            I => \tok.S_13\
        );

    \I__4290\ : InMux
    port map (
            O => \N__20513\,
            I => \tok.n3937\
        );

    \I__4289\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20502\
        );

    \I__4288\ : InMux
    port map (
            O => \N__20509\,
            I => \N__20499\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__20508\,
            I => \N__20496\
        );

    \I__4286\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20492\
        );

    \I__4285\ : InMux
    port map (
            O => \N__20506\,
            I => \N__20489\
        );

    \I__4284\ : InMux
    port map (
            O => \N__20505\,
            I => \N__20486\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__20502\,
            I => \N__20483\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__20499\,
            I => \N__20480\
        );

    \I__4281\ : InMux
    port map (
            O => \N__20496\,
            I => \N__20477\
        );

    \I__4280\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20474\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__20492\,
            I => \N__20471\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__20489\,
            I => \N__20468\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__20486\,
            I => \N__20465\
        );

    \I__4276\ : Span4Mux_h
    port map (
            O => \N__20483\,
            I => \N__20462\
        );

    \I__4275\ : Span4Mux_v
    port map (
            O => \N__20480\,
            I => \N__20457\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__20477\,
            I => \N__20457\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__20474\,
            I => \N__20453\
        );

    \I__4272\ : Span4Mux_v
    port map (
            O => \N__20471\,
            I => \N__20450\
        );

    \I__4271\ : Span4Mux_v
    port map (
            O => \N__20468\,
            I => \N__20445\
        );

    \I__4270\ : Span4Mux_v
    port map (
            O => \N__20465\,
            I => \N__20445\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__20462\,
            I => \N__20442\
        );

    \I__4268\ : Span4Mux_h
    port map (
            O => \N__20457\,
            I => \N__20439\
        );

    \I__4267\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20436\
        );

    \I__4266\ : Span4Mux_v
    port map (
            O => \N__20453\,
            I => \N__20433\
        );

    \I__4265\ : Span4Mux_v
    port map (
            O => \N__20450\,
            I => \N__20428\
        );

    \I__4264\ : Span4Mux_v
    port map (
            O => \N__20445\,
            I => \N__20428\
        );

    \I__4263\ : Span4Mux_h
    port map (
            O => \N__20442\,
            I => \N__20425\
        );

    \I__4262\ : Span4Mux_h
    port map (
            O => \N__20439\,
            I => \N__20422\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__20436\,
            I => \tok.S_14\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__20433\,
            I => \tok.S_14\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__20428\,
            I => \tok.S_14\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__20425\,
            I => \tok.S_14\
        );

    \I__4257\ : Odrv4
    port map (
            O => \N__20422\,
            I => \tok.S_14\
        );

    \I__4256\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__20408\,
            I => \tok.n5_adj_729\
        );

    \I__4254\ : InMux
    port map (
            O => \N__20405\,
            I => \tok.n3938\
        );

    \I__4253\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20396\
        );

    \I__4252\ : InMux
    port map (
            O => \N__20401\,
            I => \N__20391\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__20400\,
            I => \N__20388\
        );

    \I__4250\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20385\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__20396\,
            I => \N__20382\
        );

    \I__4248\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20379\
        );

    \I__4247\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20376\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__20391\,
            I => \N__20373\
        );

    \I__4245\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20370\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__20385\,
            I => \N__20365\
        );

    \I__4243\ : Span4Mux_v
    port map (
            O => \N__20382\,
            I => \N__20362\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__20379\,
            I => \N__20353\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__20376\,
            I => \N__20353\
        );

    \I__4240\ : Span4Mux_v
    port map (
            O => \N__20373\,
            I => \N__20353\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__20370\,
            I => \N__20353\
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__20369\,
            I => \N__20350\
        );

    \I__4237\ : InMux
    port map (
            O => \N__20368\,
            I => \N__20347\
        );

    \I__4236\ : Span4Mux_v
    port map (
            O => \N__20365\,
            I => \N__20344\
        );

    \I__4235\ : Span4Mux_h
    port map (
            O => \N__20362\,
            I => \N__20339\
        );

    \I__4234\ : Span4Mux_v
    port map (
            O => \N__20353\,
            I => \N__20339\
        );

    \I__4233\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20336\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__20347\,
            I => \N__20333\
        );

    \I__4231\ : Span4Mux_v
    port map (
            O => \N__20344\,
            I => \N__20328\
        );

    \I__4230\ : Span4Mux_v
    port map (
            O => \N__20339\,
            I => \N__20328\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__20336\,
            I => \tok.S_15\
        );

    \I__4228\ : Odrv12
    port map (
            O => \N__20333\,
            I => \tok.S_15\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__20328\,
            I => \tok.S_15\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__20321\,
            I => \N__20318\
        );

    \I__4225\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20315\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__20315\,
            I => \N__20306\
        );

    \I__4223\ : InMux
    port map (
            O => \N__20314\,
            I => \N__20302\
        );

    \I__4222\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20297\
        );

    \I__4221\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20297\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__20311\,
            I => \N__20294\
        );

    \I__4219\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20291\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__20309\,
            I => \N__20288\
        );

    \I__4217\ : Span4Mux_v
    port map (
            O => \N__20306\,
            I => \N__20284\
        );

    \I__4216\ : InMux
    port map (
            O => \N__20305\,
            I => \N__20281\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__20302\,
            I => \N__20277\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__20297\,
            I => \N__20274\
        );

    \I__4213\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20271\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__20291\,
            I => \N__20268\
        );

    \I__4211\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20265\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__20287\,
            I => \N__20262\
        );

    \I__4209\ : Span4Mux_s3_h
    port map (
            O => \N__20284\,
            I => \N__20259\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__20281\,
            I => \N__20256\
        );

    \I__4207\ : InMux
    port map (
            O => \N__20280\,
            I => \N__20253\
        );

    \I__4206\ : Span4Mux_v
    port map (
            O => \N__20277\,
            I => \N__20246\
        );

    \I__4205\ : Span4Mux_s3_h
    port map (
            O => \N__20274\,
            I => \N__20246\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__20271\,
            I => \N__20246\
        );

    \I__4203\ : Span4Mux_s3_v
    port map (
            O => \N__20268\,
            I => \N__20241\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__20265\,
            I => \N__20241\
        );

    \I__4201\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20238\
        );

    \I__4200\ : Span4Mux_h
    port map (
            O => \N__20259\,
            I => \N__20235\
        );

    \I__4199\ : Span4Mux_v
    port map (
            O => \N__20256\,
            I => \N__20230\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__20253\,
            I => \N__20230\
        );

    \I__4197\ : Span4Mux_h
    port map (
            O => \N__20246\,
            I => \N__20225\
        );

    \I__4196\ : Span4Mux_v
    port map (
            O => \N__20241\,
            I => \N__20225\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__20238\,
            I => \tok.n53\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__20235\,
            I => \tok.n53\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__20230\,
            I => \tok.n53\
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__20225\,
            I => \tok.n53\
        );

    \I__4191\ : InMux
    port map (
            O => \N__20216\,
            I => \tok.n3939\
        );

    \I__4190\ : InMux
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__4188\ : Span4Mux_v
    port map (
            O => \N__20207\,
            I => \N__20204\
        );

    \I__4187\ : Sp12to4
    port map (
            O => \N__20204\,
            I => \N__20201\
        );

    \I__4186\ : Odrv12
    port map (
            O => \N__20201\,
            I => \tok.n5_adj_750\
        );

    \I__4185\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20192\
        );

    \I__4183\ : Span4Mux_v
    port map (
            O => \N__20192\,
            I => \N__20189\
        );

    \I__4182\ : Span4Mux_h
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__4181\ : Odrv4
    port map (
            O => \N__20186\,
            I => \tok.n6_adj_812\
        );

    \I__4180\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__20180\,
            I => \N__20177\
        );

    \I__4178\ : Span12Mux_s10_v
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__4177\ : Odrv12
    port map (
            O => \N__20174\,
            I => \tok.n9_adj_836\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__20171\,
            I => \N__20166\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__20170\,
            I => \N__20163\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__20169\,
            I => \N__20159\
        );

    \I__4173\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20156\
        );

    \I__4172\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20151\
        );

    \I__4171\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20147\
        );

    \I__4170\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20144\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__20156\,
            I => \N__20140\
        );

    \I__4168\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20137\
        );

    \I__4167\ : InMux
    port map (
            O => \N__20154\,
            I => \N__20134\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__20151\,
            I => \N__20131\
        );

    \I__4165\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20128\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__20147\,
            I => \N__20123\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20123\
        );

    \I__4162\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20120\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__20140\,
            I => \N__20117\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__20137\,
            I => \N__20114\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__20134\,
            I => \N__20106\
        );

    \I__4158\ : Span4Mux_v
    port map (
            O => \N__20131\,
            I => \N__20106\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__20128\,
            I => \N__20106\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__20123\,
            I => \N__20101\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__20120\,
            I => \N__20101\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__20117\,
            I => \N__20098\
        );

    \I__4153\ : Span4Mux_v
    port map (
            O => \N__20114\,
            I => \N__20095\
        );

    \I__4152\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20092\
        );

    \I__4151\ : Span4Mux_v
    port map (
            O => \N__20106\,
            I => \N__20087\
        );

    \I__4150\ : Span4Mux_h
    port map (
            O => \N__20101\,
            I => \N__20087\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__20098\,
            I => \tok.S_1\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__20095\,
            I => \tok.S_1\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__20092\,
            I => \tok.S_1\
        );

    \I__4146\ : Odrv4
    port map (
            O => \N__20087\,
            I => \tok.S_1\
        );

    \I__4145\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__20075\,
            I => \tok.n4_adj_790\
        );

    \I__4143\ : InMux
    port map (
            O => \N__20072\,
            I => \tok.n3925\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__20069\,
            I => \N__20065\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__20068\,
            I => \N__20061\
        );

    \I__4140\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20056\
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__20064\,
            I => \N__20053\
        );

    \I__4138\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20050\
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__20060\,
            I => \N__20047\
        );

    \I__4136\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20044\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__20056\,
            I => \N__20039\
        );

    \I__4134\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20036\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__20050\,
            I => \N__20032\
        );

    \I__4132\ : InMux
    port map (
            O => \N__20047\,
            I => \N__20029\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__20044\,
            I => \N__20025\
        );

    \I__4130\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20020\
        );

    \I__4129\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20020\
        );

    \I__4128\ : Span4Mux_h
    port map (
            O => \N__20039\,
            I => \N__20017\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__20036\,
            I => \N__20014\
        );

    \I__4126\ : InMux
    port map (
            O => \N__20035\,
            I => \N__20011\
        );

    \I__4125\ : Span4Mux_h
    port map (
            O => \N__20032\,
            I => \N__20006\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__20029\,
            I => \N__20006\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__20028\,
            I => \N__20003\
        );

    \I__4122\ : Span4Mux_h
    port map (
            O => \N__20025\,
            I => \N__19998\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__20020\,
            I => \N__19998\
        );

    \I__4120\ : Span4Mux_h
    port map (
            O => \N__20017\,
            I => \N__19991\
        );

    \I__4119\ : Span4Mux_v
    port map (
            O => \N__20014\,
            I => \N__19991\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__20011\,
            I => \N__19991\
        );

    \I__4117\ : Span4Mux_v
    port map (
            O => \N__20006\,
            I => \N__19988\
        );

    \I__4116\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19985\
        );

    \I__4115\ : Span4Mux_v
    port map (
            O => \N__19998\,
            I => \N__19982\
        );

    \I__4114\ : Span4Mux_v
    port map (
            O => \N__19991\,
            I => \N__19977\
        );

    \I__4113\ : Span4Mux_h
    port map (
            O => \N__19988\,
            I => \N__19977\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__19985\,
            I => \tok.S_2\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__19982\,
            I => \tok.S_2\
        );

    \I__4110\ : Odrv4
    port map (
            O => \N__19977\,
            I => \tok.S_2\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__4108\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__19964\,
            I => \tok.n5_adj_789\
        );

    \I__4106\ : InMux
    port map (
            O => \N__19961\,
            I => \tok.n3926\
        );

    \I__4105\ : InMux
    port map (
            O => \N__19958\,
            I => \tok.n3927\
        );

    \I__4104\ : InMux
    port map (
            O => \N__19955\,
            I => \tok.n3928\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__19952\,
            I => \N__19943\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__19951\,
            I => \N__19940\
        );

    \I__4101\ : CascadeMux
    port map (
            O => \N__19950\,
            I => \N__19937\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__19949\,
            I => \N__19934\
        );

    \I__4099\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19929\
        );

    \I__4098\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19929\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__19946\,
            I => \N__19926\
        );

    \I__4096\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19923\
        );

    \I__4095\ : InMux
    port map (
            O => \N__19940\,
            I => \N__19920\
        );

    \I__4094\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19916\
        );

    \I__4093\ : InMux
    port map (
            O => \N__19934\,
            I => \N__19913\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__19929\,
            I => \N__19910\
        );

    \I__4091\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19907\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__19923\,
            I => \N__19901\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__19920\,
            I => \N__19901\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__19919\,
            I => \N__19898\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__19916\,
            I => \N__19893\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__19913\,
            I => \N__19893\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__19910\,
            I => \N__19888\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19888\
        );

    \I__4083\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19885\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__19901\,
            I => \N__19882\
        );

    \I__4081\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19879\
        );

    \I__4080\ : Span12Mux_s9_v
    port map (
            O => \N__19893\,
            I => \N__19876\
        );

    \I__4079\ : Span4Mux_v
    port map (
            O => \N__19888\,
            I => \N__19869\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__19885\,
            I => \N__19869\
        );

    \I__4077\ : Span4Mux_h
    port map (
            O => \N__19882\,
            I => \N__19869\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__19879\,
            I => \tok.S_5\
        );

    \I__4075\ : Odrv12
    port map (
            O => \N__19876\,
            I => \tok.S_5\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__19869\,
            I => \tok.S_5\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__19862\,
            I => \N__19859\
        );

    \I__4072\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__4070\ : Sp12to4
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__4069\ : Span12Mux_s6_v
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__4068\ : Odrv12
    port map (
            O => \N__19847\,
            I => \tok.n5_adj_775\
        );

    \I__4067\ : InMux
    port map (
            O => \N__19844\,
            I => \tok.n3929\
        );

    \I__4066\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__4064\ : Span12Mux_s6_v
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__4063\ : Odrv12
    port map (
            O => \N__19832\,
            I => \tok.n5_adj_773\
        );

    \I__4062\ : InMux
    port map (
            O => \N__19829\,
            I => \tok.n3930\
        );

    \I__4061\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19821\
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__19825\,
            I => \N__19818\
        );

    \I__4059\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19814\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__19821\,
            I => \N__19808\
        );

    \I__4057\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19803\
        );

    \I__4056\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19800\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__19814\,
            I => \N__19797\
        );

    \I__4054\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19794\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__19812\,
            I => \N__19791\
        );

    \I__4052\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19787\
        );

    \I__4051\ : Span4Mux_h
    port map (
            O => \N__19808\,
            I => \N__19784\
        );

    \I__4050\ : InMux
    port map (
            O => \N__19807\,
            I => \N__19779\
        );

    \I__4049\ : InMux
    port map (
            O => \N__19806\,
            I => \N__19779\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__19803\,
            I => \N__19776\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__19800\,
            I => \N__19771\
        );

    \I__4046\ : Span4Mux_s3_h
    port map (
            O => \N__19797\,
            I => \N__19766\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__19794\,
            I => \N__19766\
        );

    \I__4044\ : InMux
    port map (
            O => \N__19791\,
            I => \N__19763\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__19790\,
            I => \N__19758\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__19787\,
            I => \N__19754\
        );

    \I__4041\ : Span4Mux_s2_v
    port map (
            O => \N__19784\,
            I => \N__19749\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__19779\,
            I => \N__19749\
        );

    \I__4039\ : Span4Mux_h
    port map (
            O => \N__19776\,
            I => \N__19746\
        );

    \I__4038\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19743\
        );

    \I__4037\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19740\
        );

    \I__4036\ : Span4Mux_s3_v
    port map (
            O => \N__19771\,
            I => \N__19737\
        );

    \I__4035\ : Span4Mux_h
    port map (
            O => \N__19766\,
            I => \N__19732\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__19763\,
            I => \N__19732\
        );

    \I__4033\ : InMux
    port map (
            O => \N__19762\,
            I => \N__19729\
        );

    \I__4032\ : InMux
    port map (
            O => \N__19761\,
            I => \N__19722\
        );

    \I__4031\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19722\
        );

    \I__4030\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19722\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__19754\,
            I => \N__19717\
        );

    \I__4028\ : Span4Mux_v
    port map (
            O => \N__19749\,
            I => \N__19717\
        );

    \I__4027\ : Span4Mux_h
    port map (
            O => \N__19746\,
            I => \N__19714\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__19743\,
            I => \N__19709\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__19740\,
            I => \N__19709\
        );

    \I__4024\ : Span4Mux_h
    port map (
            O => \N__19737\,
            I => \N__19704\
        );

    \I__4023\ : Span4Mux_h
    port map (
            O => \N__19732\,
            I => \N__19704\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__19729\,
            I => \tok.A_low_7\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__19722\,
            I => \tok.A_low_7\
        );

    \I__4020\ : Odrv4
    port map (
            O => \N__19717\,
            I => \tok.A_low_7\
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__19714\,
            I => \tok.A_low_7\
        );

    \I__4018\ : Odrv12
    port map (
            O => \N__19709\,
            I => \tok.A_low_7\
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__19704\,
            I => \tok.A_low_7\
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__19691\,
            I => \N__19686\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__19690\,
            I => \N__19683\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__19689\,
            I => \N__19680\
        );

    \I__4013\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19675\
        );

    \I__4012\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19670\
        );

    \I__4011\ : InMux
    port map (
            O => \N__19680\,
            I => \N__19667\
        );

    \I__4010\ : InMux
    port map (
            O => \N__19679\,
            I => \N__19664\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__19678\,
            I => \N__19661\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__19675\,
            I => \N__19657\
        );

    \I__4007\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19652\
        );

    \I__4006\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19652\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__19670\,
            I => \N__19649\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19643\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__19664\,
            I => \N__19643\
        );

    \I__4002\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19640\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__19660\,
            I => \N__19637\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__19657\,
            I => \N__19631\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__19652\,
            I => \N__19631\
        );

    \I__3998\ : Span4Mux_v
    port map (
            O => \N__19649\,
            I => \N__19628\
        );

    \I__3997\ : InMux
    port map (
            O => \N__19648\,
            I => \N__19625\
        );

    \I__3996\ : Span4Mux_v
    port map (
            O => \N__19643\,
            I => \N__19622\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__19640\,
            I => \N__19619\
        );

    \I__3994\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19616\
        );

    \I__3993\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19613\
        );

    \I__3992\ : Span4Mux_h
    port map (
            O => \N__19631\,
            I => \N__19610\
        );

    \I__3991\ : Sp12to4
    port map (
            O => \N__19628\,
            I => \N__19599\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__19625\,
            I => \N__19599\
        );

    \I__3989\ : Sp12to4
    port map (
            O => \N__19622\,
            I => \N__19599\
        );

    \I__3988\ : Span12Mux_s7_v
    port map (
            O => \N__19619\,
            I => \N__19599\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__19616\,
            I => \N__19599\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__19613\,
            I => \tok.S_7\
        );

    \I__3985\ : Odrv4
    port map (
            O => \N__19610\,
            I => \tok.S_7\
        );

    \I__3984\ : Odrv12
    port map (
            O => \N__19599\,
            I => \tok.S_7\
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__19592\,
            I => \N__19589\
        );

    \I__3982\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__19586\,
            I => \N__19583\
        );

    \I__3980\ : Span4Mux_v
    port map (
            O => \N__19583\,
            I => \N__19580\
        );

    \I__3979\ : Span4Mux_h
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__19577\,
            I => \tok.n5_adj_752\
        );

    \I__3977\ : InMux
    port map (
            O => \N__19574\,
            I => \tok.n3931\
        );

    \I__3976\ : CascadeMux
    port map (
            O => \N__19571\,
            I => \N__19567\
        );

    \I__3975\ : InMux
    port map (
            O => \N__19570\,
            I => \N__19564\
        );

    \I__3974\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19559\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__19564\,
            I => \N__19556\
        );

    \I__3972\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19550\
        );

    \I__3971\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19546\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__19559\,
            I => \N__19541\
        );

    \I__3969\ : Span4Mux_v
    port map (
            O => \N__19556\,
            I => \N__19541\
        );

    \I__3968\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19538\
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__19554\,
            I => \N__19535\
        );

    \I__3966\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19532\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__19550\,
            I => \N__19529\
        );

    \I__3964\ : InMux
    port map (
            O => \N__19549\,
            I => \N__19526\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__19546\,
            I => \N__19523\
        );

    \I__3962\ : Span4Mux_v
    port map (
            O => \N__19541\,
            I => \N__19518\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__19538\,
            I => \N__19518\
        );

    \I__3960\ : InMux
    port map (
            O => \N__19535\,
            I => \N__19515\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__19532\,
            I => \N__19512\
        );

    \I__3958\ : Span4Mux_v
    port map (
            O => \N__19529\,
            I => \N__19507\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__19526\,
            I => \N__19507\
        );

    \I__3956\ : Span4Mux_v
    port map (
            O => \N__19523\,
            I => \N__19504\
        );

    \I__3955\ : Span4Mux_h
    port map (
            O => \N__19518\,
            I => \N__19501\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__19515\,
            I => \N__19492\
        );

    \I__3953\ : Span4Mux_v
    port map (
            O => \N__19512\,
            I => \N__19492\
        );

    \I__3952\ : Span4Mux_v
    port map (
            O => \N__19507\,
            I => \N__19492\
        );

    \I__3951\ : Span4Mux_h
    port map (
            O => \N__19504\,
            I => \N__19492\
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__19501\,
            I => \tok.S_8\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__19492\,
            I => \tok.S_8\
        );

    \I__3948\ : InMux
    port map (
            O => \N__19487\,
            I => \bfn_9_9_0_\
        );

    \I__3947\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__19481\,
            I => \N__19477\
        );

    \I__3945\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19474\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__19477\,
            I => n10_adj_875
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__19474\,
            I => n10_adj_875
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__19469\,
            I => \N__19465\
        );

    \I__3941\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19462\
        );

    \I__3940\ : InMux
    port map (
            O => \N__19465\,
            I => \N__19458\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__19462\,
            I => \N__19455\
        );

    \I__3938\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19451\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__19458\,
            I => \N__19448\
        );

    \I__3936\ : Span4Mux_v
    port map (
            O => \N__19455\,
            I => \N__19445\
        );

    \I__3935\ : InMux
    port map (
            O => \N__19454\,
            I => \N__19442\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__19451\,
            I => \c_stk_w_7_N_18_0\
        );

    \I__3933\ : Odrv12
    port map (
            O => \N__19448\,
            I => \c_stk_w_7_N_18_0\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__19445\,
            I => \c_stk_w_7_N_18_0\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__19442\,
            I => \c_stk_w_7_N_18_0\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__19433\,
            I => \N__19427\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__19432\,
            I => \N__19424\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__19431\,
            I => \N__19421\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__19430\,
            I => \N__19418\
        );

    \I__3926\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19409\
        );

    \I__3925\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19409\
        );

    \I__3924\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19409\
        );

    \I__3923\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19409\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19402\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__19408\,
            I => \N__19399\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__19407\,
            I => \N__19396\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__19406\,
            I => \N__19393\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__19405\,
            I => \N__19390\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__19402\,
            I => \N__19387\
        );

    \I__3916\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19378\
        );

    \I__3915\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19378\
        );

    \I__3914\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19378\
        );

    \I__3913\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19378\
        );

    \I__3912\ : Span4Mux_s0_v
    port map (
            O => \N__19387\,
            I => \N__19372\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__19378\,
            I => \N__19372\
        );

    \I__3910\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19368\
        );

    \I__3909\ : Span4Mux_v
    port map (
            O => \N__19372\,
            I => \N__19365\
        );

    \I__3908\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19362\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__19368\,
            I => \N__19359\
        );

    \I__3906\ : Span4Mux_h
    port map (
            O => \N__19365\,
            I => \N__19356\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__19362\,
            I => \tok.found_slot\
        );

    \I__3904\ : Odrv12
    port map (
            O => \N__19359\,
            I => \tok.found_slot\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__19356\,
            I => \tok.found_slot\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__19349\,
            I => \tok.n5_adj_655_cascade_\
        );

    \I__3901\ : InMux
    port map (
            O => \N__19346\,
            I => \N__19340\
        );

    \I__3900\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19333\
        );

    \I__3899\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19333\
        );

    \I__3898\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19333\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__19340\,
            I => \N__19330\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__19333\,
            I => \N__19327\
        );

    \I__3895\ : Span4Mux_h
    port map (
            O => \N__19330\,
            I => \N__19324\
        );

    \I__3894\ : Span4Mux_h
    port map (
            O => \N__19327\,
            I => \N__19321\
        );

    \I__3893\ : Span4Mux_h
    port map (
            O => \N__19324\,
            I => \N__19318\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__19321\,
            I => \tok.uart_tx_busy\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__19318\,
            I => \tok.uart_tx_busy\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__19313\,
            I => \N__19309\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__19312\,
            I => \N__19306\
        );

    \I__3888\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19303\
        );

    \I__3887\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19300\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__19303\,
            I => \N__19294\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__19300\,
            I => \N__19294\
        );

    \I__3884\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19291\
        );

    \I__3883\ : Span4Mux_h
    port map (
            O => \N__19294\,
            I => \N__19288\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__19291\,
            I => \tok.uart_rx_valid\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__19288\,
            I => \tok.uart_rx_valid\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__19283\,
            I => \tok.uart_stall_cascade_\
        );

    \I__3879\ : InMux
    port map (
            O => \N__19280\,
            I => \N__19270\
        );

    \I__3878\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19270\
        );

    \I__3877\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19261\
        );

    \I__3876\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19261\
        );

    \I__3875\ : InMux
    port map (
            O => \N__19276\,
            I => \N__19261\
        );

    \I__3874\ : InMux
    port map (
            O => \N__19275\,
            I => \N__19261\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__19270\,
            I => \N__19257\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__19261\,
            I => \N__19254\
        );

    \I__3871\ : InMux
    port map (
            O => \N__19260\,
            I => \N__19251\
        );

    \I__3870\ : Span4Mux_h
    port map (
            O => \N__19257\,
            I => \N__19248\
        );

    \I__3869\ : Span4Mux_s3_v
    port map (
            O => \N__19254\,
            I => \N__19243\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__19251\,
            I => \N__19243\
        );

    \I__3867\ : Sp12to4
    port map (
            O => \N__19248\,
            I => \N__19240\
        );

    \I__3866\ : Span4Mux_v
    port map (
            O => \N__19243\,
            I => \N__19237\
        );

    \I__3865\ : Odrv12
    port map (
            O => \N__19240\,
            I => \tok.n2732\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__19237\,
            I => \tok.n2732\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__19232\,
            I => \tok.n2732_cascade_\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__19229\,
            I => \N__19225\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__19228\,
            I => \N__19222\
        );

    \I__3860\ : CascadeBuf
    port map (
            O => \N__19225\,
            I => \N__19219\
        );

    \I__3859\ : CascadeBuf
    port map (
            O => \N__19222\,
            I => \N__19216\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__19219\,
            I => \N__19211\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__19216\,
            I => \N__19208\
        );

    \I__3856\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19205\
        );

    \I__3855\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19202\
        );

    \I__3854\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19199\
        );

    \I__3853\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19196\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__19205\,
            I => \N__19191\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19191\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__19199\,
            I => \N__19188\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__19196\,
            I => \N__19185\
        );

    \I__3848\ : Span4Mux_h
    port map (
            O => \N__19191\,
            I => \N__19181\
        );

    \I__3847\ : Span4Mux_h
    port map (
            O => \N__19188\,
            I => \N__19178\
        );

    \I__3846\ : Span4Mux_h
    port map (
            O => \N__19185\,
            I => \N__19175\
        );

    \I__3845\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19172\
        );

    \I__3844\ : Span4Mux_v
    port map (
            O => \N__19181\,
            I => \N__19167\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__19178\,
            I => \N__19167\
        );

    \I__3842\ : Span4Mux_h
    port map (
            O => \N__19175\,
            I => \N__19164\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__19172\,
            I => \tok.n43\
        );

    \I__3840\ : Odrv4
    port map (
            O => \N__19167\,
            I => \tok.n43\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__19164\,
            I => \tok.n43\
        );

    \I__3838\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__19154\,
            I => \tok.n5_adj_655\
        );

    \I__3836\ : SRMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__19148\,
            I => \N__19145\
        );

    \I__3834\ : Span4Mux_h
    port map (
            O => \N__19145\,
            I => \N__19139\
        );

    \I__3833\ : SRMux
    port map (
            O => \N__19144\,
            I => \N__19136\
        );

    \I__3832\ : SRMux
    port map (
            O => \N__19143\,
            I => \N__19132\
        );

    \I__3831\ : SRMux
    port map (
            O => \N__19142\,
            I => \N__19127\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__19139\,
            I => \N__19122\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__19136\,
            I => \N__19122\
        );

    \I__3828\ : SRMux
    port map (
            O => \N__19135\,
            I => \N__19119\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__19132\,
            I => \N__19115\
        );

    \I__3826\ : SRMux
    port map (
            O => \N__19131\,
            I => \N__19111\
        );

    \I__3825\ : SRMux
    port map (
            O => \N__19130\,
            I => \N__19108\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__19127\,
            I => \N__19105\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__19122\,
            I => \N__19100\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__19119\,
            I => \N__19100\
        );

    \I__3821\ : SRMux
    port map (
            O => \N__19118\,
            I => \N__19097\
        );

    \I__3820\ : Span4Mux_h
    port map (
            O => \N__19115\,
            I => \N__19093\
        );

    \I__3819\ : SRMux
    port map (
            O => \N__19114\,
            I => \N__19090\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__19111\,
            I => \N__19087\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19083\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__19105\,
            I => \N__19076\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__19100\,
            I => \N__19076\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__19097\,
            I => \N__19076\
        );

    \I__3813\ : SRMux
    port map (
            O => \N__19096\,
            I => \N__19073\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__19093\,
            I => \N__19070\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__19090\,
            I => \N__19067\
        );

    \I__3810\ : Span4Mux_v
    port map (
            O => \N__19087\,
            I => \N__19063\
        );

    \I__3809\ : SRMux
    port map (
            O => \N__19086\,
            I => \N__19060\
        );

    \I__3808\ : Span4Mux_h
    port map (
            O => \N__19083\,
            I => \N__19053\
        );

    \I__3807\ : Span4Mux_h
    port map (
            O => \N__19076\,
            I => \N__19053\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__19073\,
            I => \N__19053\
        );

    \I__3805\ : IoSpan4Mux
    port map (
            O => \N__19070\,
            I => \N__19050\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__19067\,
            I => \N__19047\
        );

    \I__3803\ : SRMux
    port map (
            O => \N__19066\,
            I => \N__19044\
        );

    \I__3802\ : Span4Mux_v
    port map (
            O => \N__19063\,
            I => \N__19039\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__19060\,
            I => \N__19039\
        );

    \I__3800\ : Span4Mux_v
    port map (
            O => \N__19053\,
            I => \N__19036\
        );

    \I__3799\ : IoSpan4Mux
    port map (
            O => \N__19050\,
            I => \N__19033\
        );

    \I__3798\ : Span4Mux_h
    port map (
            O => \N__19047\,
            I => \N__19030\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__19044\,
            I => \N__19027\
        );

    \I__3796\ : Span4Mux_v
    port map (
            O => \N__19039\,
            I => \N__19022\
        );

    \I__3795\ : Span4Mux_h
    port map (
            O => \N__19036\,
            I => \N__19022\
        );

    \I__3794\ : Span4Mux_s0_v
    port map (
            O => \N__19033\,
            I => \N__19017\
        );

    \I__3793\ : Span4Mux_v
    port map (
            O => \N__19030\,
            I => \N__19017\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__19027\,
            I => \N__19012\
        );

    \I__3791\ : Span4Mux_s0_v
    port map (
            O => \N__19022\,
            I => \N__19012\
        );

    \I__3790\ : Odrv4
    port map (
            O => \N__19017\,
            I => \tok.reset_N_2\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__19012\,
            I => \tok.reset_N_2\
        );

    \I__3788\ : InMux
    port map (
            O => \N__19007\,
            I => \N__18998\
        );

    \I__3787\ : InMux
    port map (
            O => \N__19006\,
            I => \N__18998\
        );

    \I__3786\ : InMux
    port map (
            O => \N__19005\,
            I => \N__18998\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__18998\,
            I => \tok.uart_stall\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__3783\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18980\
        );

    \I__3782\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18980\
        );

    \I__3781\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18980\
        );

    \I__3780\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18980\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__18980\,
            I => \N__18977\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__18977\,
            I => \tok.n2724\
        );

    \I__3777\ : InMux
    port map (
            O => \N__18974\,
            I => \N__18964\
        );

    \I__3776\ : InMux
    port map (
            O => \N__18973\,
            I => \N__18964\
        );

    \I__3775\ : InMux
    port map (
            O => \N__18972\,
            I => \N__18955\
        );

    \I__3774\ : InMux
    port map (
            O => \N__18971\,
            I => \N__18955\
        );

    \I__3773\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18955\
        );

    \I__3772\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18955\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__18964\,
            I => \N__18949\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__18955\,
            I => \N__18949\
        );

    \I__3769\ : InMux
    port map (
            O => \N__18954\,
            I => \N__18946\
        );

    \I__3768\ : Span4Mux_s3_v
    port map (
            O => \N__18949\,
            I => \N__18941\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__18946\,
            I => \N__18941\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__18941\,
            I => \N__18937\
        );

    \I__3765\ : InMux
    port map (
            O => \N__18940\,
            I => \N__18934\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__18937\,
            I => \tok.n4431\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__18934\,
            I => \tok.n4431\
        );

    \I__3762\ : InMux
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__18926\,
            I => \N__18923\
        );

    \I__3760\ : Span4Mux_h
    port map (
            O => \N__18923\,
            I => \N__18920\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__18920\,
            I => \tok.n5_adj_682\
        );

    \I__3758\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18908\
        );

    \I__3756\ : InMux
    port map (
            O => \N__18913\,
            I => \N__18901\
        );

    \I__3755\ : InMux
    port map (
            O => \N__18912\,
            I => \N__18901\
        );

    \I__3754\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18901\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__18908\,
            I => \tok.tc_plus_1_6\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__18901\,
            I => \tok.tc_plus_1_6\
        );

    \I__3751\ : InMux
    port map (
            O => \N__18896\,
            I => \tok.n3900\
        );

    \I__3750\ : InMux
    port map (
            O => \N__18893\,
            I => \tok.n3901\
        );

    \I__3749\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__3747\ : Span4Mux_v
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__18881\,
            I => \N__18875\
        );

    \I__3745\ : InMux
    port map (
            O => \N__18880\,
            I => \N__18872\
        );

    \I__3744\ : InMux
    port map (
            O => \N__18879\,
            I => \N__18867\
        );

    \I__3743\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18867\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__18875\,
            I => \tok.tc_plus_1_7\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__18872\,
            I => \tok.tc_plus_1_7\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__18867\,
            I => \tok.tc_plus_1_7\
        );

    \I__3739\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__18857\,
            I => \N__18853\
        );

    \I__3737\ : InMux
    port map (
            O => \N__18856\,
            I => \N__18850\
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__18853\,
            I => n92_adj_872
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__18850\,
            I => n92_adj_872
        );

    \I__3734\ : CascadeMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__3733\ : InMux
    port map (
            O => \N__18842\,
            I => \N__18837\
        );

    \I__3732\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18833\
        );

    \I__3731\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18830\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__18837\,
            I => \N__18827\
        );

    \I__3729\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18824\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__18833\,
            I => \c_stk_w_7_N_18_7\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__18830\,
            I => \c_stk_w_7_N_18_7\
        );

    \I__3726\ : Odrv4
    port map (
            O => \N__18827\,
            I => \c_stk_w_7_N_18_7\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__18824\,
            I => \c_stk_w_7_N_18_7\
        );

    \I__3724\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18811\
        );

    \I__3723\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18808\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__18811\,
            I => n92_adj_871
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__18808\,
            I => n92_adj_871
        );

    \I__3720\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18798\
        );

    \I__3719\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18795\
        );

    \I__3718\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18791\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__18798\,
            I => \N__18788\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__18795\,
            I => \N__18785\
        );

    \I__3715\ : InMux
    port map (
            O => \N__18794\,
            I => \N__18782\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__18791\,
            I => \c_stk_w_7_N_18_6\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__18788\,
            I => \c_stk_w_7_N_18_6\
        );

    \I__3712\ : Odrv4
    port map (
            O => \N__18785\,
            I => \c_stk_w_7_N_18_6\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__18782\,
            I => \c_stk_w_7_N_18_6\
        );

    \I__3710\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__18770\,
            I => n92
        );

    \I__3708\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18761\
        );

    \I__3707\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18756\
        );

    \I__3706\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18756\
        );

    \I__3705\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18753\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__18761\,
            I => \c_stk_w_7_N_18_1\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__18756\,
            I => \c_stk_w_7_N_18_1\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__18753\,
            I => \c_stk_w_7_N_18_1\
        );

    \I__3701\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18740\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__18745\,
            I => \N__18736\
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__18744\,
            I => \N__18733\
        );

    \I__3698\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18730\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__18740\,
            I => \N__18727\
        );

    \I__3696\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18722\
        );

    \I__3695\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18722\
        );

    \I__3694\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18719\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__18730\,
            I => \tok.c_stk_r_7\
        );

    \I__3692\ : Odrv4
    port map (
            O => \N__18727\,
            I => \tok.c_stk_r_7\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__18722\,
            I => \tok.c_stk_r_7\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__18719\,
            I => \tok.c_stk_r_7\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__18710\,
            I => \tok.ram.n4696_cascade_\
        );

    \I__3688\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__18704\,
            I => \tok.n4602\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__18701\,
            I => \tok.n1_adj_798_cascade_\
        );

    \I__3685\ : InMux
    port map (
            O => \N__18698\,
            I => \N__18695\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__18695\,
            I => \tok.n13_adj_799\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__3682\ : InMux
    port map (
            O => \N__18689\,
            I => \N__18686\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__3680\ : Span4Mux_h
    port map (
            O => \N__18683\,
            I => \N__18680\
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__18680\,
            I => \tok.tc_0\
        );

    \I__3678\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__18674\,
            I => \N__18668\
        );

    \I__3676\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18661\
        );

    \I__3675\ : InMux
    port map (
            O => \N__18672\,
            I => \N__18661\
        );

    \I__3674\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18661\
        );

    \I__3673\ : Span4Mux_v
    port map (
            O => \N__18668\,
            I => \N__18656\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__18661\,
            I => \N__18656\
        );

    \I__3671\ : Odrv4
    port map (
            O => \N__18656\,
            I => \tok.tc_plus_1_0\
        );

    \I__3670\ : InMux
    port map (
            O => \N__18653\,
            I => \bfn_9_5_0_\
        );

    \I__3669\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__18647\,
            I => \N__18644\
        );

    \I__3667\ : Span12Mux_s9_v
    port map (
            O => \N__18644\,
            I => \N__18638\
        );

    \I__3666\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18631\
        );

    \I__3665\ : InMux
    port map (
            O => \N__18642\,
            I => \N__18631\
        );

    \I__3664\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18631\
        );

    \I__3663\ : Odrv12
    port map (
            O => \N__18638\,
            I => \tok.tc_plus_1_1\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__18631\,
            I => \tok.tc_plus_1_1\
        );

    \I__3661\ : InMux
    port map (
            O => \N__18626\,
            I => \tok.n3895\
        );

    \I__3660\ : InMux
    port map (
            O => \N__18623\,
            I => \tok.n3896\
        );

    \I__3659\ : InMux
    port map (
            O => \N__18620\,
            I => \tok.n3897\
        );

    \I__3658\ : InMux
    port map (
            O => \N__18617\,
            I => \tok.n3898\
        );

    \I__3657\ : InMux
    port map (
            O => \N__18614\,
            I => \tok.n3899\
        );

    \I__3656\ : CascadeMux
    port map (
            O => \N__18611\,
            I => \tok.n13_adj_713_cascade_\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__18608\,
            I => \tok.C_stk.n4894_cascade_\
        );

    \I__3654\ : CascadeMux
    port map (
            O => \N__18605\,
            I => \N__18599\
        );

    \I__3653\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18595\
        );

    \I__3652\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18592\
        );

    \I__3651\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18587\
        );

    \I__3650\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18587\
        );

    \I__3649\ : InMux
    port map (
            O => \N__18598\,
            I => \N__18584\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__18595\,
            I => \tok.c_stk_r_0\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__18592\,
            I => \tok.c_stk_r_0\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__18587\,
            I => \tok.c_stk_r_0\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__18584\,
            I => \tok.c_stk_r_0\
        );

    \I__3644\ : CascadeMux
    port map (
            O => \N__18575\,
            I => \tok.ram.n4717_cascade_\
        );

    \I__3643\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__18569\,
            I => \tok.n1_adj_712\
        );

    \I__3641\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__18563\,
            I => \N__18559\
        );

    \I__3639\ : InMux
    port map (
            O => \N__18562\,
            I => \N__18556\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__18559\,
            I => \tok.C_stk.tail_7\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__18556\,
            I => \tok.C_stk.tail_7\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__18551\,
            I => \tok.C_stk.n4912_cascade_\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__3634\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__18539\,
            I => \tok.tc_6\
        );

    \I__3631\ : InMux
    port map (
            O => \N__18536\,
            I => \N__18532\
        );

    \I__3630\ : InMux
    port map (
            O => \N__18535\,
            I => \N__18529\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__18532\,
            I => \tok.tail_26\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__18529\,
            I => \tok.tail_26\
        );

    \I__3627\ : InMux
    port map (
            O => \N__18524\,
            I => \N__18520\
        );

    \I__3626\ : InMux
    port map (
            O => \N__18523\,
            I => \N__18517\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__18520\,
            I => \tok.tail_12\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__18517\,
            I => \tok.tail_12\
        );

    \I__3623\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18508\
        );

    \I__3622\ : InMux
    port map (
            O => \N__18511\,
            I => \N__18505\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__18508\,
            I => \tok.C_stk.tail_36\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__18505\,
            I => \tok.C_stk.tail_36\
        );

    \I__3619\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__3617\ : Span4Mux_s2_v
    port map (
            O => \N__18494\,
            I => \N__18490\
        );

    \I__3616\ : InMux
    port map (
            O => \N__18493\,
            I => \N__18487\
        );

    \I__3615\ : Odrv4
    port map (
            O => \N__18490\,
            I => \tok.tail_56\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__18487\,
            I => \tok.tail_56\
        );

    \I__3613\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18478\
        );

    \I__3612\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18475\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__18478\,
            I => \tok.tail_40\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__18475\,
            I => \tok.tail_40\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__3608\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__3606\ : Span4Mux_v
    port map (
            O => \N__18461\,
            I => \N__18457\
        );

    \I__3605\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18454\
        );

    \I__3604\ : Odrv4
    port map (
            O => \N__18457\,
            I => \tok.tail_48\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__18454\,
            I => \tok.tail_48\
        );

    \I__3602\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__18443\,
            I => \tok.n83_adj_704\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__18440\,
            I => \tok.n4694_cascade_\
        );

    \I__3598\ : CascadeMux
    port map (
            O => \N__18437\,
            I => \N__18433\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__18436\,
            I => \N__18430\
        );

    \I__3596\ : CascadeBuf
    port map (
            O => \N__18433\,
            I => \N__18427\
        );

    \I__3595\ : CascadeBuf
    port map (
            O => \N__18430\,
            I => \N__18424\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__18427\,
            I => \N__18421\
        );

    \I__3593\ : CascadeMux
    port map (
            O => \N__18424\,
            I => \N__18418\
        );

    \I__3592\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18415\
        );

    \I__3591\ : InMux
    port map (
            O => \N__18418\,
            I => \N__18412\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__18415\,
            I => \N__18409\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__18412\,
            I => \N__18403\
        );

    \I__3588\ : Span4Mux_h
    port map (
            O => \N__18409\,
            I => \N__18400\
        );

    \I__3587\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18397\
        );

    \I__3586\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18394\
        );

    \I__3585\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18391\
        );

    \I__3584\ : Span4Mux_v
    port map (
            O => \N__18403\,
            I => \N__18388\
        );

    \I__3583\ : Span4Mux_h
    port map (
            O => \N__18400\,
            I => \N__18385\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__18397\,
            I => \tok.n50\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__18394\,
            I => \tok.n50\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__18391\,
            I => \tok.n50\
        );

    \I__3579\ : Odrv4
    port map (
            O => \N__18388\,
            I => \tok.n50\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__18385\,
            I => \tok.n50\
        );

    \I__3577\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__18371\,
            I => \tok.n33_adj_841\
        );

    \I__3575\ : InMux
    port map (
            O => \N__18368\,
            I => \tok.n3888\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__18365\,
            I => \N__18361\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__18364\,
            I => \N__18358\
        );

    \I__3572\ : CascadeBuf
    port map (
            O => \N__18361\,
            I => \N__18355\
        );

    \I__3571\ : CascadeBuf
    port map (
            O => \N__18358\,
            I => \N__18352\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__18355\,
            I => \N__18349\
        );

    \I__3569\ : CascadeMux
    port map (
            O => \N__18352\,
            I => \N__18346\
        );

    \I__3568\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18343\
        );

    \I__3567\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18340\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__18343\,
            I => \N__18335\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__18340\,
            I => \N__18335\
        );

    \I__3564\ : Span4Mux_v
    port map (
            O => \N__18335\,
            I => \N__18329\
        );

    \I__3563\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18326\
        );

    \I__3562\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18323\
        );

    \I__3561\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18320\
        );

    \I__3560\ : Span4Mux_h
    port map (
            O => \N__18329\,
            I => \N__18317\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__18326\,
            I => \tok.n49\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__18323\,
            I => \tok.n49\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__18320\,
            I => \tok.n49\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__18317\,
            I => \tok.n49\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__3554\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__18302\,
            I => \tok.n33_adj_665\
        );

    \I__3552\ : InMux
    port map (
            O => \N__18299\,
            I => \tok.n3889\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__18296\,
            I => \N__18292\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__18295\,
            I => \N__18289\
        );

    \I__3549\ : CascadeBuf
    port map (
            O => \N__18292\,
            I => \N__18286\
        );

    \I__3548\ : CascadeBuf
    port map (
            O => \N__18289\,
            I => \N__18283\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__18286\,
            I => \N__18280\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__18283\,
            I => \N__18277\
        );

    \I__3545\ : InMux
    port map (
            O => \N__18280\,
            I => \N__18274\
        );

    \I__3544\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18270\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__18274\,
            I => \N__18267\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__18273\,
            I => \N__18264\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__18270\,
            I => \N__18257\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__18267\,
            I => \N__18257\
        );

    \I__3539\ : InMux
    port map (
            O => \N__18264\,
            I => \N__18254\
        );

    \I__3538\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18251\
        );

    \I__3537\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18248\
        );

    \I__3536\ : Span4Mux_h
    port map (
            O => \N__18257\,
            I => \N__18245\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__18254\,
            I => \tok.n47\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__18251\,
            I => \tok.n47\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__18248\,
            I => \tok.n47\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__18245\,
            I => \tok.n47\
        );

    \I__3531\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__3529\ : Span4Mux_v
    port map (
            O => \N__18230\,
            I => \N__18227\
        );

    \I__3528\ : Odrv4
    port map (
            O => \N__18227\,
            I => \tok.n33_adj_755\
        );

    \I__3527\ : InMux
    port map (
            O => \N__18224\,
            I => \tok.n3890\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__18221\,
            I => \N__18217\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__18220\,
            I => \N__18214\
        );

    \I__3524\ : CascadeBuf
    port map (
            O => \N__18217\,
            I => \N__18209\
        );

    \I__3523\ : CascadeBuf
    port map (
            O => \N__18214\,
            I => \N__18206\
        );

    \I__3522\ : InMux
    port map (
            O => \N__18213\,
            I => \N__18203\
        );

    \I__3521\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18200\
        );

    \I__3520\ : CascadeMux
    port map (
            O => \N__18209\,
            I => \N__18197\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__18206\,
            I => \N__18194\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__18203\,
            I => \N__18189\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__18200\,
            I => \N__18189\
        );

    \I__3516\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18186\
        );

    \I__3515\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18183\
        );

    \I__3514\ : Span4Mux_s2_v
    port map (
            O => \N__18189\,
            I => \N__18180\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__18186\,
            I => \N__18175\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__18183\,
            I => \N__18175\
        );

    \I__3511\ : Span4Mux_v
    port map (
            O => \N__18180\,
            I => \N__18171\
        );

    \I__3510\ : Sp12to4
    port map (
            O => \N__18175\,
            I => \N__18168\
        );

    \I__3509\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18165\
        );

    \I__3508\ : Sp12to4
    port map (
            O => \N__18171\,
            I => \N__18160\
        );

    \I__3507\ : Span12Mux_s6_v
    port map (
            O => \N__18168\,
            I => \N__18160\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__18165\,
            I => \tok.n45\
        );

    \I__3505\ : Odrv12
    port map (
            O => \N__18160\,
            I => \tok.n45\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__3503\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__18149\,
            I => \N__18146\
        );

    \I__3501\ : Span4Mux_v
    port map (
            O => \N__18146\,
            I => \N__18143\
        );

    \I__3500\ : Odrv4
    port map (
            O => \N__18143\,
            I => \tok.n33_adj_852\
        );

    \I__3499\ : InMux
    port map (
            O => \N__18140\,
            I => \tok.n3891\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__18137\,
            I => \N__18133\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__18136\,
            I => \N__18130\
        );

    \I__3496\ : CascadeBuf
    port map (
            O => \N__18133\,
            I => \N__18127\
        );

    \I__3495\ : CascadeBuf
    port map (
            O => \N__18130\,
            I => \N__18124\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__18127\,
            I => \N__18121\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__18124\,
            I => \N__18118\
        );

    \I__3492\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18115\
        );

    \I__3491\ : InMux
    port map (
            O => \N__18118\,
            I => \N__18109\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__18115\,
            I => \N__18106\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__18114\,
            I => \N__18103\
        );

    \I__3488\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18100\
        );

    \I__3487\ : InMux
    port map (
            O => \N__18112\,
            I => \N__18097\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__18109\,
            I => \N__18092\
        );

    \I__3485\ : Span4Mux_h
    port map (
            O => \N__18106\,
            I => \N__18092\
        );

    \I__3484\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18089\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__18100\,
            I => \N__18084\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__18097\,
            I => \N__18084\
        );

    \I__3481\ : Span4Mux_v
    port map (
            O => \N__18092\,
            I => \N__18081\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__18089\,
            I => \tok.n44\
        );

    \I__3479\ : Odrv12
    port map (
            O => \N__18084\,
            I => \tok.n44\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__18081\,
            I => \tok.n44\
        );

    \I__3477\ : InMux
    port map (
            O => \N__18074\,
            I => \tok.n3892\
        );

    \I__3476\ : InMux
    port map (
            O => \N__18071\,
            I => \tok.n3893\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__18068\,
            I => \N__18064\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__18067\,
            I => \N__18061\
        );

    \I__3473\ : CascadeBuf
    port map (
            O => \N__18064\,
            I => \N__18058\
        );

    \I__3472\ : CascadeBuf
    port map (
            O => \N__18061\,
            I => \N__18055\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__18058\,
            I => \N__18052\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__18055\,
            I => \N__18049\
        );

    \I__3469\ : InMux
    port map (
            O => \N__18052\,
            I => \N__18046\
        );

    \I__3468\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18041\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__18046\,
            I => \N__18038\
        );

    \I__3466\ : InMux
    port map (
            O => \N__18045\,
            I => \N__18034\
        );

    \I__3465\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18031\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__18041\,
            I => \N__18028\
        );

    \I__3463\ : Span4Mux_h
    port map (
            O => \N__18038\,
            I => \N__18025\
        );

    \I__3462\ : InMux
    port map (
            O => \N__18037\,
            I => \N__18022\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__18034\,
            I => \N__18017\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__18031\,
            I => \N__18017\
        );

    \I__3459\ : Span4Mux_v
    port map (
            O => \N__18028\,
            I => \N__18014\
        );

    \I__3458\ : Span4Mux_v
    port map (
            O => \N__18025\,
            I => \N__18011\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__18022\,
            I => \tok.n39\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__18017\,
            I => \tok.n39\
        );

    \I__3455\ : Odrv4
    port map (
            O => \N__18014\,
            I => \tok.n39\
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__18011\,
            I => \tok.n39\
        );

    \I__3453\ : InMux
    port map (
            O => \N__18002\,
            I => \tok.n3894\
        );

    \I__3452\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__17996\,
            I => \N__17993\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__17993\,
            I => \tok.n33_adj_643\
        );

    \I__3449\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17986\
        );

    \I__3448\ : InMux
    port map (
            O => \N__17989\,
            I => \N__17983\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__17986\,
            I => \tok.C_stk.tail_20\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__17983\,
            I => \tok.C_stk.tail_20\
        );

    \I__3445\ : InMux
    port map (
            O => \N__17978\,
            I => \N__17975\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__17975\,
            I => \N__17972\
        );

    \I__3443\ : Span4Mux_v
    port map (
            O => \N__17972\,
            I => \N__17969\
        );

    \I__3442\ : Span4Mux_s2_v
    port map (
            O => \N__17969\,
            I => \N__17966\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__17966\,
            I => \tok.n9_adj_689\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__17963\,
            I => \tok.n181_cascade_\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__17960\,
            I => \tok.n12_cascade_\
        );

    \I__3438\ : InMux
    port map (
            O => \N__17957\,
            I => \N__17954\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__17954\,
            I => \N__17951\
        );

    \I__3436\ : Odrv12
    port map (
            O => \N__17951\,
            I => \tok.n6_adj_653\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__17948\,
            I => \tok.n20_cascade_\
        );

    \I__3434\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17942\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__17942\,
            I => \N__17939\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__17939\,
            I => \tok.n16\
        );

    \I__3431\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17933\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__17933\,
            I => \N__17930\
        );

    \I__3429\ : Span4Mux_h
    port map (
            O => \N__17930\,
            I => \N__17927\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__17927\,
            I => \tok.n4684\
        );

    \I__3427\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17916\
        );

    \I__3426\ : InMux
    port map (
            O => \N__17923\,
            I => \N__17916\
        );

    \I__3425\ : InMux
    port map (
            O => \N__17922\,
            I => \N__17913\
        );

    \I__3424\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17910\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__17916\,
            I => \N__17905\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__17913\,
            I => \N__17899\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__17910\,
            I => \N__17899\
        );

    \I__3420\ : InMux
    port map (
            O => \N__17909\,
            I => \N__17894\
        );

    \I__3419\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17894\
        );

    \I__3418\ : Span4Mux_h
    port map (
            O => \N__17905\,
            I => \N__17885\
        );

    \I__3417\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17882\
        );

    \I__3416\ : Span4Mux_h
    port map (
            O => \N__17899\,
            I => \N__17875\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__17894\,
            I => \N__17875\
        );

    \I__3414\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17870\
        );

    \I__3413\ : InMux
    port map (
            O => \N__17892\,
            I => \N__17870\
        );

    \I__3412\ : InMux
    port map (
            O => \N__17891\,
            I => \N__17865\
        );

    \I__3411\ : InMux
    port map (
            O => \N__17890\,
            I => \N__17865\
        );

    \I__3410\ : InMux
    port map (
            O => \N__17889\,
            I => \N__17862\
        );

    \I__3409\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17859\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__17885\,
            I => \N__17854\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__17882\,
            I => \N__17854\
        );

    \I__3406\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17849\
        );

    \I__3405\ : InMux
    port map (
            O => \N__17880\,
            I => \N__17849\
        );

    \I__3404\ : Odrv4
    port map (
            O => \N__17875\,
            I => \tok.n892\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__17870\,
            I => \tok.n892\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__17865\,
            I => \tok.n892\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__17862\,
            I => \tok.n892\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__17859\,
            I => \tok.n892\
        );

    \I__3399\ : Odrv4
    port map (
            O => \N__17854\,
            I => \tok.n892\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__17849\,
            I => \tok.n892\
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__17834\,
            I => \tok.n177_cascade_\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__17831\,
            I => \tok.n12_adj_696_cascade_\
        );

    \I__3395\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__17825\,
            I => \N__17822\
        );

    \I__3393\ : Odrv12
    port map (
            O => \N__17822\,
            I => \tok.n20_adj_700\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__17819\,
            I => \N__17815\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__17818\,
            I => \N__17812\
        );

    \I__3390\ : CascadeBuf
    port map (
            O => \N__17815\,
            I => \N__17809\
        );

    \I__3389\ : CascadeBuf
    port map (
            O => \N__17812\,
            I => \N__17806\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__17809\,
            I => \N__17803\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__17806\,
            I => \N__17800\
        );

    \I__3386\ : InMux
    port map (
            O => \N__17803\,
            I => \N__17797\
        );

    \I__3385\ : InMux
    port map (
            O => \N__17800\,
            I => \N__17793\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__17797\,
            I => \N__17790\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__17796\,
            I => \N__17787\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__17793\,
            I => \N__17780\
        );

    \I__3381\ : Span4Mux_h
    port map (
            O => \N__17790\,
            I => \N__17780\
        );

    \I__3380\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17777\
        );

    \I__3379\ : InMux
    port map (
            O => \N__17786\,
            I => \N__17774\
        );

    \I__3378\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17771\
        );

    \I__3377\ : Span4Mux_v
    port map (
            O => \N__17780\,
            I => \N__17768\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__17777\,
            I => \tok.n52\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__17774\,
            I => \tok.n52\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__17771\,
            I => \tok.n52\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__17768\,
            I => \tok.n52\
        );

    \I__3372\ : InMux
    port map (
            O => \N__17759\,
            I => \N__17756\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__17756\,
            I => \tok.n33_adj_663\
        );

    \I__3370\ : InMux
    port map (
            O => \N__17753\,
            I => \bfn_8_13_0_\
        );

    \I__3369\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17745\
        );

    \I__3368\ : InMux
    port map (
            O => \N__17749\,
            I => \N__17742\
        );

    \I__3367\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17739\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__17745\,
            I => \N__17732\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__17742\,
            I => \N__17729\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__17739\,
            I => \N__17726\
        );

    \I__3363\ : InMux
    port map (
            O => \N__17738\,
            I => \N__17723\
        );

    \I__3362\ : InMux
    port map (
            O => \N__17737\,
            I => \N__17716\
        );

    \I__3361\ : InMux
    port map (
            O => \N__17736\,
            I => \N__17716\
        );

    \I__3360\ : InMux
    port map (
            O => \N__17735\,
            I => \N__17716\
        );

    \I__3359\ : Span4Mux_h
    port map (
            O => \N__17732\,
            I => \N__17710\
        );

    \I__3358\ : Span4Mux_v
    port map (
            O => \N__17729\,
            I => \N__17710\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__17726\,
            I => \N__17703\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__17723\,
            I => \N__17703\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__17716\,
            I => \N__17703\
        );

    \I__3354\ : InMux
    port map (
            O => \N__17715\,
            I => \N__17700\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__17710\,
            I => \tok.A__15__N_129\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__17703\,
            I => \tok.A__15__N_129\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__17700\,
            I => \tok.A__15__N_129\
        );

    \I__3350\ : InMux
    port map (
            O => \N__17693\,
            I => \N__17687\
        );

    \I__3349\ : InMux
    port map (
            O => \N__17692\,
            I => \N__17687\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__17687\,
            I => \tok.A_15_N_113_3\
        );

    \I__3347\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17681\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__17681\,
            I => \tok.A_3\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__17678\,
            I => \tok.n4528_cascade_\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__17675\,
            I => \tok.n892_cascade_\
        );

    \I__3343\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17669\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__17669\,
            I => \N__17666\
        );

    \I__3341\ : Span4Mux_h
    port map (
            O => \N__17666\,
            I => \N__17663\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__17663\,
            I => \tok.n10_adj_818\
        );

    \I__3339\ : InMux
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__17657\,
            I => \N__17654\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__17654\,
            I => \tok.n13_adj_842\
        );

    \I__3336\ : InMux
    port map (
            O => \N__17651\,
            I => \N__17648\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__17648\,
            I => \tok.n8_adj_666\
        );

    \I__3334\ : InMux
    port map (
            O => \N__17645\,
            I => \N__17639\
        );

    \I__3333\ : InMux
    port map (
            O => \N__17644\,
            I => \N__17636\
        );

    \I__3332\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17631\
        );

    \I__3331\ : InMux
    port map (
            O => \N__17642\,
            I => \N__17631\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__17639\,
            I => \N__17628\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__17636\,
            I => \N__17625\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__17631\,
            I => \N__17622\
        );

    \I__3327\ : Span4Mux_s3_v
    port map (
            O => \N__17628\,
            I => \N__17617\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__17625\,
            I => \N__17617\
        );

    \I__3325\ : Span4Mux_h
    port map (
            O => \N__17622\,
            I => \N__17614\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__17617\,
            I => \tok.n8_adj_777\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__17614\,
            I => \tok.n8_adj_777\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__17609\,
            I => \tok.n4502_cascade_\
        );

    \I__3321\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17603\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__17603\,
            I => \tok.n12_adj_830\
        );

    \I__3319\ : InMux
    port map (
            O => \N__17600\,
            I => \N__17597\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__17597\,
            I => \N__17594\
        );

    \I__3317\ : Span4Mux_s3_v
    port map (
            O => \N__17594\,
            I => \N__17591\
        );

    \I__3316\ : Span4Mux_v
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__17588\,
            I => \tok.n4607\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__17585\,
            I => \tok.n2616_cascade_\
        );

    \I__3313\ : InMux
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__17579\,
            I => \N__17576\
        );

    \I__3311\ : Odrv4
    port map (
            O => \N__17576\,
            I => \tok.n10_adj_849\
        );

    \I__3310\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__17567\,
            I => \tok.n12_adj_851\
        );

    \I__3307\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17560\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__17563\,
            I => \N__17557\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__17560\,
            I => \N__17554\
        );

    \I__3304\ : InMux
    port map (
            O => \N__17557\,
            I => \N__17551\
        );

    \I__3303\ : Span4Mux_h
    port map (
            O => \N__17554\,
            I => \N__17548\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__17551\,
            I => \N__17545\
        );

    \I__3301\ : Span4Mux_h
    port map (
            O => \N__17548\,
            I => \N__17540\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__17545\,
            I => \N__17540\
        );

    \I__3299\ : Span4Mux_v
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__17537\,
            I => \tok.table_rd_1\
        );

    \I__3297\ : InMux
    port map (
            O => \N__17534\,
            I => \N__17531\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__17531\,
            I => \tok.n8_adj_850\
        );

    \I__3295\ : InMux
    port map (
            O => \N__17528\,
            I => \N__17525\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__17525\,
            I => \tok.A_4\
        );

    \I__3293\ : InMux
    port map (
            O => \N__17522\,
            I => \N__17513\
        );

    \I__3292\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17510\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__17520\,
            I => \N__17505\
        );

    \I__3290\ : CascadeMux
    port map (
            O => \N__17519\,
            I => \N__17502\
        );

    \I__3289\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17490\
        );

    \I__3288\ : InMux
    port map (
            O => \N__17517\,
            I => \N__17490\
        );

    \I__3287\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17490\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__17513\,
            I => \N__17483\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__17510\,
            I => \N__17483\
        );

    \I__3284\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17480\
        );

    \I__3283\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17475\
        );

    \I__3282\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17475\
        );

    \I__3281\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17472\
        );

    \I__3280\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17463\
        );

    \I__3279\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17463\
        );

    \I__3278\ : InMux
    port map (
            O => \N__17499\,
            I => \N__17463\
        );

    \I__3277\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17463\
        );

    \I__3276\ : InMux
    port map (
            O => \N__17497\,
            I => \N__17460\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__17490\,
            I => \N__17457\
        );

    \I__3274\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17454\
        );

    \I__3273\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17451\
        );

    \I__3272\ : Span4Mux_v
    port map (
            O => \N__17483\,
            I => \N__17442\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__17480\,
            I => \N__17442\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__17475\,
            I => \N__17442\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__17472\,
            I => \N__17442\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__17463\,
            I => \N__17439\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__17460\,
            I => \N__17436\
        );

    \I__3266\ : Span4Mux_v
    port map (
            O => \N__17457\,
            I => \N__17431\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__17454\,
            I => \N__17431\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__17451\,
            I => \N__17428\
        );

    \I__3263\ : Span4Mux_v
    port map (
            O => \N__17442\,
            I => \N__17425\
        );

    \I__3262\ : Span4Mux_v
    port map (
            O => \N__17439\,
            I => \N__17416\
        );

    \I__3261\ : Span4Mux_v
    port map (
            O => \N__17436\,
            I => \N__17416\
        );

    \I__3260\ : Span4Mux_h
    port map (
            O => \N__17431\,
            I => \N__17416\
        );

    \I__3259\ : Span4Mux_h
    port map (
            O => \N__17428\,
            I => \N__17416\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__17425\,
            I => \tok.n4051\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__17416\,
            I => \tok.n4051\
        );

    \I__3256\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__17408\,
            I => \tok.A_15_N_113_4\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__17405\,
            I => \tok.A_15_N_113_4_cascade_\
        );

    \I__3253\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__17399\,
            I => \tok.A_15_N_113_0\
        );

    \I__3251\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__17393\,
            I => \tok.A_15_N_113_6\
        );

    \I__3249\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17386\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__17389\,
            I => \N__17382\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__17386\,
            I => \N__17375\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__17385\,
            I => \N__17371\
        );

    \I__3245\ : InMux
    port map (
            O => \N__17382\,
            I => \N__17361\
        );

    \I__3244\ : InMux
    port map (
            O => \N__17381\,
            I => \N__17361\
        );

    \I__3243\ : InMux
    port map (
            O => \N__17380\,
            I => \N__17361\
        );

    \I__3242\ : InMux
    port map (
            O => \N__17379\,
            I => \N__17356\
        );

    \I__3241\ : InMux
    port map (
            O => \N__17378\,
            I => \N__17356\
        );

    \I__3240\ : Span4Mux_h
    port map (
            O => \N__17375\,
            I => \N__17353\
        );

    \I__3239\ : CascadeMux
    port map (
            O => \N__17374\,
            I => \N__17350\
        );

    \I__3238\ : InMux
    port map (
            O => \N__17371\,
            I => \N__17335\
        );

    \I__3237\ : InMux
    port map (
            O => \N__17370\,
            I => \N__17335\
        );

    \I__3236\ : InMux
    port map (
            O => \N__17369\,
            I => \N__17335\
        );

    \I__3235\ : InMux
    port map (
            O => \N__17368\,
            I => \N__17335\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__17361\,
            I => \N__17332\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17329\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__17353\,
            I => \N__17326\
        );

    \I__3231\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17315\
        );

    \I__3230\ : InMux
    port map (
            O => \N__17349\,
            I => \N__17315\
        );

    \I__3229\ : InMux
    port map (
            O => \N__17348\,
            I => \N__17315\
        );

    \I__3228\ : InMux
    port map (
            O => \N__17347\,
            I => \N__17315\
        );

    \I__3227\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17315\
        );

    \I__3226\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17312\
        );

    \I__3225\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17309\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__17335\,
            I => \N__17304\
        );

    \I__3223\ : Span4Mux_h
    port map (
            O => \N__17332\,
            I => \N__17304\
        );

    \I__3222\ : Span4Mux_h
    port map (
            O => \N__17329\,
            I => \N__17297\
        );

    \I__3221\ : Span4Mux_h
    port map (
            O => \N__17326\,
            I => \N__17297\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__17315\,
            I => \N__17297\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__17312\,
            I => \N__17294\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__17309\,
            I => \N__17289\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__17304\,
            I => \N__17289\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__17297\,
            I => \N__17286\
        );

    \I__3215\ : Odrv12
    port map (
            O => \N__17294\,
            I => \tok.n23\
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__17289\,
            I => \tok.n23\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__17286\,
            I => \tok.n23\
        );

    \I__3212\ : CEMux
    port map (
            O => \N__17279\,
            I => \N__17276\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__17276\,
            I => \N__17272\
        );

    \I__3210\ : CEMux
    port map (
            O => \N__17275\,
            I => \N__17269\
        );

    \I__3209\ : Span4Mux_v
    port map (
            O => \N__17272\,
            I => \N__17262\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__17269\,
            I => \N__17262\
        );

    \I__3207\ : CEMux
    port map (
            O => \N__17268\,
            I => \N__17259\
        );

    \I__3206\ : CEMux
    port map (
            O => \N__17267\,
            I => \N__17256\
        );

    \I__3205\ : Span4Mux_v
    port map (
            O => \N__17262\,
            I => \N__17253\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__17259\,
            I => \N__17249\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__17256\,
            I => \N__17246\
        );

    \I__3202\ : Span4Mux_h
    port map (
            O => \N__17253\,
            I => \N__17243\
        );

    \I__3201\ : CEMux
    port map (
            O => \N__17252\,
            I => \N__17240\
        );

    \I__3200\ : Span4Mux_v
    port map (
            O => \N__17249\,
            I => \N__17236\
        );

    \I__3199\ : Span4Mux_v
    port map (
            O => \N__17246\,
            I => \N__17233\
        );

    \I__3198\ : Sp12to4
    port map (
            O => \N__17243\,
            I => \N__17228\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__17240\,
            I => \N__17228\
        );

    \I__3196\ : CEMux
    port map (
            O => \N__17239\,
            I => \N__17225\
        );

    \I__3195\ : Odrv4
    port map (
            O => \N__17236\,
            I => \tok.n950\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__17233\,
            I => \tok.n950\
        );

    \I__3193\ : Odrv12
    port map (
            O => \N__17228\,
            I => \tok.n950\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__17225\,
            I => \tok.n950\
        );

    \I__3191\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__17213\,
            I => \tok.n15_adj_847\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__17210\,
            I => \N__17207\
        );

    \I__3188\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17204\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__17204\,
            I => \N__17201\
        );

    \I__3186\ : Span4Mux_h
    port map (
            O => \N__17201\,
            I => \N__17197\
        );

    \I__3185\ : InMux
    port map (
            O => \N__17200\,
            I => \N__17194\
        );

    \I__3184\ : Span4Mux_v
    port map (
            O => \N__17197\,
            I => \N__17191\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__17194\,
            I => uart_rx_data_2
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__17191\,
            I => uart_rx_data_2
        );

    \I__3181\ : InMux
    port map (
            O => \N__17186\,
            I => \N__17183\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__17183\,
            I => \tok.n12_adj_843\
        );

    \I__3179\ : InMux
    port map (
            O => \N__17180\,
            I => \N__17177\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__17177\,
            I => \N__17174\
        );

    \I__3177\ : Span4Mux_h
    port map (
            O => \N__17174\,
            I => \N__17169\
        );

    \I__3176\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17166\
        );

    \I__3175\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17163\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__17169\,
            I => capture_1
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__17166\,
            I => capture_1
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__17163\,
            I => capture_1
        );

    \I__3171\ : InMux
    port map (
            O => \N__17156\,
            I => \N__17152\
        );

    \I__3170\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17149\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__17152\,
            I => uart_rx_data_0
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__17149\,
            I => uart_rx_data_0
        );

    \I__3167\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17141\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__17141\,
            I => \N__17138\
        );

    \I__3165\ : Span4Mux_h
    port map (
            O => \N__17138\,
            I => \N__17135\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__17135\,
            I => \tok.table_rd_14\
        );

    \I__3163\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17129\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__17129\,
            I => \N__17126\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__3160\ : Span4Mux_h
    port map (
            O => \N__17123\,
            I => \N__17120\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__17120\,
            I => \tok.n16_adj_730\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__17117\,
            I => \N__17114\
        );

    \I__3157\ : InMux
    port map (
            O => \N__17114\,
            I => \N__17105\
        );

    \I__3156\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17100\
        );

    \I__3155\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17100\
        );

    \I__3154\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17091\
        );

    \I__3153\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17091\
        );

    \I__3152\ : InMux
    port map (
            O => \N__17109\,
            I => \N__17091\
        );

    \I__3151\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17091\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__17105\,
            I => \N__17079\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__17100\,
            I => \N__17079\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__17091\,
            I => \N__17079\
        );

    \I__3147\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17074\
        );

    \I__3146\ : InMux
    port map (
            O => \N__17089\,
            I => \N__17074\
        );

    \I__3145\ : InMux
    port map (
            O => \N__17088\,
            I => \N__17067\
        );

    \I__3144\ : InMux
    port map (
            O => \N__17087\,
            I => \N__17067\
        );

    \I__3143\ : InMux
    port map (
            O => \N__17086\,
            I => \N__17067\
        );

    \I__3142\ : Span4Mux_s3_v
    port map (
            O => \N__17079\,
            I => \N__17060\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__17074\,
            I => \N__17060\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__17067\,
            I => \N__17060\
        );

    \I__3139\ : Span4Mux_h
    port map (
            O => \N__17060\,
            I => \N__17057\
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__17057\,
            I => \tok.n400\
        );

    \I__3137\ : InMux
    port map (
            O => \N__17054\,
            I => \N__17051\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__17051\,
            I => \N__17048\
        );

    \I__3135\ : Span4Mux_v
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__3134\ : Span4Mux_h
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__3133\ : Sp12to4
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__3132\ : Odrv12
    port map (
            O => \N__17039\,
            I => \tok.table_wr_data_0\
        );

    \I__3131\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17033\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__17033\,
            I => \tok.n2614\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__17030\,
            I => \tok.n2614_cascade_\
        );

    \I__3128\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17024\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__3126\ : Span4Mux_h
    port map (
            O => \N__17021\,
            I => \N__17018\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__17018\,
            I => \tok.n10_adj_786\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__17015\,
            I => \tok.n6_adj_848_cascade_\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__17012\,
            I => \tok.n32_cascade_\
        );

    \I__3122\ : InMux
    port map (
            O => \N__17009\,
            I => \N__17003\
        );

    \I__3121\ : InMux
    port map (
            O => \N__17008\,
            I => \N__17003\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__17003\,
            I => uart_rx_data_1
        );

    \I__3119\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16997\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__16997\,
            I => \N__16994\
        );

    \I__3117\ : Span4Mux_v
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__3116\ : Sp12to4
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__3115\ : Odrv12
    port map (
            O => \N__16988\,
            I => \tok.table_wr_data_6\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__16985\,
            I => \N__16982\
        );

    \I__3113\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16976\
        );

    \I__3112\ : InMux
    port map (
            O => \N__16981\,
            I => \N__16976\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__16976\,
            I => \N__16972\
        );

    \I__3110\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16969\
        );

    \I__3109\ : Odrv12
    port map (
            O => \N__16972\,
            I => capture_2
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__16969\,
            I => capture_2
        );

    \I__3107\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__16961\,
            I => \N__16957\
        );

    \I__3105\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16954\
        );

    \I__3104\ : Span4Mux_h
    port map (
            O => \N__16957\,
            I => \N__16948\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__16954\,
            I => \N__16948\
        );

    \I__3102\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16945\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__16948\,
            I => \N__16939\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__16945\,
            I => \N__16936\
        );

    \I__3099\ : InMux
    port map (
            O => \N__16944\,
            I => \N__16929\
        );

    \I__3098\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16929\
        );

    \I__3097\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16929\
        );

    \I__3096\ : Span4Mux_v
    port map (
            O => \N__16939\,
            I => \N__16923\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__16936\,
            I => \N__16917\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__16929\,
            I => \N__16917\
        );

    \I__3093\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16910\
        );

    \I__3092\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16910\
        );

    \I__3091\ : InMux
    port map (
            O => \N__16926\,
            I => \N__16910\
        );

    \I__3090\ : Span4Mux_h
    port map (
            O => \N__16923\,
            I => \N__16907\
        );

    \I__3089\ : InMux
    port map (
            O => \N__16922\,
            I => \N__16904\
        );

    \I__3088\ : Span4Mux_h
    port map (
            O => \N__16917\,
            I => \N__16899\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__16910\,
            I => \N__16899\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__16907\,
            I => n4005
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__16904\,
            I => n4005
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__16899\,
            I => n4005
        );

    \I__3083\ : InMux
    port map (
            O => \N__16892\,
            I => \N__16889\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__3081\ : Span4Mux_v
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__3080\ : Span4Mux_h
    port map (
            O => \N__16883\,
            I => \N__16880\
        );

    \I__3079\ : Sp12to4
    port map (
            O => \N__16880\,
            I => \N__16877\
        );

    \I__3078\ : Odrv12
    port map (
            O => \N__16877\,
            I => \tok.table_wr_data_2\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__16874\,
            I => \tok.n18_adj_844_cascade_\
        );

    \I__3076\ : InMux
    port map (
            O => \N__16871\,
            I => \N__16868\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__16868\,
            I => \N__16865\
        );

    \I__3074\ : Span12Mux_s10_v
    port map (
            O => \N__16865\,
            I => \N__16862\
        );

    \I__3073\ : Odrv12
    port map (
            O => \N__16862\,
            I => \tok.n16_adj_845\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__16859\,
            I => \tok.n20_adj_846_cascade_\
        );

    \I__3071\ : InMux
    port map (
            O => \N__16856\,
            I => \N__16852\
        );

    \I__3070\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16849\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__16852\,
            I => \tok.A_15_N_113_2\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__16849\,
            I => \tok.A_15_N_113_2\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__16844\,
            I => \N__16841\
        );

    \I__3066\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__3064\ : Span4Mux_v
    port map (
            O => \N__16835\,
            I => \N__16832\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__16832\,
            I => \tok.tc_7\
        );

    \I__3062\ : InMux
    port map (
            O => \N__16829\,
            I => \N__16826\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__3060\ : Span4Mux_v
    port map (
            O => \N__16823\,
            I => \N__16819\
        );

    \I__3059\ : InMux
    port map (
            O => \N__16822\,
            I => \N__16816\
        );

    \I__3058\ : Odrv4
    port map (
            O => \N__16819\,
            I => \tok.C_stk.tail_1\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__16816\,
            I => \tok.C_stk.tail_1\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__16811\,
            I => \tok.C_stk.n4870_cascade_\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__16808\,
            I => \tok.ram.n4714_cascade_\
        );

    \I__3054\ : InMux
    port map (
            O => \N__16805\,
            I => \N__16802\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__16802\,
            I => \N__16798\
        );

    \I__3052\ : InMux
    port map (
            O => \N__16801\,
            I => \N__16795\
        );

    \I__3051\ : Span4Mux_s1_v
    port map (
            O => \N__16798\,
            I => \N__16789\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__16795\,
            I => \N__16789\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__16794\,
            I => \N__16784\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__16789\,
            I => \N__16781\
        );

    \I__3047\ : InMux
    port map (
            O => \N__16788\,
            I => \N__16774\
        );

    \I__3046\ : InMux
    port map (
            O => \N__16787\,
            I => \N__16774\
        );

    \I__3045\ : InMux
    port map (
            O => \N__16784\,
            I => \N__16774\
        );

    \I__3044\ : Span4Mux_h
    port map (
            O => \N__16781\,
            I => \N__16771\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__16774\,
            I => \tok.c_stk_r_1\
        );

    \I__3042\ : Odrv4
    port map (
            O => \N__16771\,
            I => \tok.c_stk_r_1\
        );

    \I__3041\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16763\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__3039\ : Span4Mux_h
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__16757\,
            I => \tok.n4690\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__16754\,
            I => \tok.n1_adj_717_cascade_\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__16751\,
            I => \tok.n5_adj_718_cascade_\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__16748\,
            I => \n92_cascade_\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__3033\ : InMux
    port map (
            O => \N__16742\,
            I => \N__16739\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__16739\,
            I => \N__16736\
        );

    \I__3031\ : Span4Mux_h
    port map (
            O => \N__16736\,
            I => \N__16733\
        );

    \I__3030\ : Odrv4
    port map (
            O => \N__16733\,
            I => \tok.tc_1\
        );

    \I__3029\ : InMux
    port map (
            O => \N__16730\,
            I => \N__16727\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__16727\,
            I => \N__16724\
        );

    \I__3027\ : Span4Mux_v
    port map (
            O => \N__16724\,
            I => \N__16721\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__16721\,
            I => \tok.n28_adj_821\
        );

    \I__3025\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16715\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__16715\,
            I => \N__16712\
        );

    \I__3023\ : Span4Mux_v
    port map (
            O => \N__16712\,
            I => \N__16709\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__16709\,
            I => \N__16705\
        );

    \I__3021\ : InMux
    port map (
            O => \N__16708\,
            I => \N__16702\
        );

    \I__3020\ : Span4Mux_h
    port map (
            O => \N__16705\,
            I => \N__16698\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__16702\,
            I => \N__16695\
        );

    \I__3018\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16692\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__16698\,
            I => capture_3
        );

    \I__3016\ : Odrv12
    port map (
            O => \N__16695\,
            I => capture_3
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__16692\,
            I => capture_3
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__16685\,
            I => \N__16682\
        );

    \I__3013\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16673\
        );

    \I__3012\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16673\
        );

    \I__3011\ : InMux
    port map (
            O => \N__16680\,
            I => \N__16673\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__16673\,
            I => \tok.n847\
        );

    \I__3009\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__3007\ : Odrv4
    port map (
            O => \N__16664\,
            I => \tok.n31\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__16661\,
            I => \tok.C_stk.n4906_cascade_\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__16658\,
            I => \tok.ram.n4699_cascade_\
        );

    \I__3004\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3002\ : Span4Mux_h
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__16646\,
            I => \tok.n4649\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__16643\,
            I => \tok.n1_adj_760_cascade_\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__16640\,
            I => \tok.n13_adj_761_cascade_\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__16637\,
            I => \tok.n28_adj_834_cascade_\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__16634\,
            I => \tok.n4604_cascade_\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__16631\,
            I => \N__16628\
        );

    \I__2995\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16625\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__16622\,
            I => \tok.n34_adj_719\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__16619\,
            I => \tok.n4610_cascade_\
        );

    \I__2991\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16610\
        );

    \I__2990\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16610\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__16610\,
            I => \tok.n37\
        );

    \I__2988\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__16604\,
            I => \N__16601\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__16598\,
            I => \N__16594\
        );

    \I__2984\ : InMux
    port map (
            O => \N__16597\,
            I => \N__16591\
        );

    \I__2983\ : Span4Mux_h
    port map (
            O => \N__16594\,
            I => \N__16588\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__16591\,
            I => \tok.table_rd_7\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__16588\,
            I => \tok.table_rd_7\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \tok.n83_adj_796_cascade_\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__2978\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16573\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__16576\,
            I => \N__16570\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__16573\,
            I => \N__16567\
        );

    \I__2975\ : InMux
    port map (
            O => \N__16570\,
            I => \N__16564\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__16567\,
            I => \tok.tail_50\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__16564\,
            I => \tok.tail_50\
        );

    \I__2972\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16553\
        );

    \I__2971\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16553\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__16553\,
            I => \tok.C_stk.tail_34\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__16550\,
            I => \N__16546\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__16549\,
            I => \N__16543\
        );

    \I__2967\ : InMux
    port map (
            O => \N__16546\,
            I => \N__16540\
        );

    \I__2966\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16537\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__16540\,
            I => \tok.tail_42\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__16537\,
            I => \tok.tail_42\
        );

    \I__2963\ : InMux
    port map (
            O => \N__16532\,
            I => \N__16526\
        );

    \I__2962\ : InMux
    port map (
            O => \N__16531\,
            I => \N__16526\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__16526\,
            I => \tok.tail_28\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__16523\,
            I => \tok.n127_cascade_\
        );

    \I__2959\ : InMux
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__16517\,
            I => \N__16513\
        );

    \I__2957\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16510\
        );

    \I__2956\ : Odrv12
    port map (
            O => \N__16513\,
            I => \tok.n4446\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__16510\,
            I => \tok.n4446\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__16505\,
            I => \tok.n4394_cascade_\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__16502\,
            I => \tok.n27_adj_863_cascade_\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__16499\,
            I => \tok.n27_adj_865_cascade_\
        );

    \I__2951\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16493\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__16493\,
            I => \tok.n27_adj_664\
        );

    \I__2949\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__16487\,
            I => \N__16484\
        );

    \I__2947\ : Span4Mux_s3_v
    port map (
            O => \N__16484\,
            I => \N__16481\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__16481\,
            I => \tok.n27_adj_866\
        );

    \I__2945\ : InMux
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__16475\,
            I => \tok.uart.sender_6\
        );

    \I__2943\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16456\
        );

    \I__2942\ : InMux
    port map (
            O => \N__16471\,
            I => \N__16456\
        );

    \I__2941\ : InMux
    port map (
            O => \N__16470\,
            I => \N__16456\
        );

    \I__2940\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16456\
        );

    \I__2939\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16449\
        );

    \I__2938\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16449\
        );

    \I__2937\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16449\
        );

    \I__2936\ : SRMux
    port map (
            O => \N__16465\,
            I => \N__16444\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__16456\,
            I => \N__16439\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__16449\,
            I => \N__16439\
        );

    \I__2933\ : InMux
    port map (
            O => \N__16448\,
            I => \N__16434\
        );

    \I__2932\ : InMux
    port map (
            O => \N__16447\,
            I => \N__16434\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__16444\,
            I => \N__16431\
        );

    \I__2930\ : Span4Mux_v
    port map (
            O => \N__16439\,
            I => \N__16428\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__16434\,
            I => \N__16424\
        );

    \I__2928\ : Span4Mux_v
    port map (
            O => \N__16431\,
            I => \N__16420\
        );

    \I__2927\ : Span4Mux_h
    port map (
            O => \N__16428\,
            I => \N__16417\
        );

    \I__2926\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16414\
        );

    \I__2925\ : Span4Mux_h
    port map (
            O => \N__16424\,
            I => \N__16411\
        );

    \I__2924\ : InMux
    port map (
            O => \N__16423\,
            I => \N__16408\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__16420\,
            I => n23
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__16417\,
            I => n23
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__16414\,
            I => n23
        );

    \I__2920\ : Odrv4
    port map (
            O => \N__16411\,
            I => n23
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__16408\,
            I => n23
        );

    \I__2918\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__16394\,
            I => \N__16391\
        );

    \I__2916\ : Odrv4
    port map (
            O => \N__16391\,
            I => \tok.uart.sender_5\
        );

    \I__2915\ : CEMux
    port map (
            O => \N__16388\,
            I => \N__16383\
        );

    \I__2914\ : CEMux
    port map (
            O => \N__16387\,
            I => \N__16380\
        );

    \I__2913\ : CEMux
    port map (
            O => \N__16386\,
            I => \N__16377\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__16383\,
            I => \N__16374\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__16380\,
            I => \N__16371\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__16377\,
            I => \N__16368\
        );

    \I__2909\ : Span4Mux_h
    port map (
            O => \N__16374\,
            I => \N__16364\
        );

    \I__2908\ : Span4Mux_h
    port map (
            O => \N__16371\,
            I => \N__16359\
        );

    \I__2907\ : Span4Mux_s3_v
    port map (
            O => \N__16368\,
            I => \N__16359\
        );

    \I__2906\ : CEMux
    port map (
            O => \N__16367\,
            I => \N__16356\
        );

    \I__2905\ : Span4Mux_h
    port map (
            O => \N__16364\,
            I => \N__16353\
        );

    \I__2904\ : Span4Mux_v
    port map (
            O => \N__16359\,
            I => \N__16348\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__16356\,
            I => \N__16348\
        );

    \I__2902\ : Span4Mux_s1_h
    port map (
            O => \N__16353\,
            I => \N__16345\
        );

    \I__2901\ : Span4Mux_h
    port map (
            O => \N__16348\,
            I => \N__16342\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__16345\,
            I => \tok.uart.n964\
        );

    \I__2899\ : Odrv4
    port map (
            O => \N__16342\,
            I => \tok.uart.n964\
        );

    \I__2898\ : InMux
    port map (
            O => \N__16337\,
            I => \N__16334\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__2896\ : Span4Mux_v
    port map (
            O => \N__16331\,
            I => \N__16328\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__16328\,
            I => \tok.n16_adj_706\
        );

    \I__2894\ : InMux
    port map (
            O => \N__16325\,
            I => \N__16322\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__16322\,
            I => \tok.n14_adj_707\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__16319\,
            I => \tok.n20_adj_708_cascade_\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__16316\,
            I => \tok.n22_adj_709_cascade_\
        );

    \I__2890\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16310\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__16310\,
            I => \tok.A_15_N_113_5\
        );

    \I__2888\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16304\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__16304\,
            I => \N__16301\
        );

    \I__2886\ : Span4Mux_v
    port map (
            O => \N__16301\,
            I => \N__16298\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__16298\,
            I => \tok.n10_adj_806\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__16295\,
            I => \tok.n13_adj_813_cascade_\
        );

    \I__2883\ : InMux
    port map (
            O => \N__16292\,
            I => \N__16289\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__16289\,
            I => \tok.n18_adj_819\
        );

    \I__2881\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16283\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__16283\,
            I => \tok.n15_adj_823\
        );

    \I__2879\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16277\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__16277\,
            I => \tok.uart.sender_3\
        );

    \I__2877\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16271\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__16271\,
            I => \tok.A_0\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__16268\,
            I => \N__16265\
        );

    \I__2874\ : InMux
    port map (
            O => \N__16265\,
            I => \N__16262\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__16262\,
            I => \N__16259\
        );

    \I__2872\ : Odrv12
    port map (
            O => \N__16259\,
            I => sender_2
        );

    \I__2871\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16253\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__16253\,
            I => \N__16250\
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__16250\,
            I => \tok.A_2\
        );

    \I__2868\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__16244\,
            I => \tok.uart.sender_4\
        );

    \I__2866\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16238\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__16238\,
            I => \N__16235\
        );

    \I__2864\ : Span4Mux_h
    port map (
            O => \N__16235\,
            I => \N__16232\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__16232\,
            I => \tok.n10_adj_783\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__16229\,
            I => \tok.n14_adj_779_cascade_\
        );

    \I__2861\ : InMux
    port map (
            O => \N__16226\,
            I => \N__16223\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__16223\,
            I => \N__16220\
        );

    \I__2859\ : Span4Mux_h
    port map (
            O => \N__16220\,
            I => \N__16217\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__16217\,
            I => \tok.n20_adj_781\
        );

    \I__2857\ : CascadeMux
    port map (
            O => \N__16214\,
            I => \tok.n22_adj_784_cascade_\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__16211\,
            I => \tok.A_15_N_113_6_cascade_\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__16208\,
            I => \tok.A_6_cascade_\
        );

    \I__2854\ : InMux
    port map (
            O => \N__16205\,
            I => \N__16202\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__16202\,
            I => \N__16199\
        );

    \I__2852\ : Span4Mux_h
    port map (
            O => \N__16199\,
            I => \N__16196\
        );

    \I__2851\ : Span4Mux_v
    port map (
            O => \N__16196\,
            I => \N__16193\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__16193\,
            I => \N__16190\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__16190\,
            I => \tok.uart.sender_9\
        );

    \I__2848\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__16184\,
            I => \tok.uart.sender_8\
        );

    \I__2846\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16178\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__16178\,
            I => \tok.A_5\
        );

    \I__2844\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16172\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__16172\,
            I => \tok.uart.sender_7\
        );

    \I__2842\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16166\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__16166\,
            I => \tok.n2\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__16163\,
            I => \tok.n19_cascade_\
        );

    \I__2839\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16157\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__16157\,
            I => \N__16154\
        );

    \I__2837\ : Span4Mux_h
    port map (
            O => \N__16154\,
            I => \N__16151\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__16151\,
            I => \tok.n6_adj_684\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__16148\,
            I => \tok.n22_adj_683_cascade_\
        );

    \I__2834\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16142\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__16142\,
            I => \tok.n4544\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__16139\,
            I => \tok.A_15_N_113_0_cascade_\
        );

    \I__2831\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16133\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__16133\,
            I => \tok.n4520\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__16130\,
            I => \tok.n46_cascade_\
        );

    \I__2828\ : InMux
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__16124\,
            I => \N__16121\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__16121\,
            I => \tok.A_15_N_113_1\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__16118\,
            I => \tok.A_15_N_113_1_cascade_\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__16115\,
            I => \tok.A_1_cascade_\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__16112\,
            I => \tok.A__15__N_129_cascade_\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__16109\,
            I => \tok.n27_adj_867_cascade_\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__16106\,
            I => \N__16103\
        );

    \I__2820\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16100\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__16100\,
            I => \tok.n1\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__16097\,
            I => \tok.n14_adj_678_cascade_\
        );

    \I__2817\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16091\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__16091\,
            I => \tok.n18_adj_859\
        );

    \I__2815\ : InMux
    port map (
            O => \N__16088\,
            I => \N__16085\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__16085\,
            I => \N__16082\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__16082\,
            I => \tok.n22_adj_855\
        );

    \I__2812\ : InMux
    port map (
            O => \N__16079\,
            I => \N__16076\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__16076\,
            I => \N__16072\
        );

    \I__2810\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16069\
        );

    \I__2809\ : Span4Mux_h
    port map (
            O => \N__16072\,
            I => \N__16066\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__16069\,
            I => \tok.n880\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__16066\,
            I => \tok.n880\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__16061\,
            I => \tok.n23_cascade_\
        );

    \I__2805\ : InMux
    port map (
            O => \N__16058\,
            I => \N__16055\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__16055\,
            I => \tok.n23_adj_856\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__16052\,
            I => \N__16043\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__16051\,
            I => \N__16040\
        );

    \I__2801\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16034\
        );

    \I__2800\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16034\
        );

    \I__2799\ : InMux
    port map (
            O => \N__16048\,
            I => \N__16025\
        );

    \I__2798\ : InMux
    port map (
            O => \N__16047\,
            I => \N__16025\
        );

    \I__2797\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16025\
        );

    \I__2796\ : InMux
    port map (
            O => \N__16043\,
            I => \N__16025\
        );

    \I__2795\ : InMux
    port map (
            O => \N__16040\,
            I => \N__16020\
        );

    \I__2794\ : InMux
    port map (
            O => \N__16039\,
            I => \N__16020\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__16034\,
            I => \N__16015\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__16025\,
            I => \N__16015\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__16020\,
            I => \tok.n64\
        );

    \I__2790\ : Odrv12
    port map (
            O => \N__16015\,
            I => \tok.n64\
        );

    \I__2789\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16003\
        );

    \I__2788\ : InMux
    port map (
            O => \N__16009\,
            I => \N__16003\
        );

    \I__2787\ : InMux
    port map (
            O => \N__16008\,
            I => \N__15998\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__16003\,
            I => \N__15995\
        );

    \I__2785\ : InMux
    port map (
            O => \N__16002\,
            I => \N__15990\
        );

    \I__2784\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15990\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__15998\,
            I => \tok.n1_adj_802\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__15995\,
            I => \tok.n1_adj_802\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__15990\,
            I => \tok.n1_adj_802\
        );

    \I__2780\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15980\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__15980\,
            I => \N__15977\
        );

    \I__2778\ : Odrv12
    port map (
            O => \N__15977\,
            I => \tok.depth_2\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__15974\,
            I => \tok.depth_0_cascade_\
        );

    \I__2776\ : InMux
    port map (
            O => \N__15971\,
            I => \N__15968\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__15968\,
            I => \N__15965\
        );

    \I__2774\ : Odrv12
    port map (
            O => \N__15965\,
            I => \tok.n6_adj_853\
        );

    \I__2773\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15956\
        );

    \I__2772\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15956\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__15956\,
            I => \tok.n6_adj_832\
        );

    \I__2770\ : InMux
    port map (
            O => \N__15953\,
            I => \N__15950\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__15950\,
            I => \tok.n4504\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__15947\,
            I => \tok.n4432_cascade_\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__15944\,
            I => \N__15936\
        );

    \I__2766\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15931\
        );

    \I__2765\ : InMux
    port map (
            O => \N__15942\,
            I => \N__15931\
        );

    \I__2764\ : InMux
    port map (
            O => \N__15941\,
            I => \N__15928\
        );

    \I__2763\ : InMux
    port map (
            O => \N__15940\,
            I => \N__15921\
        );

    \I__2762\ : InMux
    port map (
            O => \N__15939\,
            I => \N__15921\
        );

    \I__2761\ : InMux
    port map (
            O => \N__15936\,
            I => \N__15921\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__15931\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__15928\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__15921\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__15914\,
            I => \tok.n1_adj_802_cascade_\
        );

    \I__2756\ : InMux
    port map (
            O => \N__15911\,
            I => \N__15902\
        );

    \I__2755\ : InMux
    port map (
            O => \N__15910\,
            I => \N__15902\
        );

    \I__2754\ : InMux
    port map (
            O => \N__15909\,
            I => \N__15902\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__15902\,
            I => \tok.n189\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__15899\,
            I => \N__15891\
        );

    \I__2751\ : InMux
    port map (
            O => \N__15898\,
            I => \N__15886\
        );

    \I__2750\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15879\
        );

    \I__2749\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15879\
        );

    \I__2748\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15879\
        );

    \I__2747\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15870\
        );

    \I__2746\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15870\
        );

    \I__2745\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15870\
        );

    \I__2744\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15870\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__15886\,
            I => \tok.n62\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__15879\,
            I => \tok.n62\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__15870\,
            I => \tok.n62\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__15863\,
            I => \tok.n189_cascade_\
        );

    \I__2739\ : InMux
    port map (
            O => \N__15860\,
            I => \N__15853\
        );

    \I__2738\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15853\
        );

    \I__2737\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15850\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__15853\,
            I => \tok.n4_adj_809\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__15850\,
            I => \tok.n4_adj_809\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__15845\,
            I => \tok.n27_adj_793_cascade_\
        );

    \I__2733\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15839\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__15839\,
            I => \tok.n25_adj_794\
        );

    \I__2731\ : InMux
    port map (
            O => \N__15836\,
            I => \N__15833\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__15833\,
            I => \tok.n26_adj_792\
        );

    \I__2729\ : InMux
    port map (
            O => \N__15830\,
            I => \N__15827\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__15827\,
            I => \tok.n28_adj_791\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__15824\,
            I => \N__15820\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__15823\,
            I => \N__15814\
        );

    \I__2725\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15808\
        );

    \I__2724\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15808\
        );

    \I__2723\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15803\
        );

    \I__2722\ : InMux
    port map (
            O => \N__15817\,
            I => \N__15803\
        );

    \I__2721\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15798\
        );

    \I__2720\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15798\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__15808\,
            I => \tok.n63\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__15803\,
            I => \tok.n63\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__15798\,
            I => \tok.n63\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__15791\,
            I => \tok.A_stk_delta_1__N_4_cascade_\
        );

    \I__2715\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15778\
        );

    \I__2714\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15778\
        );

    \I__2713\ : InMux
    port map (
            O => \N__15786\,
            I => \N__15771\
        );

    \I__2712\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15771\
        );

    \I__2711\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15771\
        );

    \I__2710\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15768\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__15778\,
            I => \tok.n61\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__15771\,
            I => \tok.n61\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__15768\,
            I => \tok.n61\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__15761\,
            I => \tok.n4_adj_809_cascade_\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__15758\,
            I => \tok.depth_3_cascade_\
        );

    \I__2704\ : InMux
    port map (
            O => \N__15755\,
            I => \N__15752\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__15752\,
            I => \tok.depth_1\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__15749\,
            I => \tok.n4554_cascade_\
        );

    \I__2701\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15736\
        );

    \I__2700\ : InMux
    port map (
            O => \N__15745\,
            I => \N__15733\
        );

    \I__2699\ : InMux
    port map (
            O => \N__15744\,
            I => \N__15728\
        );

    \I__2698\ : InMux
    port map (
            O => \N__15743\,
            I => \N__15725\
        );

    \I__2697\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15721\
        );

    \I__2696\ : InMux
    port map (
            O => \N__15741\,
            I => \N__15716\
        );

    \I__2695\ : InMux
    port map (
            O => \N__15740\,
            I => \N__15713\
        );

    \I__2694\ : InMux
    port map (
            O => \N__15739\,
            I => \N__15709\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__15736\,
            I => \N__15706\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__15733\,
            I => \N__15703\
        );

    \I__2691\ : InMux
    port map (
            O => \N__15732\,
            I => \N__15700\
        );

    \I__2690\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15697\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__15728\,
            I => \N__15692\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__15725\,
            I => \N__15692\
        );

    \I__2687\ : InMux
    port map (
            O => \N__15724\,
            I => \N__15689\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__15721\,
            I => \N__15686\
        );

    \I__2685\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15683\
        );

    \I__2684\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15678\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__15716\,
            I => \N__15673\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__15713\,
            I => \N__15673\
        );

    \I__2681\ : InMux
    port map (
            O => \N__15712\,
            I => \N__15670\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__15709\,
            I => \N__15667\
        );

    \I__2679\ : Span4Mux_s3_h
    port map (
            O => \N__15706\,
            I => \N__15658\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__15703\,
            I => \N__15658\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__15700\,
            I => \N__15658\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__15697\,
            I => \N__15658\
        );

    \I__2675\ : Span4Mux_s3_h
    port map (
            O => \N__15692\,
            I => \N__15653\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__15689\,
            I => \N__15653\
        );

    \I__2673\ : Span4Mux_v
    port map (
            O => \N__15686\,
            I => \N__15650\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__15683\,
            I => \N__15647\
        );

    \I__2671\ : InMux
    port map (
            O => \N__15682\,
            I => \N__15644\
        );

    \I__2670\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15641\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__15678\,
            I => \N__15638\
        );

    \I__2668\ : Span12Mux_s7_h
    port map (
            O => \N__15673\,
            I => \N__15635\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__15670\,
            I => \N__15632\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__15667\,
            I => \N__15627\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__15658\,
            I => \N__15627\
        );

    \I__2664\ : Span4Mux_h
    port map (
            O => \N__15653\,
            I => \N__15624\
        );

    \I__2663\ : Span4Mux_h
    port map (
            O => \N__15650\,
            I => \N__15615\
        );

    \I__2662\ : Span4Mux_v
    port map (
            O => \N__15647\,
            I => \N__15615\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__15644\,
            I => \N__15615\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__15641\,
            I => \N__15615\
        );

    \I__2659\ : Odrv12
    port map (
            O => \N__15638\,
            I => \tok.n237\
        );

    \I__2658\ : Odrv12
    port map (
            O => \N__15635\,
            I => \tok.n237\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__15632\,
            I => \tok.n237\
        );

    \I__2656\ : Odrv4
    port map (
            O => \N__15627\,
            I => \tok.n237\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__15624\,
            I => \tok.n237\
        );

    \I__2654\ : Odrv4
    port map (
            O => \N__15615\,
            I => \tok.n237\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__15602\,
            I => \tok.n875_cascade_\
        );

    \I__2652\ : InMux
    port map (
            O => \N__15599\,
            I => \N__15594\
        );

    \I__2651\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15591\
        );

    \I__2650\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15588\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__15594\,
            I => \N__15585\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__15591\,
            I => \tok.n2562\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__15588\,
            I => \tok.n2562\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__15585\,
            I => \tok.n2562\
        );

    \I__2645\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15572\
        );

    \I__2644\ : InMux
    port map (
            O => \N__15577\,
            I => \N__15572\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__15572\,
            I => \tok.n2503\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__15569\,
            I => \tok.n2562_cascade_\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__15566\,
            I => \tok.n4474_cascade_\
        );

    \I__2640\ : InMux
    port map (
            O => \N__15563\,
            I => \N__15560\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__15560\,
            I => \tok.n875\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__15557\,
            I => \tok.n20_adj_772_cascade_\
        );

    \I__2637\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15548\
        );

    \I__2636\ : InMux
    port map (
            O => \N__15553\,
            I => \N__15548\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__15548\,
            I => \tok.tail_9\
        );

    \I__2634\ : InMux
    port map (
            O => \N__15545\,
            I => \N__15539\
        );

    \I__2633\ : InMux
    port map (
            O => \N__15544\,
            I => \N__15539\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__15539\,
            I => \tok.C_stk.tail_17\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__15536\,
            I => \N__15533\
        );

    \I__2630\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15527\
        );

    \I__2629\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15527\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__15527\,
            I => \N__15524\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__15524\,
            I => \tok.tail_25\
        );

    \I__2626\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15515\
        );

    \I__2625\ : InMux
    port map (
            O => \N__15520\,
            I => \N__15515\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__15515\,
            I => \tok.C_stk.tail_33\
        );

    \I__2623\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15508\
        );

    \I__2622\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15505\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__15508\,
            I => \tok.tail_57\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__15505\,
            I => \tok.tail_57\
        );

    \I__2619\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15494\
        );

    \I__2618\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15494\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__15494\,
            I => \tok.tail_41\
        );

    \I__2616\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15487\
        );

    \I__2615\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15484\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__15487\,
            I => \tok.tail_49\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__15484\,
            I => \tok.tail_49\
        );

    \I__2612\ : InMux
    port map (
            O => \N__15479\,
            I => \N__15475\
        );

    \I__2611\ : InMux
    port map (
            O => \N__15478\,
            I => \N__15472\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__15475\,
            I => \tok.tail_58\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__15472\,
            I => \tok.tail_58\
        );

    \I__2608\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15464\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__15464\,
            I => \N__15461\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__15461\,
            I => \tok.n16_adj_820\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__15458\,
            I => \tok.n20_adj_822_cascade_\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__15455\,
            I => \tok.A_15_N_113_5_cascade_\
        );

    \I__2603\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15449\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__15449\,
            I => \N__15446\
        );

    \I__2601\ : Span4Mux_v
    port map (
            O => \N__15446\,
            I => \N__15443\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__15443\,
            I => \tok.n297\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__15440\,
            I => \N__15437\
        );

    \I__2598\ : InMux
    port map (
            O => \N__15437\,
            I => \N__15434\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__15434\,
            I => \tok.n208\
        );

    \I__2596\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15428\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__15425\,
            I => \N__15422\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__15422\,
            I => \tok.n20_adj_858\
        );

    \I__2592\ : InMux
    port map (
            O => \N__15419\,
            I => \N__15416\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__15416\,
            I => \N__15413\
        );

    \I__2590\ : Span4Mux_h
    port map (
            O => \N__15413\,
            I => \N__15410\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__15410\,
            I => \tok.n299\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__15407\,
            I => \tok.n27_adj_644_cascade_\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__15404\,
            I => \tok.n2_adj_720_cascade_\
        );

    \I__2586\ : InMux
    port map (
            O => \N__15401\,
            I => \N__15398\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__15398\,
            I => \tok.n14_adj_722\
        );

    \I__2584\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15392\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__15392\,
            I => \N__15389\
        );

    \I__2582\ : Span12Mux_s11_v
    port map (
            O => \N__15389\,
            I => \N__15386\
        );

    \I__2581\ : Odrv12
    port map (
            O => \N__15386\,
            I => \tok.n6_adj_731\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__15383\,
            I => \tok.n13_adj_726_cascade_\
        );

    \I__2579\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__15377\,
            I => \N__15374\
        );

    \I__2577\ : Odrv12
    port map (
            O => \N__15374\,
            I => \tok.n12_adj_723\
        );

    \I__2576\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15368\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__15368\,
            I => \N__15365\
        );

    \I__2574\ : Span4Mux_v
    port map (
            O => \N__15365\,
            I => \N__15362\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__15362\,
            I => \tok.n4661\
        );

    \I__2572\ : CascadeMux
    port map (
            O => \N__15359\,
            I => \tok.n20_adj_732_cascade_\
        );

    \I__2571\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__15353\,
            I => \N__15350\
        );

    \I__2569\ : Odrv12
    port map (
            O => \N__15350\,
            I => \tok.n4658\
        );

    \I__2568\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__15344\,
            I => \tok.n9_adj_728\
        );

    \I__2566\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15338\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__15338\,
            I => \N__15335\
        );

    \I__2564\ : Span4Mux_v
    port map (
            O => \N__15335\,
            I => \N__15332\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__15332\,
            I => \tok.n184\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__2561\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15323\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__15323\,
            I => \N__15319\
        );

    \I__2559\ : InMux
    port map (
            O => \N__15322\,
            I => \N__15316\
        );

    \I__2558\ : Span4Mux_h
    port map (
            O => \N__15319\,
            I => \N__15313\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__15316\,
            I => uart_rx_data_5
        );

    \I__2556\ : Odrv4
    port map (
            O => \N__15313\,
            I => uart_rx_data_5
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__15308\,
            I => \tok.n12_adj_815_cascade_\
        );

    \I__2554\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15302\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__15302\,
            I => \tok.n4653\
        );

    \I__2552\ : InMux
    port map (
            O => \N__15299\,
            I => \N__15296\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__15296\,
            I => \tok.n4671\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__15293\,
            I => \N__15290\
        );

    \I__2549\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15287\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__15287\,
            I => \tok.n18_adj_672\
        );

    \I__2547\ : InMux
    port map (
            O => \N__15284\,
            I => \N__15281\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__15281\,
            I => \N__15278\
        );

    \I__2545\ : Span4Mux_v
    port map (
            O => \N__15278\,
            I => \N__15275\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__15275\,
            I => \tok.n6_adj_676\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__15272\,
            I => \tok.n20_adj_674_cascade_\
        );

    \I__2542\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15266\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__15266\,
            I => \N__15263\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__15263\,
            I => \N__15260\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__15260\,
            I => \tok.n16_adj_673\
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__15257\,
            I => \tok.n4676_cascade_\
        );

    \I__2537\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15251\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__15251\,
            I => \tok.n12_adj_744\
        );

    \I__2535\ : InMux
    port map (
            O => \N__15248\,
            I => \N__15245\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__15245\,
            I => \tok.n4524\
        );

    \I__2533\ : InMux
    port map (
            O => \N__15242\,
            I => \N__15239\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__15239\,
            I => \tok.n12_adj_670\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__15236\,
            I => \tok.n15_cascade_\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__2529\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15227\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__15227\,
            I => \tok.n183\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \N__15221\
        );

    \I__2526\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15217\
        );

    \I__2525\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15214\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__15217\,
            I => \N__15211\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__15214\,
            I => \N__15208\
        );

    \I__2522\ : Span4Mux_h
    port map (
            O => \N__15211\,
            I => \N__15205\
        );

    \I__2521\ : Span4Mux_v
    port map (
            O => \N__15208\,
            I => \N__15202\
        );

    \I__2520\ : Span4Mux_v
    port map (
            O => \N__15205\,
            I => \N__15199\
        );

    \I__2519\ : Odrv4
    port map (
            O => \N__15202\,
            I => \tok.table_rd_6\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__15199\,
            I => \tok.table_rd_6\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__15194\,
            I => \tok.n16_adj_778_cascade_\
        );

    \I__2516\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15188\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__15188\,
            I => \N__15185\
        );

    \I__2514\ : Span4Mux_h
    port map (
            O => \N__15185\,
            I => \N__15182\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__15182\,
            I => \tok.n6_adj_780\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__15179\,
            I => \N__15176\
        );

    \I__2511\ : InMux
    port map (
            O => \N__15176\,
            I => \N__15173\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__15173\,
            I => \N__15170\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__15170\,
            I => \tok.table_rd_13\
        );

    \I__2508\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15164\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__15164\,
            I => \N__15161\
        );

    \I__2506\ : Span4Mux_h
    port map (
            O => \N__15161\,
            I => \N__15158\
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__15158\,
            I => \tok.table_rd_10\
        );

    \I__2504\ : InMux
    port map (
            O => \N__15155\,
            I => \N__15152\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__15152\,
            I => \tok.n10_adj_671\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__15149\,
            I => \tok.n14_adj_669_cascade_\
        );

    \I__2501\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15143\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__15143\,
            I => \N__15140\
        );

    \I__2499\ : Span4Mux_h
    port map (
            O => \N__15140\,
            I => \N__15137\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__15137\,
            I => \tok.table_rd_11\
        );

    \I__2497\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15131\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__15131\,
            I => \N__15128\
        );

    \I__2495\ : Span4Mux_h
    port map (
            O => \N__15128\,
            I => \N__15125\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__15125\,
            I => \tok.n16_adj_691\
        );

    \I__2493\ : InMux
    port map (
            O => \N__15122\,
            I => \N__15118\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__15121\,
            I => \N__15115\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__15118\,
            I => \N__15112\
        );

    \I__2490\ : InMux
    port map (
            O => \N__15115\,
            I => \N__15109\
        );

    \I__2489\ : Span4Mux_h
    port map (
            O => \N__15112\,
            I => \N__15106\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__15109\,
            I => \tok.key_rd_4\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__15106\,
            I => \tok.key_rd_4\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__15101\,
            I => \N__15098\
        );

    \I__2485\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15095\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__15095\,
            I => \N__15091\
        );

    \I__2483\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15088\
        );

    \I__2482\ : Span4Mux_h
    port map (
            O => \N__15091\,
            I => \N__15085\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__15088\,
            I => \tok.key_rd_1\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__15085\,
            I => \tok.key_rd_1\
        );

    \I__2479\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__15077\,
            I => \tok.n18_adj_756\
        );

    \I__2477\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15071\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__15071\,
            I => \N__15068\
        );

    \I__2475\ : Span4Mux_h
    port map (
            O => \N__15068\,
            I => \N__15064\
        );

    \I__2474\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15061\
        );

    \I__2473\ : Span4Mux_s3_h
    port map (
            O => \N__15064\,
            I => \N__15058\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__15061\,
            I => \tok.key_rd_0\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__15058\,
            I => \tok.key_rd_0\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__15053\,
            I => \N__15050\
        );

    \I__2469\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15047\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__15047\,
            I => \N__15044\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__15044\,
            I => \N__15040\
        );

    \I__2466\ : InMux
    port map (
            O => \N__15043\,
            I => \N__15037\
        );

    \I__2465\ : Span4Mux_h
    port map (
            O => \N__15040\,
            I => \N__15034\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__15037\,
            I => \tok.key_rd_6\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__15034\,
            I => \tok.key_rd_6\
        );

    \I__2462\ : InMux
    port map (
            O => \N__15029\,
            I => \N__15026\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__15026\,
            I => \N__15023\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__15023\,
            I => \tok.n4645\
        );

    \I__2459\ : InMux
    port map (
            O => \N__15020\,
            I => \N__15017\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__15017\,
            I => \N__15014\
        );

    \I__2457\ : Span4Mux_h
    port map (
            O => \N__15014\,
            I => \N__15011\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__15011\,
            I => \tok.n13_adj_657\
        );

    \I__2455\ : InMux
    port map (
            O => \N__15008\,
            I => \N__15005\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__15005\,
            I => \tok.n10_adj_656\
        );

    \I__2453\ : InMux
    port map (
            O => \N__15002\,
            I => \N__14999\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__14999\,
            I => \N__14996\
        );

    \I__2451\ : Span4Mux_h
    port map (
            O => \N__14996\,
            I => \N__14993\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__14993\,
            I => \tok.table_rd_9\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__14990\,
            I => \tok.n30_cascade_\
        );

    \I__2448\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14984\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__14984\,
            I => \N__14981\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__14981\,
            I => \N__14978\
        );

    \I__2445\ : Span4Mux_h
    port map (
            O => \N__14978\,
            I => \N__14975\
        );

    \I__2444\ : Odrv4
    port map (
            O => \N__14975\,
            I => \tok.n12_adj_659\
        );

    \I__2443\ : CEMux
    port map (
            O => \N__14972\,
            I => \N__14969\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__14969\,
            I => \N__14966\
        );

    \I__2441\ : Odrv12
    port map (
            O => \N__14966\,
            I => \tok.uart.n922\
        );

    \I__2440\ : InMux
    port map (
            O => \N__14963\,
            I => \N__14960\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__14960\,
            I => \N__14957\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__14957\,
            I => \N__14954\
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__14954\,
            I => \tok.n301\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__14951\,
            I => \tok.n19_adj_860_cascade_\
        );

    \I__2435\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14945\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__14945\,
            I => \tok.n17_adj_861\
        );

    \I__2433\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14939\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__14939\,
            I => \tok.n29_adj_864\
        );

    \I__2431\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14933\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__14933\,
            I => \N__14930\
        );

    \I__2429\ : Span4Mux_h
    port map (
            O => \N__14930\,
            I => \N__14926\
        );

    \I__2428\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14923\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__14926\,
            I => \N__14918\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__14923\,
            I => \N__14918\
        );

    \I__2425\ : Span4Mux_h
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__2424\ : Span4Mux_s2_h
    port map (
            O => \N__14915\,
            I => \N__14911\
        );

    \I__2423\ : InMux
    port map (
            O => \N__14914\,
            I => \N__14908\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__14911\,
            I => capture_8
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__14908\,
            I => capture_8
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__14903\,
            I => \N__14900\
        );

    \I__2419\ : InMux
    port map (
            O => \N__14900\,
            I => \N__14896\
        );

    \I__2418\ : InMux
    port map (
            O => \N__14899\,
            I => \N__14893\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__14896\,
            I => uart_rx_data_7
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__14893\,
            I => uart_rx_data_7
        );

    \I__2415\ : InMux
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__2413\ : Span4Mux_v
    port map (
            O => \N__14882\,
            I => \N__14879\
        );

    \I__2412\ : Span4Mux_h
    port map (
            O => \N__14879\,
            I => \N__14876\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__14876\,
            I => \tok.table_wr_data_10\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__14873\,
            I => \N__14870\
        );

    \I__2409\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14867\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__14867\,
            I => \N__14864\
        );

    \I__2407\ : Span4Mux_h
    port map (
            O => \N__14864\,
            I => \N__14861\
        );

    \I__2406\ : Span4Mux_v
    port map (
            O => \N__14861\,
            I => \N__14858\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__14858\,
            I => \tok.n293\
        );

    \I__2404\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14852\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__14852\,
            I => \N__14849\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__14849\,
            I => \tok.n2634\
        );

    \I__2401\ : SRMux
    port map (
            O => \N__14846\,
            I => \N__14842\
        );

    \I__2400\ : SRMux
    port map (
            O => \N__14845\,
            I => \N__14839\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__14842\,
            I => \N__14834\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__14839\,
            I => \N__14834\
        );

    \I__2397\ : Span4Mux_v
    port map (
            O => \N__14834\,
            I => \N__14831\
        );

    \I__2396\ : Span4Mux_s3_h
    port map (
            O => \N__14831\,
            I => \N__14828\
        );

    \I__2395\ : Span4Mux_h
    port map (
            O => \N__14828\,
            I => \N__14825\
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__14825\,
            I => \tok.write_slot\
        );

    \I__2393\ : InMux
    port map (
            O => \N__14822\,
            I => \N__14819\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__14819\,
            I => \N__14816\
        );

    \I__2391\ : Span4Mux_h
    port map (
            O => \N__14816\,
            I => \N__14813\
        );

    \I__2390\ : Span4Mux_s3_h
    port map (
            O => \N__14813\,
            I => \N__14810\
        );

    \I__2389\ : Span4Mux_h
    port map (
            O => \N__14810\,
            I => \N__14807\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__14807\,
            I => \tok.table_wr_data_5\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__14804\,
            I => \tok.n83_adj_716_cascade_\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__14801\,
            I => \tok.n12_adj_740_cascade_\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__14798\,
            I => \tok.n12_adj_801_cascade_\
        );

    \I__2384\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14792\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__14792\,
            I => \tok.n284\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__14789\,
            I => \tok.n284_cascade_\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__14786\,
            I => \tok.n182_cascade_\
        );

    \I__2380\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14780\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__14780\,
            I => \N__14777\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__14777\,
            I => \N__14774\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__14774\,
            I => \tok.n12_adj_766\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__14771\,
            I => \N__14768\
        );

    \I__2375\ : InMux
    port map (
            O => \N__14768\,
            I => \N__14765\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__14765\,
            I => \N__14762\
        );

    \I__2373\ : Span4Mux_h
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__2372\ : Odrv4
    port map (
            O => \N__14759\,
            I => \tok.n24_adj_854\
        );

    \I__2371\ : InMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__14753\,
            I => \N__14750\
        );

    \I__2369\ : Span12Mux_s9_h
    port map (
            O => \N__14750\,
            I => \N__14747\
        );

    \I__2368\ : Odrv12
    port map (
            O => \N__14747\,
            I => \tok.n21_adj_857\
        );

    \I__2367\ : CascadeMux
    port map (
            O => \N__14744\,
            I => \tok.n30_adj_862_cascade_\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__14741\,
            I => \n29_cascade_\
        );

    \I__2365\ : CEMux
    port map (
            O => \N__14738\,
            I => \N__14733\
        );

    \I__2364\ : CEMux
    port map (
            O => \N__14737\,
            I => \N__14730\
        );

    \I__2363\ : CEMux
    port map (
            O => \N__14736\,
            I => \N__14723\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__14733\,
            I => \N__14717\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__14730\,
            I => \N__14717\
        );

    \I__2360\ : CEMux
    port map (
            O => \N__14729\,
            I => \N__14714\
        );

    \I__2359\ : CEMux
    port map (
            O => \N__14728\,
            I => \N__14709\
        );

    \I__2358\ : CEMux
    port map (
            O => \N__14727\,
            I => \N__14704\
        );

    \I__2357\ : CEMux
    port map (
            O => \N__14726\,
            I => \N__14700\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__14723\,
            I => \N__14697\
        );

    \I__2355\ : CEMux
    port map (
            O => \N__14722\,
            I => \N__14694\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__14717\,
            I => \N__14689\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__14714\,
            I => \N__14689\
        );

    \I__2352\ : CEMux
    port map (
            O => \N__14713\,
            I => \N__14686\
        );

    \I__2351\ : CEMux
    port map (
            O => \N__14712\,
            I => \N__14683\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__14709\,
            I => \N__14677\
        );

    \I__2349\ : CEMux
    port map (
            O => \N__14708\,
            I => \N__14674\
        );

    \I__2348\ : CEMux
    port map (
            O => \N__14707\,
            I => \N__14671\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__14704\,
            I => \N__14668\
        );

    \I__2346\ : CEMux
    port map (
            O => \N__14703\,
            I => \N__14665\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__14700\,
            I => \N__14661\
        );

    \I__2344\ : Span4Mux_s3_h
    port map (
            O => \N__14697\,
            I => \N__14656\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__14694\,
            I => \N__14656\
        );

    \I__2342\ : Span4Mux_s2_h
    port map (
            O => \N__14689\,
            I => \N__14651\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__14686\,
            I => \N__14651\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__14683\,
            I => \N__14648\
        );

    \I__2339\ : CEMux
    port map (
            O => \N__14682\,
            I => \N__14645\
        );

    \I__2338\ : CEMux
    port map (
            O => \N__14681\,
            I => \N__14642\
        );

    \I__2337\ : CEMux
    port map (
            O => \N__14680\,
            I => \N__14639\
        );

    \I__2336\ : Span4Mux_h
    port map (
            O => \N__14677\,
            I => \N__14634\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__14674\,
            I => \N__14634\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__14671\,
            I => \N__14631\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__14668\,
            I => \N__14626\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__14665\,
            I => \N__14626\
        );

    \I__2331\ : CEMux
    port map (
            O => \N__14664\,
            I => \N__14623\
        );

    \I__2330\ : Span4Mux_h
    port map (
            O => \N__14661\,
            I => \N__14620\
        );

    \I__2329\ : Span4Mux_h
    port map (
            O => \N__14656\,
            I => \N__14617\
        );

    \I__2328\ : Span4Mux_h
    port map (
            O => \N__14651\,
            I => \N__14606\
        );

    \I__2327\ : Span4Mux_v
    port map (
            O => \N__14648\,
            I => \N__14606\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__14645\,
            I => \N__14606\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__14642\,
            I => \N__14606\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__14639\,
            I => \N__14606\
        );

    \I__2323\ : Span4Mux_v
    port map (
            O => \N__14634\,
            I => \N__14597\
        );

    \I__2322\ : Span4Mux_h
    port map (
            O => \N__14631\,
            I => \N__14597\
        );

    \I__2321\ : Span4Mux_s2_v
    port map (
            O => \N__14626\,
            I => \N__14597\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__14623\,
            I => \N__14597\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__14620\,
            I => \tok.A_stk.rd_15__N_301\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__14617\,
            I => \tok.A_stk.rd_15__N_301\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__14606\,
            I => \tok.A_stk.rd_15__N_301\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__14597\,
            I => \tok.A_stk.rd_15__N_301\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__14588\,
            I => \tok.n83_adj_735_cascade_\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__14585\,
            I => \tok.n7_cascade_\
        );

    \I__2313\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14579\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__14579\,
            I => \tok.n4516\
        );

    \I__2311\ : InMux
    port map (
            O => \N__14576\,
            I => \N__14573\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__14573\,
            I => \N__14569\
        );

    \I__2309\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14566\
        );

    \I__2308\ : Span12Mux_s6_h
    port map (
            O => \N__14569\,
            I => \N__14563\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__14566\,
            I => capture_0
        );

    \I__2306\ : Odrv12
    port map (
            O => \N__14563\,
            I => capture_0
        );

    \I__2305\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14554\
        );

    \I__2304\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14551\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__14554\,
            I => \tok.n17\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__14551\,
            I => \tok.n17\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__14546\,
            I => \tok.n4_adj_654_cascade_\
        );

    \I__2300\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14491\
        );

    \I__2299\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14491\
        );

    \I__2298\ : InMux
    port map (
            O => \N__14541\,
            I => \N__14491\
        );

    \I__2297\ : InMux
    port map (
            O => \N__14540\,
            I => \N__14491\
        );

    \I__2296\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14491\
        );

    \I__2295\ : InMux
    port map (
            O => \N__14538\,
            I => \N__14491\
        );

    \I__2294\ : InMux
    port map (
            O => \N__14537\,
            I => \N__14491\
        );

    \I__2293\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14469\
        );

    \I__2292\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14469\
        );

    \I__2291\ : InMux
    port map (
            O => \N__14534\,
            I => \N__14469\
        );

    \I__2290\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14469\
        );

    \I__2289\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14469\
        );

    \I__2288\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14469\
        );

    \I__2287\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14469\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__14529\,
            I => \N__14451\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__14528\,
            I => \N__14448\
        );

    \I__2284\ : InMux
    port map (
            O => \N__14527\,
            I => \N__14431\
        );

    \I__2283\ : InMux
    port map (
            O => \N__14526\,
            I => \N__14431\
        );

    \I__2282\ : InMux
    port map (
            O => \N__14525\,
            I => \N__14431\
        );

    \I__2281\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14431\
        );

    \I__2280\ : InMux
    port map (
            O => \N__14523\,
            I => \N__14431\
        );

    \I__2279\ : InMux
    port map (
            O => \N__14522\,
            I => \N__14431\
        );

    \I__2278\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14388\
        );

    \I__2277\ : InMux
    port map (
            O => \N__14520\,
            I => \N__14388\
        );

    \I__2276\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14388\
        );

    \I__2275\ : InMux
    port map (
            O => \N__14518\,
            I => \N__14388\
        );

    \I__2274\ : InMux
    port map (
            O => \N__14517\,
            I => \N__14388\
        );

    \I__2273\ : InMux
    port map (
            O => \N__14516\,
            I => \N__14388\
        );

    \I__2272\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14388\
        );

    \I__2271\ : InMux
    port map (
            O => \N__14514\,
            I => \N__14378\
        );

    \I__2270\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14375\
        );

    \I__2269\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14360\
        );

    \I__2268\ : InMux
    port map (
            O => \N__14511\,
            I => \N__14360\
        );

    \I__2267\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14360\
        );

    \I__2266\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14360\
        );

    \I__2265\ : InMux
    port map (
            O => \N__14508\,
            I => \N__14360\
        );

    \I__2264\ : InMux
    port map (
            O => \N__14507\,
            I => \N__14360\
        );

    \I__2263\ : InMux
    port map (
            O => \N__14506\,
            I => \N__14360\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__14491\,
            I => \N__14357\
        );

    \I__2261\ : InMux
    port map (
            O => \N__14490\,
            I => \N__14342\
        );

    \I__2260\ : InMux
    port map (
            O => \N__14489\,
            I => \N__14342\
        );

    \I__2259\ : InMux
    port map (
            O => \N__14488\,
            I => \N__14342\
        );

    \I__2258\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14342\
        );

    \I__2257\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14342\
        );

    \I__2256\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14342\
        );

    \I__2255\ : InMux
    port map (
            O => \N__14484\,
            I => \N__14342\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__14469\,
            I => \N__14339\
        );

    \I__2253\ : InMux
    port map (
            O => \N__14468\,
            I => \N__14330\
        );

    \I__2252\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14315\
        );

    \I__2251\ : InMux
    port map (
            O => \N__14466\,
            I => \N__14315\
        );

    \I__2250\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14315\
        );

    \I__2249\ : InMux
    port map (
            O => \N__14464\,
            I => \N__14315\
        );

    \I__2248\ : InMux
    port map (
            O => \N__14463\,
            I => \N__14315\
        );

    \I__2247\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14315\
        );

    \I__2246\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14315\
        );

    \I__2245\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14300\
        );

    \I__2244\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14300\
        );

    \I__2243\ : InMux
    port map (
            O => \N__14458\,
            I => \N__14300\
        );

    \I__2242\ : InMux
    port map (
            O => \N__14457\,
            I => \N__14300\
        );

    \I__2241\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14300\
        );

    \I__2240\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14300\
        );

    \I__2239\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14300\
        );

    \I__2238\ : InMux
    port map (
            O => \N__14451\,
            I => \N__14295\
        );

    \I__2237\ : InMux
    port map (
            O => \N__14448\,
            I => \N__14295\
        );

    \I__2236\ : InMux
    port map (
            O => \N__14447\,
            I => \N__14286\
        );

    \I__2235\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14286\
        );

    \I__2234\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14286\
        );

    \I__2233\ : InMux
    port map (
            O => \N__14444\,
            I => \N__14286\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__14431\,
            I => \N__14283\
        );

    \I__2231\ : InMux
    port map (
            O => \N__14430\,
            I => \N__14268\
        );

    \I__2230\ : InMux
    port map (
            O => \N__14429\,
            I => \N__14268\
        );

    \I__2229\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14268\
        );

    \I__2228\ : InMux
    port map (
            O => \N__14427\,
            I => \N__14268\
        );

    \I__2227\ : InMux
    port map (
            O => \N__14426\,
            I => \N__14268\
        );

    \I__2226\ : InMux
    port map (
            O => \N__14425\,
            I => \N__14268\
        );

    \I__2225\ : InMux
    port map (
            O => \N__14424\,
            I => \N__14268\
        );

    \I__2224\ : InMux
    port map (
            O => \N__14423\,
            I => \N__14253\
        );

    \I__2223\ : InMux
    port map (
            O => \N__14422\,
            I => \N__14253\
        );

    \I__2222\ : InMux
    port map (
            O => \N__14421\,
            I => \N__14253\
        );

    \I__2221\ : InMux
    port map (
            O => \N__14420\,
            I => \N__14253\
        );

    \I__2220\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14253\
        );

    \I__2219\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14253\
        );

    \I__2218\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14253\
        );

    \I__2217\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14217\
        );

    \I__2216\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14217\
        );

    \I__2215\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14217\
        );

    \I__2214\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14217\
        );

    \I__2213\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14217\
        );

    \I__2212\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14217\
        );

    \I__2211\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14217\
        );

    \I__2210\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14202\
        );

    \I__2209\ : InMux
    port map (
            O => \N__14408\,
            I => \N__14202\
        );

    \I__2208\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14202\
        );

    \I__2207\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14202\
        );

    \I__2206\ : InMux
    port map (
            O => \N__14405\,
            I => \N__14202\
        );

    \I__2205\ : InMux
    port map (
            O => \N__14404\,
            I => \N__14202\
        );

    \I__2204\ : InMux
    port map (
            O => \N__14403\,
            I => \N__14202\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__14388\,
            I => \N__14199\
        );

    \I__2202\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14184\
        );

    \I__2201\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14184\
        );

    \I__2200\ : InMux
    port map (
            O => \N__14385\,
            I => \N__14184\
        );

    \I__2199\ : InMux
    port map (
            O => \N__14384\,
            I => \N__14184\
        );

    \I__2198\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14184\
        );

    \I__2197\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14184\
        );

    \I__2196\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14184\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__14378\,
            I => \N__14179\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__14375\,
            I => \N__14179\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__14360\,
            I => \N__14174\
        );

    \I__2192\ : Span4Mux_s2_h
    port map (
            O => \N__14357\,
            I => \N__14174\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14171\
        );

    \I__2190\ : Span4Mux_s2_h
    port map (
            O => \N__14339\,
            I => \N__14168\
        );

    \I__2189\ : InMux
    port map (
            O => \N__14338\,
            I => \N__14155\
        );

    \I__2188\ : InMux
    port map (
            O => \N__14337\,
            I => \N__14155\
        );

    \I__2187\ : InMux
    port map (
            O => \N__14336\,
            I => \N__14155\
        );

    \I__2186\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14155\
        );

    \I__2185\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14155\
        );

    \I__2184\ : InMux
    port map (
            O => \N__14333\,
            I => \N__14155\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__14330\,
            I => \N__14148\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__14315\,
            I => \N__14148\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__14300\,
            I => \N__14148\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__14295\,
            I => \N__14137\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__14286\,
            I => \N__14137\
        );

    \I__2178\ : Span4Mux_s3_v
    port map (
            O => \N__14283\,
            I => \N__14137\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__14268\,
            I => \N__14137\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__14253\,
            I => \N__14137\
        );

    \I__2175\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14119\
        );

    \I__2174\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14119\
        );

    \I__2173\ : InMux
    port map (
            O => \N__14250\,
            I => \N__14119\
        );

    \I__2172\ : InMux
    port map (
            O => \N__14249\,
            I => \N__14119\
        );

    \I__2171\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14119\
        );

    \I__2170\ : InMux
    port map (
            O => \N__14247\,
            I => \N__14119\
        );

    \I__2169\ : InMux
    port map (
            O => \N__14246\,
            I => \N__14119\
        );

    \I__2168\ : InMux
    port map (
            O => \N__14245\,
            I => \N__14104\
        );

    \I__2167\ : InMux
    port map (
            O => \N__14244\,
            I => \N__14104\
        );

    \I__2166\ : InMux
    port map (
            O => \N__14243\,
            I => \N__14104\
        );

    \I__2165\ : InMux
    port map (
            O => \N__14242\,
            I => \N__14104\
        );

    \I__2164\ : InMux
    port map (
            O => \N__14241\,
            I => \N__14104\
        );

    \I__2163\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14104\
        );

    \I__2162\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14104\
        );

    \I__2161\ : InMux
    port map (
            O => \N__14238\,
            I => \N__14089\
        );

    \I__2160\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14089\
        );

    \I__2159\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14089\
        );

    \I__2158\ : InMux
    port map (
            O => \N__14235\,
            I => \N__14089\
        );

    \I__2157\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14089\
        );

    \I__2156\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14089\
        );

    \I__2155\ : InMux
    port map (
            O => \N__14232\,
            I => \N__14089\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__14217\,
            I => \N__14082\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__14202\,
            I => \N__14082\
        );

    \I__2152\ : Span4Mux_h
    port map (
            O => \N__14199\,
            I => \N__14082\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__14184\,
            I => \N__14075\
        );

    \I__2150\ : Span4Mux_h
    port map (
            O => \N__14179\,
            I => \N__14075\
        );

    \I__2149\ : Span4Mux_h
    port map (
            O => \N__14174\,
            I => \N__14075\
        );

    \I__2148\ : Span4Mux_h
    port map (
            O => \N__14171\,
            I => \N__14070\
        );

    \I__2147\ : Span4Mux_h
    port map (
            O => \N__14168\,
            I => \N__14070\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__14155\,
            I => \N__14063\
        );

    \I__2145\ : Span4Mux_s3_h
    port map (
            O => \N__14148\,
            I => \N__14063\
        );

    \I__2144\ : Span4Mux_v
    port map (
            O => \N__14137\,
            I => \N__14063\
        );

    \I__2143\ : InMux
    port map (
            O => \N__14136\,
            I => \N__14056\
        );

    \I__2142\ : InMux
    port map (
            O => \N__14135\,
            I => \N__14056\
        );

    \I__2141\ : InMux
    port map (
            O => \N__14134\,
            I => \N__14056\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__14119\,
            I => n786
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__14104\,
            I => n786
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__14089\,
            I => n786
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__14082\,
            I => n786
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__14075\,
            I => n786
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__14070\,
            I => n786
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__14063\,
            I => n786
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__14056\,
            I => n786
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__14039\,
            I => \N__14035\
        );

    \I__2131\ : InMux
    port map (
            O => \N__14038\,
            I => \N__14030\
        );

    \I__2130\ : InMux
    port map (
            O => \N__14035\,
            I => \N__14030\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__14030\,
            I => \tok.A_stk.tail_31\
        );

    \I__2128\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14021\
        );

    \I__2127\ : InMux
    port map (
            O => \N__14026\,
            I => \N__14021\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__14021\,
            I => \tok.A_stk.tail_15\
        );

    \I__2125\ : InMux
    port map (
            O => \N__14018\,
            I => \N__14012\
        );

    \I__2124\ : InMux
    port map (
            O => \N__14017\,
            I => \N__14012\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__14012\,
            I => \tok.A_stk.tail_79\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__14009\,
            I => \N__14006\
        );

    \I__2121\ : InMux
    port map (
            O => \N__14006\,
            I => \N__14000\
        );

    \I__2120\ : InMux
    port map (
            O => \N__14005\,
            I => \N__14000\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__14000\,
            I => \tok.A_stk.tail_95\
        );

    \I__2118\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13993\
        );

    \I__2117\ : InMux
    port map (
            O => \N__13996\,
            I => \N__13990\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__13993\,
            I => tail_111
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__13990\,
            I => tail_111
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__13985\,
            I => \N__13982\
        );

    \I__2113\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13978\
        );

    \I__2112\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13975\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__13978\,
            I => \N__13972\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__13975\,
            I => \N__13969\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__13972\,
            I => tail_127
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__13969\,
            I => tail_127
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__2106\ : InMux
    port map (
            O => \N__13961\,
            I => \N__13957\
        );

    \I__2105\ : InMux
    port map (
            O => \N__13960\,
            I => \N__13954\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__13957\,
            I => tail_97
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__13954\,
            I => tail_97
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__13949\,
            I => \N__13946\
        );

    \I__2101\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13942\
        );

    \I__2100\ : InMux
    port map (
            O => \N__13945\,
            I => \N__13939\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__13942\,
            I => tail_113
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__13939\,
            I => tail_113
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__13934\,
            I => \N__13918\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__13933\,
            I => \N__13915\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__13932\,
            I => \N__13912\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__13931\,
            I => \N__13901\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__13930\,
            I => \N__13898\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__13929\,
            I => \N__13895\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__13928\,
            I => \N__13867\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__13927\,
            I => \N__13864\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__13926\,
            I => \N__13861\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__13925\,
            I => \N__13854\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__13924\,
            I => \N__13851\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__13923\,
            I => \N__13848\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__13922\,
            I => \N__13843\
        );

    \I__2084\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13821\
        );

    \I__2083\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13821\
        );

    \I__2082\ : InMux
    port map (
            O => \N__13915\,
            I => \N__13821\
        );

    \I__2081\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13821\
        );

    \I__2080\ : InMux
    port map (
            O => \N__13911\,
            I => \N__13821\
        );

    \I__2079\ : InMux
    port map (
            O => \N__13910\,
            I => \N__13821\
        );

    \I__2078\ : InMux
    port map (
            O => \N__13909\,
            I => \N__13821\
        );

    \I__2077\ : InMux
    port map (
            O => \N__13908\,
            I => \N__13818\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__13907\,
            I => \N__13810\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__13906\,
            I => \N__13807\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__13905\,
            I => \N__13804\
        );

    \I__2073\ : InMux
    port map (
            O => \N__13904\,
            I => \N__13785\
        );

    \I__2072\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13785\
        );

    \I__2071\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13785\
        );

    \I__2070\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13785\
        );

    \I__2069\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13785\
        );

    \I__2068\ : InMux
    port map (
            O => \N__13893\,
            I => \N__13785\
        );

    \I__2067\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13785\
        );

    \I__2066\ : InMux
    port map (
            O => \N__13891\,
            I => \N__13772\
        );

    \I__2065\ : InMux
    port map (
            O => \N__13890\,
            I => \N__13772\
        );

    \I__2064\ : InMux
    port map (
            O => \N__13889\,
            I => \N__13772\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__13888\,
            I => \N__13764\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__13887\,
            I => \N__13761\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__13886\,
            I => \N__13758\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__13885\,
            I => \N__13752\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__13884\,
            I => \N__13749\
        );

    \I__2058\ : InMux
    port map (
            O => \N__13883\,
            I => \N__13730\
        );

    \I__2057\ : InMux
    port map (
            O => \N__13882\,
            I => \N__13730\
        );

    \I__2056\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13730\
        );

    \I__2055\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13730\
        );

    \I__2054\ : InMux
    port map (
            O => \N__13879\,
            I => \N__13730\
        );

    \I__2053\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13730\
        );

    \I__2052\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13730\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__13876\,
            I => \N__13716\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__13875\,
            I => \N__13712\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__13874\,
            I => \N__13709\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__13873\,
            I => \N__13706\
        );

    \I__2047\ : InMux
    port map (
            O => \N__13872\,
            I => \N__13696\
        );

    \I__2046\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13696\
        );

    \I__2045\ : InMux
    port map (
            O => \N__13870\,
            I => \N__13696\
        );

    \I__2044\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13683\
        );

    \I__2043\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13683\
        );

    \I__2042\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13683\
        );

    \I__2041\ : InMux
    port map (
            O => \N__13860\,
            I => \N__13683\
        );

    \I__2040\ : InMux
    port map (
            O => \N__13859\,
            I => \N__13683\
        );

    \I__2039\ : InMux
    port map (
            O => \N__13858\,
            I => \N__13683\
        );

    \I__2038\ : InMux
    port map (
            O => \N__13857\,
            I => \N__13670\
        );

    \I__2037\ : InMux
    port map (
            O => \N__13854\,
            I => \N__13670\
        );

    \I__2036\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13670\
        );

    \I__2035\ : InMux
    port map (
            O => \N__13848\,
            I => \N__13670\
        );

    \I__2034\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13670\
        );

    \I__2033\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13670\
        );

    \I__2032\ : InMux
    port map (
            O => \N__13843\,
            I => \N__13667\
        );

    \I__2031\ : InMux
    port map (
            O => \N__13842\,
            I => \N__13660\
        );

    \I__2030\ : InMux
    port map (
            O => \N__13841\,
            I => \N__13660\
        );

    \I__2029\ : InMux
    port map (
            O => \N__13840\,
            I => \N__13660\
        );

    \I__2028\ : InMux
    port map (
            O => \N__13839\,
            I => \N__13651\
        );

    \I__2027\ : InMux
    port map (
            O => \N__13838\,
            I => \N__13651\
        );

    \I__2026\ : InMux
    port map (
            O => \N__13837\,
            I => \N__13651\
        );

    \I__2025\ : InMux
    port map (
            O => \N__13836\,
            I => \N__13651\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__13821\,
            I => \N__13646\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__13818\,
            I => \N__13646\
        );

    \I__2022\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13635\
        );

    \I__2021\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13632\
        );

    \I__2020\ : InMux
    port map (
            O => \N__13815\,
            I => \N__13619\
        );

    \I__2019\ : InMux
    port map (
            O => \N__13814\,
            I => \N__13619\
        );

    \I__2018\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13619\
        );

    \I__2017\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13619\
        );

    \I__2016\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13619\
        );

    \I__2015\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13619\
        );

    \I__2014\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13610\
        );

    \I__2013\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13610\
        );

    \I__2012\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13610\
        );

    \I__2011\ : InMux
    port map (
            O => \N__13800\,
            I => \N__13610\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__13785\,
            I => \N__13607\
        );

    \I__2009\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13594\
        );

    \I__2008\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13594\
        );

    \I__2007\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13594\
        );

    \I__2006\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13594\
        );

    \I__2005\ : InMux
    port map (
            O => \N__13780\,
            I => \N__13594\
        );

    \I__2004\ : InMux
    port map (
            O => \N__13779\,
            I => \N__13594\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__13772\,
            I => \N__13591\
        );

    \I__2002\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13582\
        );

    \I__2001\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13582\
        );

    \I__2000\ : InMux
    port map (
            O => \N__13769\,
            I => \N__13582\
        );

    \I__1999\ : InMux
    port map (
            O => \N__13768\,
            I => \N__13582\
        );

    \I__1998\ : InMux
    port map (
            O => \N__13767\,
            I => \N__13567\
        );

    \I__1997\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13567\
        );

    \I__1996\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13567\
        );

    \I__1995\ : InMux
    port map (
            O => \N__13758\,
            I => \N__13567\
        );

    \I__1994\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13567\
        );

    \I__1993\ : InMux
    port map (
            O => \N__13756\,
            I => \N__13567\
        );

    \I__1992\ : InMux
    port map (
            O => \N__13755\,
            I => \N__13567\
        );

    \I__1991\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13554\
        );

    \I__1990\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13554\
        );

    \I__1989\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13554\
        );

    \I__1988\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13554\
        );

    \I__1987\ : InMux
    port map (
            O => \N__13746\,
            I => \N__13554\
        );

    \I__1986\ : InMux
    port map (
            O => \N__13745\,
            I => \N__13554\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__13730\,
            I => \N__13551\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__13729\,
            I => \N__13548\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__13728\,
            I => \N__13545\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__13727\,
            I => \N__13542\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__13726\,
            I => \N__13539\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__13725\,
            I => \N__13533\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__13724\,
            I => \N__13530\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__13723\,
            I => \N__13527\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__13722\,
            I => \N__13520\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__13721\,
            I => \N__13517\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__13720\,
            I => \N__13514\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__13719\,
            I => \N__13508\
        );

    \I__1973\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13497\
        );

    \I__1972\ : InMux
    port map (
            O => \N__13715\,
            I => \N__13482\
        );

    \I__1971\ : InMux
    port map (
            O => \N__13712\,
            I => \N__13482\
        );

    \I__1970\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13482\
        );

    \I__1969\ : InMux
    port map (
            O => \N__13706\,
            I => \N__13482\
        );

    \I__1968\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13482\
        );

    \I__1967\ : InMux
    port map (
            O => \N__13704\,
            I => \N__13482\
        );

    \I__1966\ : InMux
    port map (
            O => \N__13703\,
            I => \N__13482\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__13696\,
            I => \N__13473\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__13683\,
            I => \N__13473\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__13670\,
            I => \N__13473\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__13667\,
            I => \N__13473\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__13660\,
            I => \N__13466\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__13651\,
            I => \N__13466\
        );

    \I__1959\ : Span4Mux_s2_h
    port map (
            O => \N__13646\,
            I => \N__13466\
        );

    \I__1958\ : InMux
    port map (
            O => \N__13645\,
            I => \N__13463\
        );

    \I__1957\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13448\
        );

    \I__1956\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13448\
        );

    \I__1955\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13448\
        );

    \I__1954\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13448\
        );

    \I__1953\ : InMux
    port map (
            O => \N__13640\,
            I => \N__13448\
        );

    \I__1952\ : InMux
    port map (
            O => \N__13639\,
            I => \N__13448\
        );

    \I__1951\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13448\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__13635\,
            I => \N__13443\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__13632\,
            I => \N__13443\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__13619\,
            I => \N__13436\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__13610\,
            I => \N__13436\
        );

    \I__1946\ : Span4Mux_s2_h
    port map (
            O => \N__13607\,
            I => \N__13436\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__13594\,
            I => \N__13433\
        );

    \I__1944\ : Span4Mux_s3_h
    port map (
            O => \N__13591\,
            I => \N__13426\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__13582\,
            I => \N__13426\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__13567\,
            I => \N__13426\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__13554\,
            I => \N__13421\
        );

    \I__1940\ : Span4Mux_s3_h
    port map (
            O => \N__13551\,
            I => \N__13421\
        );

    \I__1939\ : InMux
    port map (
            O => \N__13548\,
            I => \N__13406\
        );

    \I__1938\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13406\
        );

    \I__1937\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13406\
        );

    \I__1936\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13406\
        );

    \I__1935\ : InMux
    port map (
            O => \N__13538\,
            I => \N__13406\
        );

    \I__1934\ : InMux
    port map (
            O => \N__13537\,
            I => \N__13406\
        );

    \I__1933\ : InMux
    port map (
            O => \N__13536\,
            I => \N__13406\
        );

    \I__1932\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13393\
        );

    \I__1931\ : InMux
    port map (
            O => \N__13530\,
            I => \N__13393\
        );

    \I__1930\ : InMux
    port map (
            O => \N__13527\,
            I => \N__13393\
        );

    \I__1929\ : InMux
    port map (
            O => \N__13526\,
            I => \N__13393\
        );

    \I__1928\ : InMux
    port map (
            O => \N__13525\,
            I => \N__13393\
        );

    \I__1927\ : InMux
    port map (
            O => \N__13524\,
            I => \N__13393\
        );

    \I__1926\ : InMux
    port map (
            O => \N__13523\,
            I => \N__13378\
        );

    \I__1925\ : InMux
    port map (
            O => \N__13520\,
            I => \N__13378\
        );

    \I__1924\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13378\
        );

    \I__1923\ : InMux
    port map (
            O => \N__13514\,
            I => \N__13378\
        );

    \I__1922\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13378\
        );

    \I__1921\ : InMux
    port map (
            O => \N__13512\,
            I => \N__13378\
        );

    \I__1920\ : InMux
    port map (
            O => \N__13511\,
            I => \N__13378\
        );

    \I__1919\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13373\
        );

    \I__1918\ : InMux
    port map (
            O => \N__13507\,
            I => \N__13373\
        );

    \I__1917\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13358\
        );

    \I__1916\ : InMux
    port map (
            O => \N__13505\,
            I => \N__13358\
        );

    \I__1915\ : InMux
    port map (
            O => \N__13504\,
            I => \N__13358\
        );

    \I__1914\ : InMux
    port map (
            O => \N__13503\,
            I => \N__13358\
        );

    \I__1913\ : InMux
    port map (
            O => \N__13502\,
            I => \N__13358\
        );

    \I__1912\ : InMux
    port map (
            O => \N__13501\,
            I => \N__13358\
        );

    \I__1911\ : InMux
    port map (
            O => \N__13500\,
            I => \N__13358\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__13497\,
            I => \N__13351\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__13482\,
            I => \N__13351\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__13473\,
            I => \N__13351\
        );

    \I__1907\ : Span4Mux_h
    port map (
            O => \N__13466\,
            I => \N__13348\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__13463\,
            I => \N__13339\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__13448\,
            I => \N__13339\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__13443\,
            I => \N__13339\
        );

    \I__1903\ : Span4Mux_h
    port map (
            O => \N__13436\,
            I => \N__13339\
        );

    \I__1902\ : Span4Mux_s3_h
    port map (
            O => \N__13433\,
            I => \N__13332\
        );

    \I__1901\ : Span4Mux_v
    port map (
            O => \N__13426\,
            I => \N__13332\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__13421\,
            I => \N__13332\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__13406\,
            I => n29
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__13393\,
            I => n29
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__13378\,
            I => n29
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__13373\,
            I => n29
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__13358\,
            I => n29
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__13351\,
            I => n29
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__13348\,
            I => n29
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__13339\,
            I => n29
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__13332\,
            I => n29
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__13313\,
            I => \tok.n2_adj_685_cascade_\
        );

    \I__1889\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13307\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__13307\,
            I => \tok.n14_adj_686\
        );

    \I__1887\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13301\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__13301\,
            I => \N__13297\
        );

    \I__1885\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13294\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__13297\,
            I => sender_1
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__13294\,
            I => sender_1
        );

    \I__1882\ : IoInMux
    port map (
            O => \N__13289\,
            I => \N__13286\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__13286\,
            I => \N__13283\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__13283\,
            I => tx_c
        );

    \I__1879\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13277\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__13277\,
            I => reset_c
        );

    \I__1877\ : InMux
    port map (
            O => \N__13274\,
            I => \N__13268\
        );

    \I__1876\ : InMux
    port map (
            O => \N__13273\,
            I => \N__13268\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__13268\,
            I => \tok.A_stk.tail_63\
        );

    \I__1874\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13259\
        );

    \I__1873\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13259\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__13259\,
            I => \tok.A_stk.tail_47\
        );

    \I__1871\ : InMux
    port map (
            O => \N__13256\,
            I => \N__13253\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__13253\,
            I => \N__13250\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__13250\,
            I => \tok.n6_adj_667\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__13247\,
            I => \N__13244\
        );

    \I__1867\ : InMux
    port map (
            O => \N__13244\,
            I => \N__13241\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__13241\,
            I => \tok.n294\
        );

    \I__1865\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13235\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__13235\,
            I => \N__13232\
        );

    \I__1863\ : Span4Mux_h
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__1862\ : Span4Mux_h
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__1861\ : Sp12to4
    port map (
            O => \N__13226\,
            I => \N__13223\
        );

    \I__1860\ : Odrv12
    port map (
            O => \N__13223\,
            I => \tok.table_wr_data_3\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__13220\,
            I => \N__13217\
        );

    \I__1858\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13214\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__13214\,
            I => \tok.n298\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__13211\,
            I => \N__13208\
        );

    \I__1855\ : InMux
    port map (
            O => \N__13208\,
            I => \N__13205\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__13205\,
            I => \tok.n289\
        );

    \I__1853\ : InMux
    port map (
            O => \N__13202\,
            I => \N__13199\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__13199\,
            I => \tok.n6_adj_814\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__13196\,
            I => \tok.n34_cascade_\
        );

    \I__1850\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13190\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__13190\,
            I => \N__13187\
        );

    \I__1848\ : Span4Mux_h
    port map (
            O => \N__13187\,
            I => \N__13184\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__13184\,
            I => \tok.n13\
        );

    \I__1846\ : InMux
    port map (
            O => \N__13181\,
            I => \N__13178\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__13178\,
            I => \tok.n4656\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__13175\,
            I => \tok.n20_adj_754_cascade_\
        );

    \I__1843\ : InMux
    port map (
            O => \N__13172\,
            I => \N__13169\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__13169\,
            I => \N__13166\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__13166\,
            I => \tok.n9_adj_749\
        );

    \I__1840\ : InMux
    port map (
            O => \N__13163\,
            I => \N__13160\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__13160\,
            I => \N__13157\
        );

    \I__1838\ : Span4Mux_v
    port map (
            O => \N__13157\,
            I => \N__13154\
        );

    \I__1837\ : Span4Mux_h
    port map (
            O => \N__13154\,
            I => \N__13151\
        );

    \I__1836\ : Span4Mux_s1_h
    port map (
            O => \N__13151\,
            I => \N__13148\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__13148\,
            I => \tok.table_rd_15\
        );

    \I__1834\ : InMux
    port map (
            O => \N__13145\,
            I => \N__13142\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__13142\,
            I => \tok.n16_adj_751\
        );

    \I__1832\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13136\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__13136\,
            I => \tok.n17_adj_774\
        );

    \I__1830\ : InMux
    port map (
            O => \N__13133\,
            I => \N__13130\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__13130\,
            I => \N__13127\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__13127\,
            I => \tok.n10_adj_705\
        );

    \I__1827\ : InMux
    port map (
            O => \N__13124\,
            I => \N__13121\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__13121\,
            I => \tok.n6_adj_692\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__13118\,
            I => \tok.n13_adj_688_cascade_\
        );

    \I__1824\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13112\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__13112\,
            I => \tok.n12_adj_687\
        );

    \I__1822\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13106\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__13106\,
            I => \N__13103\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__13103\,
            I => \tok.n4674\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__13100\,
            I => \tok.n20_adj_693_cascade_\
        );

    \I__1818\ : InMux
    port map (
            O => \N__13097\,
            I => \tok.n3949\
        );

    \I__1817\ : InMux
    port map (
            O => \N__13094\,
            I => \tok.n3950\
        );

    \I__1816\ : InMux
    port map (
            O => \N__13091\,
            I => \tok.n3951\
        );

    \I__1815\ : InMux
    port map (
            O => \N__13088\,
            I => \tok.n3952\
        );

    \I__1814\ : InMux
    port map (
            O => \N__13085\,
            I => \tok.n3953\
        );

    \I__1813\ : InMux
    port map (
            O => \N__13082\,
            I => \tok.n3954\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__13079\,
            I => \tok.n2_adj_739_cascade_\
        );

    \I__1811\ : InMux
    port map (
            O => \N__13076\,
            I => \N__13073\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__13073\,
            I => \N__13070\
        );

    \I__1809\ : Span4Mux_v
    port map (
            O => \N__13070\,
            I => \N__13067\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__13067\,
            I => \tok.n6_adj_753\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__13064\,
            I => \tok.n14_adj_741_cascade_\
        );

    \I__1806\ : InMux
    port map (
            O => \N__13061\,
            I => \N__13058\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__13058\,
            I => \N__13055\
        );

    \I__1804\ : Span4Mux_h
    port map (
            O => \N__13055\,
            I => \N__13052\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__13052\,
            I => \tok.n13_adj_748\
        );

    \I__1802\ : InMux
    port map (
            O => \N__13049\,
            I => \tok.n3940\
        );

    \I__1801\ : InMux
    port map (
            O => \N__13046\,
            I => \tok.n3941\
        );

    \I__1800\ : InMux
    port map (
            O => \N__13043\,
            I => \tok.n3942\
        );

    \I__1799\ : InMux
    port map (
            O => \N__13040\,
            I => \tok.n3943\
        );

    \I__1798\ : InMux
    port map (
            O => \N__13037\,
            I => \tok.n3944\
        );

    \I__1797\ : InMux
    port map (
            O => \N__13034\,
            I => \tok.n3945\
        );

    \I__1796\ : InMux
    port map (
            O => \N__13031\,
            I => \N__13028\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__13028\,
            I => \N__13025\
        );

    \I__1794\ : Odrv12
    port map (
            O => \N__13025\,
            I => \tok.n10_adj_764\
        );

    \I__1793\ : InMux
    port map (
            O => \N__13022\,
            I => \tok.n3946\
        );

    \I__1792\ : InMux
    port map (
            O => \N__13019\,
            I => \bfn_5_9_0_\
        );

    \I__1791\ : InMux
    port map (
            O => \N__13016\,
            I => \tok.n3948\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__13013\,
            I => \N__13010\
        );

    \I__1789\ : InMux
    port map (
            O => \N__13010\,
            I => \N__13004\
        );

    \I__1788\ : InMux
    port map (
            O => \N__13009\,
            I => \N__13004\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__13004\,
            I => \tok.A_stk.tail_4\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__13001\,
            I => \N__12998\
        );

    \I__1785\ : InMux
    port map (
            O => \N__12998\,
            I => \N__12995\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__12995\,
            I => \tok.n23_adj_677\
        );

    \I__1783\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12989\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__12989\,
            I => \tok.n24\
        );

    \I__1781\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12983\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__12983\,
            I => \tok.n26_adj_805\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__12980\,
            I => \tok.n30_adj_824_cascade_\
        );

    \I__1778\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12974\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__12974\,
            I => \tok.found_slot_N_145\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__12971\,
            I => \tok.n4642_cascade_\
        );

    \I__1775\ : InMux
    port map (
            O => \N__12968\,
            I => \N__12964\
        );

    \I__1774\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12961\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__12964\,
            I => \N__12958\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__12961\,
            I => \tok.key_rd_13\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__12958\,
            I => \tok.key_rd_13\
        );

    \I__1770\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12950\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__12950\,
            I => \tok.n14_adj_804\
        );

    \I__1768\ : InMux
    port map (
            O => \N__12947\,
            I => \N__12944\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__12944\,
            I => \tok.n27_adj_734\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__12941\,
            I => \N__12937\
        );

    \I__1765\ : InMux
    port map (
            O => \N__12940\,
            I => \N__12934\
        );

    \I__1764\ : InMux
    port map (
            O => \N__12937\,
            I => \N__12931\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__12934\,
            I => \N__12926\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__12931\,
            I => \N__12926\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__12926\,
            I => \tok.key_rd_12\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__12923\,
            I => \N__12920\
        );

    \I__1759\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12916\
        );

    \I__1758\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12913\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__12916\,
            I => \N__12910\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__12913\,
            I => \N__12907\
        );

    \I__1755\ : Odrv12
    port map (
            O => \N__12910\,
            I => \tok.key_rd_10\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__12907\,
            I => \tok.key_rd_10\
        );

    \I__1753\ : InMux
    port map (
            O => \N__12902\,
            I => \N__12899\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__12899\,
            I => \tok.n21_adj_714\
        );

    \I__1751\ : InMux
    port map (
            O => \N__12896\,
            I => \N__12890\
        );

    \I__1750\ : InMux
    port map (
            O => \N__12895\,
            I => \N__12890\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__12890\,
            I => \N__12887\
        );

    \I__1748\ : Span4Mux_h
    port map (
            O => \N__12887\,
            I => \N__12884\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__12884\,
            I => \tok.key_rd_2\
        );

    \I__1746\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12878\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__12878\,
            I => \N__12874\
        );

    \I__1744\ : InMux
    port map (
            O => \N__12877\,
            I => \N__12871\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__12874\,
            I => \N__12868\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__12871\,
            I => \N__12865\
        );

    \I__1741\ : Span4Mux_h
    port map (
            O => \N__12868\,
            I => \N__12860\
        );

    \I__1740\ : Span4Mux_v
    port map (
            O => \N__12865\,
            I => \N__12860\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__12860\,
            I => \tok.key_rd_7\
        );

    \I__1738\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12854\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__12854\,
            I => \tok.n22\
        );

    \I__1736\ : InMux
    port map (
            O => \N__12851\,
            I => \bfn_5_8_0_\
        );

    \I__1735\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12842\
        );

    \I__1734\ : InMux
    port map (
            O => \N__12847\,
            I => \N__12842\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__12842\,
            I => \tok.A_stk.tail_21\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__12839\,
            I => \N__12836\
        );

    \I__1731\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12830\
        );

    \I__1730\ : InMux
    port map (
            O => \N__12835\,
            I => \N__12830\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__12830\,
            I => \tok.A_stk.tail_5\
        );

    \I__1728\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12823\
        );

    \I__1727\ : InMux
    port map (
            O => \N__12826\,
            I => \N__12820\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__12823\,
            I => \N__12817\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__12820\,
            I => tail_116
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__12817\,
            I => tail_116
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__12812\,
            I => \N__12809\
        );

    \I__1722\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12806\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__12806\,
            I => \N__12802\
        );

    \I__1720\ : InMux
    port map (
            O => \N__12805\,
            I => \N__12799\
        );

    \I__1719\ : Sp12to4
    port map (
            O => \N__12802\,
            I => \N__12796\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__12799\,
            I => tail_100
        );

    \I__1717\ : Odrv12
    port map (
            O => \N__12796\,
            I => tail_100
        );

    \I__1716\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12785\
        );

    \I__1715\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12785\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__12785\,
            I => \tok.A_stk.tail_84\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__12782\,
            I => \N__12778\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__12781\,
            I => \N__12775\
        );

    \I__1711\ : InMux
    port map (
            O => \N__12778\,
            I => \N__12770\
        );

    \I__1710\ : InMux
    port map (
            O => \N__12775\,
            I => \N__12770\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__12770\,
            I => \tok.A_stk.tail_68\
        );

    \I__1708\ : InMux
    port map (
            O => \N__12767\,
            I => \N__12761\
        );

    \I__1707\ : InMux
    port map (
            O => \N__12766\,
            I => \N__12761\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__12761\,
            I => \tok.A_stk.tail_52\
        );

    \I__1705\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12752\
        );

    \I__1704\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12752\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__12752\,
            I => \tok.A_stk.tail_36\
        );

    \I__1702\ : InMux
    port map (
            O => \N__12749\,
            I => \N__12743\
        );

    \I__1701\ : InMux
    port map (
            O => \N__12748\,
            I => \N__12743\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__12743\,
            I => \tok.A_stk.tail_20\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__12740\,
            I => \N__12736\
        );

    \I__1698\ : InMux
    port map (
            O => \N__12739\,
            I => \N__12733\
        );

    \I__1697\ : InMux
    port map (
            O => \N__12736\,
            I => \N__12730\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__12733\,
            I => tail_117
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__12730\,
            I => tail_117
        );

    \I__1694\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12721\
        );

    \I__1693\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12718\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__12721\,
            I => tail_101
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__12718\,
            I => tail_101
        );

    \I__1690\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12707\
        );

    \I__1689\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12707\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__12707\,
            I => \tok.A_stk.tail_67\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__12704\,
            I => \N__12700\
        );

    \I__1686\ : InMux
    port map (
            O => \N__12703\,
            I => \N__12697\
        );

    \I__1685\ : InMux
    port map (
            O => \N__12700\,
            I => \N__12694\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__12697\,
            I => tail_99
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__12694\,
            I => tail_99
        );

    \I__1682\ : InMux
    port map (
            O => \N__12689\,
            I => \N__12683\
        );

    \I__1681\ : InMux
    port map (
            O => \N__12688\,
            I => \N__12683\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__12683\,
            I => \tok.A_stk.tail_83\
        );

    \I__1679\ : InMux
    port map (
            O => \N__12680\,
            I => \N__12676\
        );

    \I__1678\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12673\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__12676\,
            I => \tok.A_stk.tail_35\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__12673\,
            I => \tok.A_stk.tail_35\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__12668\,
            I => \N__12664\
        );

    \I__1674\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12661\
        );

    \I__1673\ : InMux
    port map (
            O => \N__12664\,
            I => \N__12658\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__12661\,
            I => \tok.A_stk.tail_3\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__12658\,
            I => \tok.A_stk.tail_3\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__12653\,
            I => \N__12649\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__12652\,
            I => \N__12646\
        );

    \I__1668\ : InMux
    port map (
            O => \N__12649\,
            I => \N__12643\
        );

    \I__1667\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12640\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__12643\,
            I => \tok.A_stk.tail_19\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__12640\,
            I => \tok.A_stk.tail_19\
        );

    \I__1664\ : InMux
    port map (
            O => \N__12635\,
            I => \N__12631\
        );

    \I__1663\ : InMux
    port map (
            O => \N__12634\,
            I => \N__12628\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__12631\,
            I => \tok.A_stk.tail_85\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__12628\,
            I => \tok.A_stk.tail_85\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__12623\,
            I => \N__12619\
        );

    \I__1659\ : InMux
    port map (
            O => \N__12622\,
            I => \N__12616\
        );

    \I__1658\ : InMux
    port map (
            O => \N__12619\,
            I => \N__12613\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__12616\,
            I => \tok.A_stk.tail_69\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__12613\,
            I => \tok.A_stk.tail_69\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__12608\,
            I => \N__12604\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__12607\,
            I => \N__12601\
        );

    \I__1653\ : InMux
    port map (
            O => \N__12604\,
            I => \N__12596\
        );

    \I__1652\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12596\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__12596\,
            I => \tok.A_stk.tail_53\
        );

    \I__1650\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12587\
        );

    \I__1649\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12587\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__12587\,
            I => \N__12584\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__12584\,
            I => \tok.A_stk.tail_37\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__12581\,
            I => \N__12577\
        );

    \I__1645\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12572\
        );

    \I__1644\ : InMux
    port map (
            O => \N__12577\,
            I => \N__12572\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__12572\,
            I => \tok.A_stk.tail_49\
        );

    \I__1642\ : InMux
    port map (
            O => \N__12569\,
            I => \N__12563\
        );

    \I__1641\ : InMux
    port map (
            O => \N__12568\,
            I => \N__12563\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__12563\,
            I => \tok.A_stk.tail_65\
        );

    \I__1639\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12554\
        );

    \I__1638\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12554\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__12554\,
            I => \tok.A_stk.tail_81\
        );

    \I__1636\ : InMux
    port map (
            O => \N__12551\,
            I => \N__12545\
        );

    \I__1635\ : InMux
    port map (
            O => \N__12550\,
            I => \N__12545\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__12545\,
            I => \tok.A_stk.tail_1\
        );

    \I__1633\ : InMux
    port map (
            O => \N__12542\,
            I => \N__12538\
        );

    \I__1632\ : InMux
    port map (
            O => \N__12541\,
            I => \N__12535\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__12538\,
            I => tail_115
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__12535\,
            I => tail_115
        );

    \I__1629\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12524\
        );

    \I__1628\ : InMux
    port map (
            O => \N__12529\,
            I => \N__12524\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__12524\,
            I => \tok.A_stk.tail_51\
        );

    \I__1626\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12515\
        );

    \I__1625\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12515\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__12515\,
            I => \tok.A_stk.tail_92\
        );

    \I__1623\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12506\
        );

    \I__1622\ : InMux
    port map (
            O => \N__12511\,
            I => \N__12506\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__12506\,
            I => \tok.A_stk.tail_76\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__12503\,
            I => \N__12500\
        );

    \I__1619\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12496\
        );

    \I__1618\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12493\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__12496\,
            I => \N__12490\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__12493\,
            I => \tok.A_stk.tail_60\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__12490\,
            I => \tok.A_stk.tail_60\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__12485\,
            I => \N__12481\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__12484\,
            I => \N__12478\
        );

    \I__1612\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12473\
        );

    \I__1611\ : InMux
    port map (
            O => \N__12478\,
            I => \N__12473\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__12473\,
            I => \tok.A_stk.tail_44\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__12470\,
            I => \N__12466\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__12469\,
            I => \N__12463\
        );

    \I__1607\ : InMux
    port map (
            O => \N__12466\,
            I => \N__12458\
        );

    \I__1606\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12458\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__12458\,
            I => \tok.A_stk.tail_28\
        );

    \I__1604\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12451\
        );

    \I__1603\ : InMux
    port map (
            O => \N__12454\,
            I => \N__12448\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__12451\,
            I => \tok.A_stk.tail_12\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__12448\,
            I => \tok.A_stk.tail_12\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__12443\,
            I => \N__12439\
        );

    \I__1599\ : InMux
    port map (
            O => \N__12442\,
            I => \N__12434\
        );

    \I__1598\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12434\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__12434\,
            I => \tok.A_stk.tail_17\
        );

    \I__1596\ : InMux
    port map (
            O => \N__12431\,
            I => \N__12425\
        );

    \I__1595\ : InMux
    port map (
            O => \N__12430\,
            I => \N__12425\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__12425\,
            I => \tok.A_stk.tail_33\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__12422\,
            I => \N__12419\
        );

    \I__1592\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12416\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__12413\,
            I => \tok.n290\
        );

    \I__1589\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12407\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__12407\,
            I => \N__12404\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__12404\,
            I => \tok.n6_adj_701\
        );

    \I__1586\ : InMux
    port map (
            O => \N__12401\,
            I => \tok.n3921\
        );

    \I__1585\ : InMux
    port map (
            O => \N__12398\,
            I => \tok.n3922\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__12395\,
            I => \N__12392\
        );

    \I__1583\ : InMux
    port map (
            O => \N__12392\,
            I => \N__12389\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__12389\,
            I => \N__12386\
        );

    \I__1581\ : Odrv12
    port map (
            O => \N__12386\,
            I => \tok.n288\
        );

    \I__1580\ : InMux
    port map (
            O => \N__12383\,
            I => \tok.n3923\
        );

    \I__1579\ : InMux
    port map (
            O => \N__12380\,
            I => \bfn_4_13_0_\
        );

    \I__1578\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12374\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__12374\,
            I => \tok.n292\
        );

    \I__1576\ : InMux
    port map (
            O => \N__12371\,
            I => \N__12368\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__12368\,
            I => \tok.n287\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__12365\,
            I => \N__12361\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__12364\,
            I => \N__12358\
        );

    \I__1572\ : InMux
    port map (
            O => \N__12361\,
            I => \N__12355\
        );

    \I__1571\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12352\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__12355\,
            I => tail_124
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__12352\,
            I => tail_124
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__12347\,
            I => \N__12343\
        );

    \I__1567\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12340\
        );

    \I__1566\ : InMux
    port map (
            O => \N__12343\,
            I => \N__12337\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__12340\,
            I => tail_108
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__12337\,
            I => tail_108
        );

    \I__1563\ : InMux
    port map (
            O => \N__12332\,
            I => \tok.n3913\
        );

    \I__1562\ : InMux
    port map (
            O => \N__12329\,
            I => \tok.n3914\
        );

    \I__1561\ : InMux
    port map (
            O => \N__12326\,
            I => \tok.n3915\
        );

    \I__1560\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12320\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__12320\,
            I => \N__12317\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__12317\,
            I => \tok.n295\
        );

    \I__1557\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12311\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__12311\,
            I => \N__12308\
        );

    \I__1555\ : Span4Mux_h
    port map (
            O => \N__12308\,
            I => \N__12305\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__12305\,
            I => \tok.n6_adj_768\
        );

    \I__1553\ : InMux
    port map (
            O => \N__12302\,
            I => \tok.n3916\
        );

    \I__1552\ : InMux
    port map (
            O => \N__12299\,
            I => \bfn_4_12_0_\
        );

    \I__1551\ : InMux
    port map (
            O => \N__12296\,
            I => \tok.n3918\
        );

    \I__1550\ : InMux
    port map (
            O => \N__12293\,
            I => \tok.n3919\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__12290\,
            I => \N__12287\
        );

    \I__1548\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12284\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__12284\,
            I => \N__12281\
        );

    \I__1546\ : Span4Mux_v
    port map (
            O => \N__12281\,
            I => \N__12278\
        );

    \I__1545\ : Odrv4
    port map (
            O => \N__12278\,
            I => \tok.n291\
        );

    \I__1544\ : InMux
    port map (
            O => \N__12275\,
            I => \tok.n3920\
        );

    \I__1543\ : InMux
    port map (
            O => \N__12272\,
            I => \N__12263\
        );

    \I__1542\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12263\
        );

    \I__1541\ : InMux
    port map (
            O => \N__12270\,
            I => \N__12263\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__12263\,
            I => capture_7
        );

    \I__1539\ : InMux
    port map (
            O => \N__12260\,
            I => \N__12257\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__12257\,
            I => \N__12252\
        );

    \I__1537\ : InMux
    port map (
            O => \N__12256\,
            I => \N__12247\
        );

    \I__1536\ : InMux
    port map (
            O => \N__12255\,
            I => \N__12247\
        );

    \I__1535\ : Odrv12
    port map (
            O => \N__12252\,
            I => capture_6
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__12247\,
            I => capture_6
        );

    \I__1533\ : SRMux
    port map (
            O => \N__12242\,
            I => \N__12236\
        );

    \I__1532\ : SRMux
    port map (
            O => \N__12241\,
            I => \N__12233\
        );

    \I__1531\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12227\
        );

    \I__1530\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12227\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__12236\,
            I => \N__12224\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__12233\,
            I => \N__12221\
        );

    \I__1527\ : InMux
    port map (
            O => \N__12232\,
            I => \N__12218\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__12227\,
            I => \N__12215\
        );

    \I__1525\ : Span4Mux_h
    port map (
            O => \N__12224\,
            I => \N__12210\
        );

    \I__1524\ : Span4Mux_v
    port map (
            O => \N__12221\,
            I => \N__12210\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__12218\,
            I => \N__12207\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__12215\,
            I => \N__12203\
        );

    \I__1521\ : Span4Mux_s1_h
    port map (
            O => \N__12210\,
            I => \N__12198\
        );

    \I__1520\ : Span4Mux_h
    port map (
            O => \N__12207\,
            I => \N__12198\
        );

    \I__1519\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12195\
        );

    \I__1518\ : Span4Mux_h
    port map (
            O => \N__12203\,
            I => \N__12192\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__12198\,
            I => txtick
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__12195\,
            I => txtick
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__12192\,
            I => txtick
        );

    \I__1514\ : InMux
    port map (
            O => \N__12185\,
            I => \bfn_4_11_0_\
        );

    \I__1513\ : InMux
    port map (
            O => \N__12182\,
            I => \tok.n3910\
        );

    \I__1512\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12176\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__12176\,
            I => \N__12173\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__12173\,
            I => \tok.n300\
        );

    \I__1509\ : InMux
    port map (
            O => \N__12170\,
            I => \tok.n3911\
        );

    \I__1508\ : InMux
    port map (
            O => \N__12167\,
            I => \tok.n3912\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__12164\,
            I => \tok.uart.n6_cascade_\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__12161\,
            I => \n23_cascade_\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__12158\,
            I => \N__12155\
        );

    \I__1504\ : InMux
    port map (
            O => \N__12155\,
            I => \N__12144\
        );

    \I__1503\ : InMux
    port map (
            O => \N__12154\,
            I => \N__12144\
        );

    \I__1502\ : InMux
    port map (
            O => \N__12153\,
            I => \N__12144\
        );

    \I__1501\ : InMux
    port map (
            O => \N__12152\,
            I => \N__12139\
        );

    \I__1500\ : InMux
    port map (
            O => \N__12151\,
            I => \N__12139\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__12144\,
            I => \N__12136\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__12139\,
            I => \tok.uart.sentbits_0\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__12136\,
            I => \tok.uart.sentbits_0\
        );

    \I__1496\ : InMux
    port map (
            O => \N__12131\,
            I => \N__12121\
        );

    \I__1495\ : InMux
    port map (
            O => \N__12130\,
            I => \N__12121\
        );

    \I__1494\ : InMux
    port map (
            O => \N__12129\,
            I => \N__12121\
        );

    \I__1493\ : InMux
    port map (
            O => \N__12128\,
            I => \N__12118\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__12121\,
            I => \N__12115\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__12118\,
            I => \tok.uart.sentbits_1\
        );

    \I__1490\ : Odrv4
    port map (
            O => \N__12115\,
            I => \tok.uart.sentbits_1\
        );

    \I__1489\ : CEMux
    port map (
            O => \N__12110\,
            I => \N__12106\
        );

    \I__1488\ : CEMux
    port map (
            O => \N__12109\,
            I => \N__12103\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__12106\,
            I => \N__12100\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__12103\,
            I => \N__12097\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__12100\,
            I => \tok.uart.n978\
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__12097\,
            I => \tok.uart.n978\
        );

    \I__1483\ : SRMux
    port map (
            O => \N__12092\,
            I => \N__12089\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__12089\,
            I => \N__12085\
        );

    \I__1481\ : SRMux
    port map (
            O => \N__12088\,
            I => \N__12082\
        );

    \I__1480\ : Span4Mux_s3_h
    port map (
            O => \N__12085\,
            I => \N__12077\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__12082\,
            I => \N__12077\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__12077\,
            I => \tok.uart.n1083\
        );

    \I__1477\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12070\
        );

    \I__1476\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12067\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__12070\,
            I => \tok.key_rd_14\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__12067\,
            I => \tok.key_rd_14\
        );

    \I__1473\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12058\
        );

    \I__1472\ : InMux
    port map (
            O => \N__12061\,
            I => \N__12055\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__12058\,
            I => \tok.key_rd_11\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__12055\,
            I => \tok.key_rd_11\
        );

    \I__1469\ : InMux
    port map (
            O => \N__12050\,
            I => \N__12047\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__12047\,
            I => \N__12044\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__12044\,
            I => \tok.table_wr_data_11\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__12041\,
            I => \N__12038\
        );

    \I__1465\ : InMux
    port map (
            O => \N__12038\,
            I => \N__12034\
        );

    \I__1464\ : InMux
    port map (
            O => \N__12037\,
            I => \N__12031\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__12034\,
            I => \tok.key_rd_15\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__12031\,
            I => \tok.key_rd_15\
        );

    \I__1461\ : InMux
    port map (
            O => \N__12026\,
            I => \N__12022\
        );

    \I__1460\ : InMux
    port map (
            O => \N__12025\,
            I => \N__12019\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__12022\,
            I => \tok.key_rd_9\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__12019\,
            I => \tok.key_rd_9\
        );

    \I__1457\ : InMux
    port map (
            O => \N__12014\,
            I => \N__12011\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__12011\,
            I => \N__12008\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__12008\,
            I => \tok.table_wr_data_7\
        );

    \I__1454\ : InMux
    port map (
            O => \N__12005\,
            I => \N__12002\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__12002\,
            I => \N__11999\
        );

    \I__1452\ : Span4Mux_h
    port map (
            O => \N__11999\,
            I => \N__11996\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__11996\,
            I => \tok.table_wr_data_4\
        );

    \I__1450\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11990\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__11990\,
            I => \N__11987\
        );

    \I__1448\ : Span4Mux_v
    port map (
            O => \N__11987\,
            I => \N__11984\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__11984\,
            I => \tok.table_wr_data_1\
        );

    \I__1446\ : InMux
    port map (
            O => \N__11981\,
            I => \N__11978\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__11978\,
            I => \N__11975\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__11975\,
            I => \N__11972\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__11972\,
            I => \tok.n15_adj_771\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__11969\,
            I => \N__11965\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__11968\,
            I => \N__11962\
        );

    \I__1440\ : InMux
    port map (
            O => \N__11965\,
            I => \N__11957\
        );

    \I__1439\ : InMux
    port map (
            O => \N__11962\,
            I => \N__11957\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__11957\,
            I => \tok.A_stk.tail_38\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__11954\,
            I => \N__11950\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__11953\,
            I => \N__11947\
        );

    \I__1435\ : InMux
    port map (
            O => \N__11950\,
            I => \N__11942\
        );

    \I__1434\ : InMux
    port map (
            O => \N__11947\,
            I => \N__11942\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__11942\,
            I => \tok.A_stk.tail_22\
        );

    \I__1432\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11933\
        );

    \I__1431\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11933\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__11933\,
            I => \tok.A_stk.tail_6\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__11930\,
            I => \tok.n20_adj_803_cascade_\
        );

    \I__1428\ : InMux
    port map (
            O => \N__11927\,
            I => \N__11921\
        );

    \I__1427\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11921\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__11921\,
            I => \tok.key_rd_5\
        );

    \I__1425\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11912\
        );

    \I__1424\ : InMux
    port map (
            O => \N__11917\,
            I => \N__11912\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__11912\,
            I => \tok.key_rd_3\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__11909\,
            I => \N__11905\
        );

    \I__1421\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11900\
        );

    \I__1420\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11900\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__11900\,
            I => \tok.key_rd_8\
        );

    \I__1418\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11894\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__11894\,
            I => \tok.n28\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__11891\,
            I => \tok.n25_cascade_\
        );

    \I__1415\ : InMux
    port map (
            O => \N__11888\,
            I => \N__11885\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__11885\,
            I => \tok.n26\
        );

    \I__1413\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11876\
        );

    \I__1412\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11876\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__11876\,
            I => \tok.A_stk.tail_77\
        );

    \I__1410\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11867\
        );

    \I__1409\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11867\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__11867\,
            I => \tok.A_stk.tail_61\
        );

    \I__1407\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11858\
        );

    \I__1406\ : InMux
    port map (
            O => \N__11863\,
            I => \N__11858\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__11858\,
            I => \tok.A_stk.tail_45\
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__11855\,
            I => \N__11851\
        );

    \I__1403\ : InMux
    port map (
            O => \N__11854\,
            I => \N__11846\
        );

    \I__1402\ : InMux
    port map (
            O => \N__11851\,
            I => \N__11846\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__11846\,
            I => \tok.A_stk.tail_29\
        );

    \I__1400\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11839\
        );

    \I__1399\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11836\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__11839\,
            I => \tok.A_stk.tail_13\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__11836\,
            I => \tok.A_stk.tail_13\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__11831\,
            I => \N__11828\
        );

    \I__1395\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11824\
        );

    \I__1394\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11821\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__11824\,
            I => \N__11818\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__11821\,
            I => tail_118
        );

    \I__1391\ : Odrv12
    port map (
            O => \N__11818\,
            I => tail_118
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__11813\,
            I => \N__11810\
        );

    \I__1389\ : InMux
    port map (
            O => \N__11810\,
            I => \N__11806\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__11809\,
            I => \N__11803\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__11806\,
            I => \N__11800\
        );

    \I__1386\ : InMux
    port map (
            O => \N__11803\,
            I => \N__11797\
        );

    \I__1385\ : Span4Mux_h
    port map (
            O => \N__11800\,
            I => \N__11794\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__11797\,
            I => tail_102
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__11794\,
            I => tail_102
        );

    \I__1382\ : InMux
    port map (
            O => \N__11789\,
            I => \N__11783\
        );

    \I__1381\ : InMux
    port map (
            O => \N__11788\,
            I => \N__11783\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__11783\,
            I => \tok.A_stk.tail_86\
        );

    \I__1379\ : InMux
    port map (
            O => \N__11780\,
            I => \N__11774\
        );

    \I__1378\ : InMux
    port map (
            O => \N__11779\,
            I => \N__11774\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__11774\,
            I => \tok.A_stk.tail_70\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__11771\,
            I => \N__11767\
        );

    \I__1375\ : InMux
    port map (
            O => \N__11770\,
            I => \N__11762\
        );

    \I__1374\ : InMux
    port map (
            O => \N__11767\,
            I => \N__11762\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__11762\,
            I => \tok.A_stk.tail_54\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__1371\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11752\
        );

    \I__1370\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11749\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__11752\,
            I => tail_98
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__11749\,
            I => tail_98
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__11744\,
            I => \N__11740\
        );

    \I__1366\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11737\
        );

    \I__1365\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11734\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__11737\,
            I => tail_114
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__11734\,
            I => tail_114
        );

    \I__1362\ : InMux
    port map (
            O => \N__11729\,
            I => \N__11725\
        );

    \I__1361\ : InMux
    port map (
            O => \N__11728\,
            I => \N__11722\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__11725\,
            I => tail_125
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__11722\,
            I => tail_125
        );

    \I__1358\ : InMux
    port map (
            O => \N__11717\,
            I => \N__11713\
        );

    \I__1357\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11710\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__11713\,
            I => tail_109
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__11710\,
            I => tail_109
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__11705\,
            I => \N__11702\
        );

    \I__1353\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11696\
        );

    \I__1352\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11696\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__11696\,
            I => \tok.A_stk.tail_93\
        );

    \I__1350\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11687\
        );

    \I__1349\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11687\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__11687\,
            I => \tok.A_stk.tail_18\
        );

    \I__1347\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11678\
        );

    \I__1346\ : InMux
    port map (
            O => \N__11683\,
            I => \N__11678\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__11678\,
            I => \tok.A_stk.tail_34\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__11675\,
            I => \N__11671\
        );

    \I__1343\ : InMux
    port map (
            O => \N__11674\,
            I => \N__11666\
        );

    \I__1342\ : InMux
    port map (
            O => \N__11671\,
            I => \N__11666\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__11666\,
            I => \tok.A_stk.tail_50\
        );

    \I__1340\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11657\
        );

    \I__1339\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11657\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__11657\,
            I => \tok.A_stk.tail_66\
        );

    \I__1337\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11648\
        );

    \I__1336\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11648\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__11648\,
            I => \tok.A_stk.tail_82\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__11645\,
            I => \N__11642\
        );

    \I__1333\ : InMux
    port map (
            O => \N__11642\,
            I => \N__11638\
        );

    \I__1332\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11635\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__11638\,
            I => \tok.A_stk.tail_2\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__11635\,
            I => \tok.A_stk.tail_2\
        );

    \I__1329\ : InMux
    port map (
            O => \N__11630\,
            I => \N__11626\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__11629\,
            I => \N__11623\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__11626\,
            I => \N__11620\
        );

    \I__1326\ : InMux
    port map (
            O => \N__11623\,
            I => \N__11617\
        );

    \I__1325\ : Span4Mux_h
    port map (
            O => \N__11620\,
            I => \N__11614\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__11617\,
            I => tail_110
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__11614\,
            I => tail_110
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__11609\,
            I => \N__11605\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__11608\,
            I => \N__11602\
        );

    \I__1320\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11599\
        );

    \I__1319\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11596\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__11599\,
            I => \N__11593\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__11596\,
            I => \N__11590\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__11593\,
            I => tail_126
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__11590\,
            I => tail_126
        );

    \I__1314\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11582\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__11582\,
            I => \tok.n4\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__11579\,
            I => \tok.n206_cascade_\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__11576\,
            I => \tok.n204_cascade_\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__11573\,
            I => \tok.n16_adj_699_cascade_\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__11570\,
            I => \N__11567\
        );

    \I__1308\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11564\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__11564\,
            I => \tok.n4667\
        );

    \I__1306\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11556\
        );

    \I__1305\ : InMux
    port map (
            O => \N__11560\,
            I => \N__11553\
        );

    \I__1304\ : InMux
    port map (
            O => \N__11559\,
            I => \N__11550\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__11556\,
            I => \N__11547\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__11553\,
            I => capture_9
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__11550\,
            I => capture_9
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__11547\,
            I => capture_9
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__11540\,
            I => \tok.n4508_cascade_\
        );

    \I__1298\ : InMux
    port map (
            O => \N__11537\,
            I => \N__11534\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__11534\,
            I => \tok.n4680\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__11531\,
            I => \tok.n16_adj_660_cascade_\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__11528\,
            I => \tok.uart.n3994_cascade_\
        );

    \I__1294\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11522\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__11522\,
            I => \N__11518\
        );

    \I__1292\ : InMux
    port map (
            O => \N__11521\,
            I => \N__11515\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__11518\,
            I => n795
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__11515\,
            I => n795
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__11510\,
            I => \tok.uart.n4506_cascade_\
        );

    \I__1288\ : SRMux
    port map (
            O => \N__11507\,
            I => \N__11504\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__11504\,
            I => \N__11501\
        );

    \I__1286\ : Span4Mux_s2_h
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__11498\,
            I => \tok.uart.rxclkcounter_6__N_477\
        );

    \I__1284\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11492\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__11492\,
            I => \tok.uart.n4438\
        );

    \I__1282\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11483\
        );

    \I__1281\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11483\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__11483\,
            I => \tok.uart.n2\
        );

    \I__1279\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__11477\,
            I => \N__11474\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__11474\,
            I => \tok.n16_adj_769\
        );

    \I__1276\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11465\
        );

    \I__1275\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11462\
        );

    \I__1274\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11457\
        );

    \I__1273\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11457\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__11465\,
            I => \tok.uart.bytephase_1\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__11462\,
            I => \tok.uart.bytephase_1\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__11457\,
            I => \tok.uart.bytephase_1\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__11450\,
            I => \N__11444\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__11449\,
            I => \N__11441\
        );

    \I__1267\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11438\
        );

    \I__1266\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11435\
        );

    \I__1265\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11430\
        );

    \I__1264\ : InMux
    port map (
            O => \N__11441\,
            I => \N__11430\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__11438\,
            I => \tok.uart.bytephase_5\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__11435\,
            I => \tok.uart.bytephase_5\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__11430\,
            I => \tok.uart.bytephase_5\
        );

    \I__1260\ : InMux
    port map (
            O => \N__11423\,
            I => \N__11417\
        );

    \I__1259\ : InMux
    port map (
            O => \N__11422\,
            I => \N__11414\
        );

    \I__1258\ : InMux
    port map (
            O => \N__11421\,
            I => \N__11409\
        );

    \I__1257\ : InMux
    port map (
            O => \N__11420\,
            I => \N__11409\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__11417\,
            I => \tok.uart.bytephase_3\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__11414\,
            I => \tok.uart.bytephase_3\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__11409\,
            I => \tok.uart.bytephase_3\
        );

    \I__1253\ : InMux
    port map (
            O => \N__11402\,
            I => \N__11396\
        );

    \I__1252\ : InMux
    port map (
            O => \N__11401\,
            I => \N__11393\
        );

    \I__1251\ : InMux
    port map (
            O => \N__11400\,
            I => \N__11388\
        );

    \I__1250\ : InMux
    port map (
            O => \N__11399\,
            I => \N__11388\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__11396\,
            I => \tok.uart.bytephase_0\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__11393\,
            I => \tok.uart.bytephase_0\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__11388\,
            I => \tok.uart.bytephase_0\
        );

    \I__1246\ : InMux
    port map (
            O => \N__11381\,
            I => \N__11376\
        );

    \I__1245\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11373\
        );

    \I__1244\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11370\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__11376\,
            I => \tok.uart.bytephase_2\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__11373\,
            I => \tok.uart.bytephase_2\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__11370\,
            I => \tok.uart.bytephase_2\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__11363\,
            I => \tok.uart.n13_cascade_\
        );

    \I__1239\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11354\
        );

    \I__1238\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11351\
        );

    \I__1237\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11346\
        );

    \I__1236\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11346\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__11354\,
            I => \tok.uart.bytephase_4\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__11351\,
            I => \tok.uart.bytephase_4\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__11346\,
            I => \tok.uart.bytephase_4\
        );

    \I__1232\ : SRMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__11336\,
            I => \N__11332\
        );

    \I__1230\ : InMux
    port map (
            O => \N__11335\,
            I => \N__11329\
        );

    \I__1229\ : Odrv12
    port map (
            O => \N__11332\,
            I => \bytephase_5__N_510\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__11329\,
            I => \bytephase_5__N_510\
        );

    \I__1227\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11320\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__11323\,
            I => \N__11317\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__11320\,
            I => \N__11313\
        );

    \I__1224\ : InMux
    port map (
            O => \N__11317\,
            I => \N__11308\
        );

    \I__1223\ : InMux
    port map (
            O => \N__11316\,
            I => \N__11308\
        );

    \I__1222\ : Span4Mux_s3_h
    port map (
            O => \N__11313\,
            I => \N__11303\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__11308\,
            I => \N__11303\
        );

    \I__1220\ : Span4Mux_v
    port map (
            O => \N__11303\,
            I => \N__11300\
        );

    \I__1219\ : IoSpan4Mux
    port map (
            O => \N__11300\,
            I => \N__11297\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__11297\,
            I => rx_c
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__11294\,
            I => \tok.n18_adj_767_cascade_\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__11291\,
            I => \tok.n20_adj_770_cascade_\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__11288\,
            I => \tok.A_15_N_113_7_cascade_\
        );

    \I__1214\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11282\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__11282\,
            I => \tok.A_15_N_84_7\
        );

    \I__1212\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__11276\,
            I => \tok.A_15_N_113_7\
        );

    \I__1210\ : InMux
    port map (
            O => \N__11273\,
            I => \N__11267\
        );

    \I__1209\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11267\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__11267\,
            I => \tok.uart.sentbits_3\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__11264\,
            I => \N__11259\
        );

    \I__1206\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11252\
        );

    \I__1205\ : InMux
    port map (
            O => \N__11262\,
            I => \N__11252\
        );

    \I__1204\ : InMux
    port map (
            O => \N__11259\,
            I => \N__11252\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__11252\,
            I => \tok.uart.sentbits_2\
        );

    \I__1202\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11245\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__11248\,
            I => \N__11242\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__11245\,
            I => \N__11239\
        );

    \I__1199\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11236\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__11239\,
            I => tail_106
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__11236\,
            I => tail_106
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__11231\,
            I => \N__11228\
        );

    \I__1195\ : InMux
    port map (
            O => \N__11228\,
            I => \N__11222\
        );

    \I__1194\ : InMux
    port map (
            O => \N__11227\,
            I => \N__11222\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__11222\,
            I => \tok.A_stk.tail_90\
        );

    \I__1192\ : InMux
    port map (
            O => \N__11219\,
            I => \N__11213\
        );

    \I__1191\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11213\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__11213\,
            I => \tok.A_stk.tail_74\
        );

    \I__1189\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11204\
        );

    \I__1188\ : InMux
    port map (
            O => \N__11209\,
            I => \N__11204\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__11204\,
            I => \tok.A_stk.tail_58\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__11201\,
            I => \N__11197\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__11200\,
            I => \N__11194\
        );

    \I__1184\ : InMux
    port map (
            O => \N__11197\,
            I => \N__11189\
        );

    \I__1183\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11189\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__11189\,
            I => \tok.A_stk.tail_42\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__11186\,
            I => \N__11182\
        );

    \I__1180\ : InMux
    port map (
            O => \N__11185\,
            I => \N__11177\
        );

    \I__1179\ : InMux
    port map (
            O => \N__11182\,
            I => \N__11177\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__11177\,
            I => \tok.A_stk.tail_26\
        );

    \I__1177\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11168\
        );

    \I__1176\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11168\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__11168\,
            I => \tok.A_stk.tail_10\
        );

    \I__1174\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11162\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__11162\,
            I => \tok.n2_adj_763\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__11159\,
            I => \tok.n13_adj_765_cascade_\
        );

    \I__1171\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11152\
        );

    \I__1170\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11149\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__11152\,
            I => \tok.A_stk.tail_8\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__11149\,
            I => \tok.A_stk.tail_8\
        );

    \I__1167\ : InMux
    port map (
            O => \N__11144\,
            I => \N__11140\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__11143\,
            I => \N__11137\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__11140\,
            I => \N__11134\
        );

    \I__1164\ : InMux
    port map (
            O => \N__11137\,
            I => \N__11131\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__11134\,
            I => tail_96
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__11131\,
            I => tail_96
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__11126\,
            I => \N__11123\
        );

    \I__1160\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11119\
        );

    \I__1159\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11116\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__11119\,
            I => \N__11113\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__11116\,
            I => tail_112
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__11113\,
            I => tail_112
        );

    \I__1155\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__11105\,
            I => \N__11101\
        );

    \I__1153\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11098\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__11101\,
            I => tail_105
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__11098\,
            I => tail_105
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__1149\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11086\
        );

    \I__1148\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11083\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__11086\,
            I => \N__11080\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__11083\,
            I => tail_121
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__11080\,
            I => tail_121
        );

    \I__1144\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11071\
        );

    \I__1143\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11068\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__11071\,
            I => tail_104
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__11068\,
            I => tail_104
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__11063\,
            I => \N__11060\
        );

    \I__1139\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11056\
        );

    \I__1138\ : InMux
    port map (
            O => \N__11059\,
            I => \N__11053\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__11056\,
            I => \N__11050\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__11053\,
            I => tail_120
        );

    \I__1135\ : Odrv4
    port map (
            O => \N__11050\,
            I => tail_120
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__11045\,
            I => \N__11042\
        );

    \I__1133\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11039\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__11039\,
            I => \N__11035\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__11038\,
            I => \N__11032\
        );

    \I__1130\ : Span4Mux_v
    port map (
            O => \N__11035\,
            I => \N__11029\
        );

    \I__1129\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11026\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__11029\,
            I => tail_103
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__11026\,
            I => tail_103
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__11021\,
            I => \N__11018\
        );

    \I__1125\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11015\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__11015\,
            I => \N__11011\
        );

    \I__1123\ : InMux
    port map (
            O => \N__11014\,
            I => \N__11008\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__11011\,
            I => \N__11005\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__11008\,
            I => tail_119
        );

    \I__1120\ : Odrv4
    port map (
            O => \N__11005\,
            I => tail_119
        );

    \I__1119\ : InMux
    port map (
            O => \N__11000\,
            I => \N__10997\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__10997\,
            I => \N__10994\
        );

    \I__1117\ : Span4Mux_h
    port map (
            O => \N__10994\,
            I => \N__10991\
        );

    \I__1116\ : Odrv4
    port map (
            O => \N__10991\,
            I => \tok.table_wr_data_12\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__10988\,
            I => \N__10985\
        );

    \I__1114\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10981\
        );

    \I__1113\ : InMux
    port map (
            O => \N__10984\,
            I => \N__10978\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__10981\,
            I => \N__10975\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__10978\,
            I => tail_122
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__10975\,
            I => tail_122
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__10970\,
            I => \N__10966\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__10969\,
            I => \N__10963\
        );

    \I__1107\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10958\
        );

    \I__1106\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10958\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__10958\,
            I => \tok.A_stk.tail_30\
        );

    \I__1104\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10951\
        );

    \I__1103\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10948\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__10951\,
            I => \tok.A_stk.tail_14\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__10948\,
            I => \tok.A_stk.tail_14\
        );

    \I__1100\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10937\
        );

    \I__1099\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10937\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__10937\,
            I => \tok.A_stk.tail_88\
        );

    \I__1097\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10928\
        );

    \I__1096\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10928\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__10928\,
            I => \tok.A_stk.tail_72\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__10925\,
            I => \N__10921\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__10924\,
            I => \N__10918\
        );

    \I__1092\ : InMux
    port map (
            O => \N__10921\,
            I => \N__10913\
        );

    \I__1091\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10913\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__10913\,
            I => \N__10910\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__10910\,
            I => \tok.A_stk.tail_56\
        );

    \I__1088\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10901\
        );

    \I__1087\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10901\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__10901\,
            I => \tok.A_stk.tail_40\
        );

    \I__1085\ : InMux
    port map (
            O => \N__10898\,
            I => \N__10892\
        );

    \I__1084\ : InMux
    port map (
            O => \N__10897\,
            I => \N__10892\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__10892\,
            I => \tok.A_stk.tail_24\
        );

    \I__1082\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10883\
        );

    \I__1081\ : InMux
    port map (
            O => \N__10888\,
            I => \N__10883\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__10883\,
            I => \tok.A_stk.tail_64\
        );

    \I__1079\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10874\
        );

    \I__1078\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10874\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__10874\,
            I => \tok.A_stk.tail_80\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__1075\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10864\
        );

    \I__1074\ : InMux
    port map (
            O => \N__10867\,
            I => \N__10861\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__10864\,
            I => \tok.A_stk.tail_0\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__10861\,
            I => \tok.A_stk.tail_0\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__1070\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10847\
        );

    \I__1069\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10847\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__10844\,
            I => \tok.A_stk.tail_94\
        );

    \I__1066\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10835\
        );

    \I__1065\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10835\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__10835\,
            I => \tok.A_stk.tail_78\
        );

    \I__1063\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10826\
        );

    \I__1062\ : InMux
    port map (
            O => \N__10831\,
            I => \N__10826\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__10826\,
            I => \tok.A_stk.tail_62\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__10823\,
            I => \N__10819\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__10822\,
            I => \N__10816\
        );

    \I__1058\ : InMux
    port map (
            O => \N__10819\,
            I => \N__10811\
        );

    \I__1057\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10811\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__10811\,
            I => \tok.A_stk.tail_46\
        );

    \I__1055\ : InMux
    port map (
            O => \N__10808\,
            I => \tok.uart.n3963\
        );

    \I__1054\ : InMux
    port map (
            O => \N__10805\,
            I => \tok.uart.n3964\
        );

    \I__1053\ : InMux
    port map (
            O => \N__10802\,
            I => \tok.uart.n3965\
        );

    \I__1052\ : InMux
    port map (
            O => \N__10799\,
            I => \tok.uart.n3966\
        );

    \I__1051\ : InMux
    port map (
            O => \N__10796\,
            I => \tok.uart.n3967\
        );

    \I__1050\ : CEMux
    port map (
            O => \N__10793\,
            I => \N__10790\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__10790\,
            I => \N__10787\
        );

    \I__1048\ : Span4Mux_v
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__1047\ : Odrv4
    port map (
            O => \N__10784\,
            I => n940
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__1045\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10772\
        );

    \I__1044\ : InMux
    port map (
            O => \N__10777\,
            I => \N__10772\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__10772\,
            I => \tok.A_stk.tail_16\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__10769\,
            I => \N__10765\
        );

    \I__1041\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10762\
        );

    \I__1040\ : InMux
    port map (
            O => \N__10765\,
            I => \N__10759\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__10762\,
            I => \tok.A_stk.tail_32\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__10759\,
            I => \tok.A_stk.tail_32\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__10754\,
            I => \N__10750\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__10753\,
            I => \N__10747\
        );

    \I__1035\ : InMux
    port map (
            O => \N__10750\,
            I => \N__10742\
        );

    \I__1034\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10742\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__10742\,
            I => \tok.A_stk.tail_48\
        );

    \I__1032\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10736\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__10736\,
            I => \N__10733\
        );

    \I__1030\ : Odrv4
    port map (
            O => \N__10733\,
            I => \tok.table_wr_data_8\
        );

    \I__1029\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10727\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__1027\ : Span4Mux_v
    port map (
            O => \N__10724\,
            I => \N__10721\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__10721\,
            I => \tok.table_wr_data_15\
        );

    \I__1025\ : InMux
    port map (
            O => \N__10718\,
            I => \N__10715\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__10715\,
            I => \N__10712\
        );

    \I__1023\ : Span4Mux_h
    port map (
            O => \N__10712\,
            I => \N__10709\
        );

    \I__1022\ : Span4Mux_s1_h
    port map (
            O => \N__10709\,
            I => \N__10706\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__10706\,
            I => \tok.table_wr_data_14\
        );

    \I__1020\ : InMux
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__10697\,
            I => \tok.table_wr_data_13\
        );

    \I__1017\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10691\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__1015\ : Odrv4
    port map (
            O => \N__10688\,
            I => \tok.uart.n12\
        );

    \I__1014\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10681\
        );

    \I__1013\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10678\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__10681\,
            I => \tok.uart.rxclkcounter_6\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__10678\,
            I => \tok.uart.rxclkcounter_6\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__10673\,
            I => \N__10669\
        );

    \I__1009\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10666\
        );

    \I__1008\ : InMux
    port map (
            O => \N__10669\,
            I => \N__10663\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__10666\,
            I => \tok.uart.rxclkcounter_5\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__10663\,
            I => \tok.uart.rxclkcounter_5\
        );

    \I__1005\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10654\
        );

    \I__1004\ : InMux
    port map (
            O => \N__10657\,
            I => \N__10651\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__10654\,
            I => \tok.uart.rxclkcounter_2\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__10651\,
            I => \tok.uart.rxclkcounter_2\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__10646\,
            I => \n795_cascade_\
        );

    \I__1000\ : InMux
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__998\ : Span4Mux_h
    port map (
            O => \N__10637\,
            I => \N__10634\
        );

    \I__997\ : Odrv4
    port map (
            O => \N__10634\,
            I => \tok.table_wr_data_9\
        );

    \I__996\ : InMux
    port map (
            O => \N__10631\,
            I => \bfn_1_10_0_\
        );

    \I__995\ : SRMux
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__993\ : Span4Mux_h
    port map (
            O => \N__10622\,
            I => \N__10619\
        );

    \I__992\ : Span4Mux_s0_h
    port map (
            O => \N__10619\,
            I => \N__10616\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__10616\,
            I => \tok.uart.n1081\
        );

    \I__990\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10609\
        );

    \I__989\ : InMux
    port map (
            O => \N__10612\,
            I => \N__10606\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__10609\,
            I => \tok.uart.rxclkcounter_0\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__10606\,
            I => \tok.uart.rxclkcounter_0\
        );

    \I__986\ : InMux
    port map (
            O => \N__10601\,
            I => \bfn_1_8_0_\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__10598\,
            I => \N__10595\
        );

    \I__984\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10591\
        );

    \I__983\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10588\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__10591\,
            I => \N__10585\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__10588\,
            I => \tok.uart.rxclkcounter_1\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__10585\,
            I => \tok.uart.rxclkcounter_1\
        );

    \I__979\ : InMux
    port map (
            O => \N__10580\,
            I => \tok.uart.n3968\
        );

    \I__978\ : InMux
    port map (
            O => \N__10577\,
            I => \tok.uart.n3969\
        );

    \I__977\ : InMux
    port map (
            O => \N__10574\,
            I => \N__10570\
        );

    \I__976\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10567\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__10570\,
            I => \tok.uart.rxclkcounter_3\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__10567\,
            I => \tok.uart.rxclkcounter_3\
        );

    \I__973\ : InMux
    port map (
            O => \N__10562\,
            I => \tok.uart.n3970\
        );

    \I__972\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10555\
        );

    \I__971\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10552\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__10555\,
            I => \tok.uart.rxclkcounter_4\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__10552\,
            I => \tok.uart.rxclkcounter_4\
        );

    \I__968\ : InMux
    port map (
            O => \N__10547\,
            I => \tok.uart.n3971\
        );

    \I__967\ : InMux
    port map (
            O => \N__10544\,
            I => \tok.uart.n3972\
        );

    \I__966\ : InMux
    port map (
            O => \N__10541\,
            I => \tok.uart.n3973\
        );

    \I__965\ : InMux
    port map (
            O => \N__10538\,
            I => \tok.uart.n3960\
        );

    \I__964\ : InMux
    port map (
            O => \N__10535\,
            I => \tok.uart.n3961\
        );

    \I__963\ : InMux
    port map (
            O => \N__10532\,
            I => \bfn_1_6_0_\
        );

    \I__962\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10525\
        );

    \I__961\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10522\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__10525\,
            I => \N__10519\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__10522\,
            I => \tok.uart.txclkcounter_3\
        );

    \I__958\ : Odrv4
    port map (
            O => \N__10519\,
            I => \tok.uart.txclkcounter_3\
        );

    \I__957\ : InMux
    port map (
            O => \N__10514\,
            I => \N__10510\
        );

    \I__956\ : InMux
    port map (
            O => \N__10513\,
            I => \N__10507\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__10510\,
            I => \N__10504\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__10507\,
            I => \tok.uart.txclkcounter_5\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__10504\,
            I => \tok.uart.txclkcounter_5\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__10499\,
            I => \N__10496\
        );

    \I__951\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10492\
        );

    \I__950\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10489\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__10492\,
            I => \N__10486\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__10489\,
            I => \tok.uart.txclkcounter_0\
        );

    \I__947\ : Odrv12
    port map (
            O => \N__10486\,
            I => \tok.uart.txclkcounter_0\
        );

    \I__946\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10477\
        );

    \I__945\ : InMux
    port map (
            O => \N__10480\,
            I => \N__10474\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__10477\,
            I => \N__10471\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__10474\,
            I => \tok.uart.txclkcounter_2\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__10471\,
            I => \tok.uart.txclkcounter_2\
        );

    \I__941\ : InMux
    port map (
            O => \N__10466\,
            I => \N__10462\
        );

    \I__940\ : InMux
    port map (
            O => \N__10465\,
            I => \N__10459\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10456\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__10459\,
            I => \tok.uart.txclkcounter_6\
        );

    \I__937\ : Odrv4
    port map (
            O => \N__10456\,
            I => \tok.uart.txclkcounter_6\
        );

    \I__936\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10447\
        );

    \I__935\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10444\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__10447\,
            I => \N__10441\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__10444\,
            I => \tok.uart.txclkcounter_1\
        );

    \I__932\ : Odrv12
    port map (
            O => \N__10441\,
            I => \tok.uart.txclkcounter_1\
        );

    \I__931\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10432\
        );

    \I__930\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10429\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__10432\,
            I => \N__10426\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__10429\,
            I => \tok.uart.txclkcounter_7\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__10426\,
            I => \tok.uart.txclkcounter_7\
        );

    \I__926\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10417\
        );

    \I__925\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10414\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__10417\,
            I => \N__10411\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__10414\,
            I => \tok.uart.txclkcounter_8\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__10411\,
            I => \tok.uart.txclkcounter_8\
        );

    \I__921\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10402\
        );

    \I__920\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10399\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__10402\,
            I => \N__10396\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__10399\,
            I => \tok.uart.txclkcounter_4\
        );

    \I__917\ : Odrv4
    port map (
            O => \N__10396\,
            I => \tok.uart.txclkcounter_4\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__10391\,
            I => \tok.uart.n14_cascade_\
        );

    \I__915\ : InMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__10385\,
            I => \tok.uart.n15_adj_640\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__10382\,
            I => \txtick_cascade_\
        );

    \I__912\ : InMux
    port map (
            O => \N__10379\,
            I => \N__10373\
        );

    \I__911\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10373\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__10373\,
            I => \tok.A_stk.tail_43\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__10370\,
            I => \N__10366\
        );

    \I__908\ : InMux
    port map (
            O => \N__10369\,
            I => \N__10361\
        );

    \I__907\ : InMux
    port map (
            O => \N__10366\,
            I => \N__10361\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__10361\,
            I => \tok.A_stk.tail_27\
        );

    \I__905\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10354\
        );

    \I__904\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10351\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__10354\,
            I => \tok.A_stk.tail_11\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__10351\,
            I => \tok.A_stk.tail_11\
        );

    \I__901\ : InMux
    port map (
            O => \N__10346\,
            I => \bfn_1_5_0_\
        );

    \I__900\ : InMux
    port map (
            O => \N__10343\,
            I => \tok.uart.n3955\
        );

    \I__899\ : InMux
    port map (
            O => \N__10340\,
            I => \tok.uart.n3956\
        );

    \I__898\ : InMux
    port map (
            O => \N__10337\,
            I => \tok.uart.n3957\
        );

    \I__897\ : InMux
    port map (
            O => \N__10334\,
            I => \tok.uart.n3958\
        );

    \I__896\ : InMux
    port map (
            O => \N__10331\,
            I => \tok.uart.n3959\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__10328\,
            I => \N__10324\
        );

    \I__894\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10321\
        );

    \I__893\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10318\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__10321\,
            I => \tok.A_stk.tail_39\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__10318\,
            I => \tok.A_stk.tail_39\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__10313\,
            I => \N__10309\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__10312\,
            I => \N__10306\
        );

    \I__888\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10301\
        );

    \I__887\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10301\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__10301\,
            I => \tok.A_stk.tail_23\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__10298\,
            I => \N__10295\
        );

    \I__884\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10289\
        );

    \I__883\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10289\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__10289\,
            I => \tok.A_stk.tail_7\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \N__10282\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__10285\,
            I => \N__10279\
        );

    \I__879\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10276\
        );

    \I__878\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10273\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__10276\,
            I => tail_123
        );

    \I__876\ : LocalMux
    port map (
            O => \N__10273\,
            I => tail_123
        );

    \I__875\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10264\
        );

    \I__874\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10261\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__10264\,
            I => tail_107
        );

    \I__872\ : LocalMux
    port map (
            O => \N__10261\,
            I => tail_107
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__870\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10247\
        );

    \I__869\ : InMux
    port map (
            O => \N__10252\,
            I => \N__10247\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__10247\,
            I => \tok.A_stk.tail_91\
        );

    \I__867\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10238\
        );

    \I__866\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10238\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__10238\,
            I => \tok.A_stk.tail_75\
        );

    \I__864\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10229\
        );

    \I__863\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10229\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__10229\,
            I => \tok.A_stk.tail_59\
        );

    \I__861\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10220\
        );

    \I__860\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10220\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__10220\,
            I => \tok.A_stk.tail_73\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__10217\,
            I => \N__10213\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__10216\,
            I => \N__10210\
        );

    \I__856\ : InMux
    port map (
            O => \N__10213\,
            I => \N__10205\
        );

    \I__855\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10205\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__10205\,
            I => \N__10202\
        );

    \I__853\ : Odrv4
    port map (
            O => \N__10202\,
            I => \tok.A_stk.tail_57\
        );

    \I__852\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10193\
        );

    \I__851\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10193\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__10193\,
            I => \tok.A_stk.tail_41\
        );

    \I__849\ : InMux
    port map (
            O => \N__10190\,
            I => \N__10184\
        );

    \I__848\ : InMux
    port map (
            O => \N__10189\,
            I => \N__10184\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__10184\,
            I => \tok.A_stk.tail_25\
        );

    \I__846\ : InMux
    port map (
            O => \N__10181\,
            I => \N__10177\
        );

    \I__845\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10174\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__10177\,
            I => \tok.A_stk.tail_9\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__10174\,
            I => \tok.A_stk.tail_9\
        );

    \I__842\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10163\
        );

    \I__841\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10163\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__10163\,
            I => \tok.A_stk.tail_87\
        );

    \I__839\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10154\
        );

    \I__838\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10154\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__10154\,
            I => \tok.A_stk.tail_71\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__835\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10144\
        );

    \I__834\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10141\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__10144\,
            I => \tok.A_stk.tail_55\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__10141\,
            I => \tok.A_stk.tail_55\
        );

    \I__831\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10130\
        );

    \I__830\ : InMux
    port map (
            O => \N__10135\,
            I => \N__10130\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__10130\,
            I => \tok.A_stk.tail_89\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.uart.n3962\,
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n3917\,
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n3924_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n3909\,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n3947\,
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n3932\,
            carryinitout => \bfn_9_9_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \OSCInst0\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b01"
        )
    port map (
            CLKHFPU => \N__21701\,
            CLKHFEN => \N__21700\,
            CLKHF => clk
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i123_LC_0_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__10268\,
            in1 => \N__13908\,
            in2 => \N__10286\,
            in3 => \N__14468\,
            lcout => tail_123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i105_LC_0_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10135\,
            in1 => \N__13892\,
            in2 => \N__11093\,
            in3 => \N__14541\,
            lcout => tail_105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26199\,
            ce => \N__14736\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i89_LC_0_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14539\,
            in1 => \N__11104\,
            in2 => \N__13931\,
            in3 => \N__10225\,
            lcout => \tok.A_stk.tail_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26199\,
            ce => \N__14736\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i73_LC_0_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10136\,
            in1 => \N__13894\,
            in2 => \N__10216\,
            in3 => \N__14543\,
            lcout => \tok.A_stk.tail_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26199\,
            ce => \N__14736\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i57_LC_0_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14538\,
            in1 => \N__10198\,
            in2 => \N__13930\,
            in3 => \N__10226\,
            lcout => \tok.A_stk.tail_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26199\,
            ce => \N__14736\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i41_LC_0_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10189\,
            in1 => \N__13893\,
            in2 => \N__10217\,
            in3 => \N__14542\,
            lcout => \tok.A_stk.tail_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26199\,
            ce => \N__14736\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i25_LC_0_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14537\,
            in1 => \N__10181\,
            in2 => \N__13929\,
            in3 => \N__10199\,
            lcout => \tok.A_stk.tail_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26199\,
            ce => \N__14736\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i9_LC_0_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10190\,
            in1 => \N__14540\,
            in2 => \N__21145\,
            in3 => \N__13904\,
            lcout => \tok.A_stk.tail_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26199\,
            ce => \N__14736\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i9_LC_0_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10180\,
            in1 => \N__15746\,
            in2 => \_gnd_net_\,
            in3 => \N__22651\,
            lcout => \tok.S_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26199\,
            ce => \N__14736\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i103_LC_0_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13878\,
            in1 => \N__10168\,
            in2 => \N__11021\,
            in3 => \N__14534\,
            lcout => tail_103,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26203\,
            ce => \N__14728\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i87_LC_0_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14532\,
            in1 => \N__10159\,
            in2 => \N__11038\,
            in3 => \N__13883\,
            lcout => \tok.A_stk.tail_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26203\,
            ce => \N__14728\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i71_LC_0_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13880\,
            in1 => \N__10169\,
            in2 => \N__10151\,
            in3 => \N__14536\,
            lcout => \tok.A_stk.tail_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26203\,
            ce => \N__14728\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i55_LC_0_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14531\,
            in1 => \N__10160\,
            in2 => \N__10328\,
            in3 => \N__13882\,
            lcout => \tok.A_stk.tail_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26203\,
            ce => \N__14728\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i39_LC_0_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13879\,
            in1 => \N__10147\,
            in2 => \N__10312\,
            in3 => \N__14535\,
            lcout => \tok.A_stk.tail_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26203\,
            ce => \N__14728\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i23_LC_0_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14530\,
            in1 => \N__10327\,
            in2 => \N__10298\,
            in3 => \N__13881\,
            lcout => \tok.A_stk.tail_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26203\,
            ce => \N__14728\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i7_LC_0_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__13877\,
            in1 => \N__14533\,
            in2 => \N__10313\,
            in3 => \N__19636\,
            lcout => \tok.A_stk.tail_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26203\,
            ce => \N__14728\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i7_LC_0_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10294\,
            in1 => \N__15742\,
            in2 => \_gnd_net_\,
            in3 => \N__19811\,
            lcout => \tok.S_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26203\,
            ce => \N__14728\,
            sr => \_gnd_net_\
        );

    \tok.uart.i2_3_lut_LC_0_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__11521\,
            in1 => \N__11471\,
            in2 => \_gnd_net_\,
            in3 => \N__11401\,
            lcout => n4005,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i107_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10252\,
            in1 => \N__13909\,
            in2 => \N__10285\,
            in3 => \N__14465\,
            lcout => tail_107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26197\,
            ce => \N__14729\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i91_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14463\,
            in1 => \N__10267\,
            in2 => \N__13934\,
            in3 => \N__10243\,
            lcout => \tok.A_stk.tail_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26197\,
            ce => \N__14729\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i75_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10234\,
            in1 => \N__13911\,
            in2 => \N__10256\,
            in3 => \N__14467\,
            lcout => \tok.A_stk.tail_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26197\,
            ce => \N__14729\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i59_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14462\,
            in1 => \N__10378\,
            in2 => \N__13933\,
            in3 => \N__10244\,
            lcout => \tok.A_stk.tail_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26197\,
            ce => \N__14729\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i43_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10235\,
            in1 => \N__13910\,
            in2 => \N__10370\,
            in3 => \N__14466\,
            lcout => \tok.A_stk.tail_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26197\,
            ce => \N__14729\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i27_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14461\,
            in1 => \N__10358\,
            in2 => \N__13932\,
            in3 => \N__10379\,
            lcout => \tok.A_stk.tail_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26197\,
            ce => \N__14729\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i11_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10369\,
            in1 => \N__14464\,
            in2 => \N__20843\,
            in3 => \N__13921\,
            lcout => \tok.A_stk.tail_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26197\,
            ce => \N__14729\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i11_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10357\,
            in1 => \N__15744\,
            in2 => \_gnd_net_\,
            in3 => \N__21440\,
            lcout => \tok.S_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26197\,
            ce => \N__14729\,
            sr => \_gnd_net_\
        );

    \tok.uart.txclkcounter_144__i0_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10495\,
            in2 => \_gnd_net_\,
            in3 => \N__10346\,
            lcout => \tok.uart.txclkcounter_0\,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => \tok.uart.n3955\,
            clk => \N__26200\,
            ce => 'H',
            sr => \N__12241\
        );

    \tok.uart.txclkcounter_144__i1_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10450\,
            in2 => \_gnd_net_\,
            in3 => \N__10343\,
            lcout => \tok.uart.txclkcounter_1\,
            ltout => OPEN,
            carryin => \tok.uart.n3955\,
            carryout => \tok.uart.n3956\,
            clk => \N__26200\,
            ce => 'H',
            sr => \N__12241\
        );

    \tok.uart.txclkcounter_144__i2_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10480\,
            in2 => \_gnd_net_\,
            in3 => \N__10340\,
            lcout => \tok.uart.txclkcounter_2\,
            ltout => OPEN,
            carryin => \tok.uart.n3956\,
            carryout => \tok.uart.n3957\,
            clk => \N__26200\,
            ce => 'H',
            sr => \N__12241\
        );

    \tok.uart.txclkcounter_144__i3_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10528\,
            in2 => \_gnd_net_\,
            in3 => \N__10337\,
            lcout => \tok.uart.txclkcounter_3\,
            ltout => OPEN,
            carryin => \tok.uart.n3957\,
            carryout => \tok.uart.n3958\,
            clk => \N__26200\,
            ce => 'H',
            sr => \N__12241\
        );

    \tok.uart.txclkcounter_144__i4_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10405\,
            in2 => \_gnd_net_\,
            in3 => \N__10334\,
            lcout => \tok.uart.txclkcounter_4\,
            ltout => OPEN,
            carryin => \tok.uart.n3958\,
            carryout => \tok.uart.n3959\,
            clk => \N__26200\,
            ce => 'H',
            sr => \N__12241\
        );

    \tok.uart.txclkcounter_144__i5_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10513\,
            in2 => \_gnd_net_\,
            in3 => \N__10331\,
            lcout => \tok.uart.txclkcounter_5\,
            ltout => OPEN,
            carryin => \tok.uart.n3959\,
            carryout => \tok.uart.n3960\,
            clk => \N__26200\,
            ce => 'H',
            sr => \N__12241\
        );

    \tok.uart.txclkcounter_144__i6_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10465\,
            in2 => \_gnd_net_\,
            in3 => \N__10538\,
            lcout => \tok.uart.txclkcounter_6\,
            ltout => OPEN,
            carryin => \tok.uart.n3960\,
            carryout => \tok.uart.n3961\,
            clk => \N__26200\,
            ce => 'H',
            sr => \N__12241\
        );

    \tok.uart.txclkcounter_144__i7_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10435\,
            in2 => \_gnd_net_\,
            in3 => \N__10535\,
            lcout => \tok.uart.txclkcounter_7\,
            ltout => OPEN,
            carryin => \tok.uart.n3961\,
            carryout => \tok.uart.n3962\,
            clk => \N__26200\,
            ce => 'H',
            sr => \N__12241\
        );

    \tok.uart.txclkcounter_144__i8_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10420\,
            in2 => \_gnd_net_\,
            in3 => \N__10532\,
            lcout => \tok.uart.txclkcounter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26204\,
            ce => 'H',
            sr => \N__12242\
        );

    \tok.uart.i6_4_lut_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10529\,
            in1 => \N__10514\,
            in2 => \N__10499\,
            in3 => \N__10481\,
            lcout => \tok.uart.n15_adj_640\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1014_2_lut_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12206\,
            in2 => \_gnd_net_\,
            in3 => \N__16447\,
            lcout => \tok.uart.n1081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i5_3_lut_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__10466\,
            in1 => \N__10451\,
            in2 => \_gnd_net_\,
            in3 => \N__10436\,
            lcout => OPEN,
            ltout => \tok.uart.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i4705_4_lut_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10421\,
            in1 => \N__10406\,
            in2 => \N__10391\,
            in3 => \N__10388\,
            lcout => txtick,
            ltout => \txtick_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i4701_2_lut_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__16448\,
            in1 => \_gnd_net_\,
            in2 => \N__10382\,
            in3 => \_gnd_net_\,
            lcout => \tok.uart.n964\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i10_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17345\,
            in1 => \N__19648\,
            in2 => \_gnd_net_\,
            in3 => \N__11285\,
            lcout => \tok.uart.sender_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26208\,
            ce => \N__16367\,
            sr => \N__10628\
        );

    \tok.uart.i5_4_lut_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__10612\,
            in1 => \N__10558\,
            in2 => \N__10598\,
            in3 => \N__10573\,
            lcout => \tok.uart.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rxclkcounter_147__i0_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10613\,
            in2 => \_gnd_net_\,
            in3 => \N__10601\,
            lcout => \tok.uart.rxclkcounter_0\,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => \tok.uart.n3968\,
            clk => \N__26213\,
            ce => 'H',
            sr => \N__11507\
        );

    \tok.uart.rxclkcounter_147__i1_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10594\,
            in2 => \_gnd_net_\,
            in3 => \N__10580\,
            lcout => \tok.uart.rxclkcounter_1\,
            ltout => OPEN,
            carryin => \tok.uart.n3968\,
            carryout => \tok.uart.n3969\,
            clk => \N__26213\,
            ce => 'H',
            sr => \N__11507\
        );

    \tok.uart.rxclkcounter_147__i2_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10658\,
            in2 => \_gnd_net_\,
            in3 => \N__10577\,
            lcout => \tok.uart.rxclkcounter_2\,
            ltout => OPEN,
            carryin => \tok.uart.n3969\,
            carryout => \tok.uart.n3970\,
            clk => \N__26213\,
            ce => 'H',
            sr => \N__11507\
        );

    \tok.uart.rxclkcounter_147__i3_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10574\,
            in2 => \_gnd_net_\,
            in3 => \N__10562\,
            lcout => \tok.uart.rxclkcounter_3\,
            ltout => OPEN,
            carryin => \tok.uart.n3970\,
            carryout => \tok.uart.n3971\,
            clk => \N__26213\,
            ce => 'H',
            sr => \N__11507\
        );

    \tok.uart.rxclkcounter_147__i4_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10559\,
            in2 => \_gnd_net_\,
            in3 => \N__10547\,
            lcout => \tok.uart.rxclkcounter_4\,
            ltout => OPEN,
            carryin => \tok.uart.n3971\,
            carryout => \tok.uart.n3972\,
            clk => \N__26213\,
            ce => 'H',
            sr => \N__11507\
        );

    \tok.uart.rxclkcounter_147__i5_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10672\,
            in2 => \_gnd_net_\,
            in3 => \N__10544\,
            lcout => \tok.uart.rxclkcounter_5\,
            ltout => OPEN,
            carryin => \tok.uart.n3972\,
            carryout => \tok.uart.n3973\,
            clk => \N__26213\,
            ce => 'H',
            sr => \N__11507\
        );

    \tok.uart.rxclkcounter_147__i6_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10685\,
            in2 => \_gnd_net_\,
            in3 => \N__10541\,
            lcout => \tok.uart.rxclkcounter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26213\,
            ce => 'H',
            sr => \N__11507\
        );

    \tok.i2577_2_lut_3_lut_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__23899\,
            in1 => \_gnd_net_\,
            in2 => \N__29327\,
            in3 => \N__19553\,
            lcout => \tok.table_wr_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2570_2_lut_3_lut_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20402\,
            in1 => \N__29317\,
            in2 => \_gnd_net_\,
            in3 => \N__23895\,
            lcout => \tok.table_wr_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2571_2_lut_3_lut_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__23896\,
            in1 => \_gnd_net_\,
            in2 => \N__29326\,
            in3 => \N__20507\,
            lcout => \tok.table_wr_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2572_2_lut_3_lut_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20596\,
            in1 => \N__29321\,
            in2 => \_gnd_net_\,
            in3 => \N__23897\,
            lcout => \tok.table_wr_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i6_4_lut_adj_28_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__10694\,
            in1 => \N__10684\,
            in2 => \N__10673\,
            in3 => \N__10657\,
            lcout => n795,
            ltout => \n795_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10646\,
            in3 => \N__11335\,
            lcout => n940,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i8_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14914\,
            in1 => \N__11560\,
            in2 => \_gnd_net_\,
            in3 => \N__16922\,
            lcout => capture_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2576_2_lut_3_lut_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__21158\,
            in1 => \N__29322\,
            in2 => \_gnd_net_\,
            in3 => \N__23898\,
            lcout => \tok.table_wr_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.bytephase__i0_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11402\,
            in2 => \_gnd_net_\,
            in3 => \N__10631\,
            lcout => \tok.uart.bytephase_0\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \tok.uart.n3963\,
            clk => \N__26227\,
            ce => \N__10793\,
            sr => \N__11339\
        );

    \tok.uart.bytephase__i1_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11470\,
            in2 => \_gnd_net_\,
            in3 => \N__10808\,
            lcout => \tok.uart.bytephase_1\,
            ltout => OPEN,
            carryin => \tok.uart.n3963\,
            carryout => \tok.uart.n3964\,
            clk => \N__26227\,
            ce => \N__10793\,
            sr => \N__11339\
        );

    \tok.uart.bytephase__i2_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11381\,
            in2 => \_gnd_net_\,
            in3 => \N__10805\,
            lcout => \tok.uart.bytephase_2\,
            ltout => OPEN,
            carryin => \tok.uart.n3964\,
            carryout => \tok.uart.n3965\,
            clk => \N__26227\,
            ce => \N__10793\,
            sr => \N__11339\
        );

    \tok.uart.bytephase__i3_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11423\,
            in2 => \_gnd_net_\,
            in3 => \N__10802\,
            lcout => \tok.uart.bytephase_3\,
            ltout => OPEN,
            carryin => \tok.uart.n3965\,
            carryout => \tok.uart.n3966\,
            clk => \N__26227\,
            ce => \N__10793\,
            sr => \N__11339\
        );

    \tok.uart.bytephase__i4_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11360\,
            in2 => \_gnd_net_\,
            in3 => \N__10799\,
            lcout => \tok.uart.bytephase_4\,
            ltout => OPEN,
            carryin => \tok.uart.n3966\,
            carryout => \tok.uart.n3967\,
            clk => \N__26227\,
            ce => \N__10793\,
            sr => \N__11339\
        );

    \tok.uart.bytephase__i5_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11448\,
            in2 => \_gnd_net_\,
            in3 => \N__10796\,
            lcout => \tok.uart.bytephase_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26227\,
            ce => \N__10793\,
            sr => \N__11339\
        );

    \tok.A_stk.tail_i0_i16_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10768\,
            in1 => \N__13816\,
            in2 => \N__10871\,
            in3 => \N__14514\,
            lcout => \tok.A_stk.tail_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26196\,
            ce => \N__14726\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i0_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__13779\,
            in1 => \N__14525\,
            in2 => \N__10781\,
            in3 => \N__29518\,
            lcout => \tok.A_stk.tail_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26198\,
            ce => \N__14707\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i32_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14522\,
            in1 => \N__10777\,
            in2 => \N__10754\,
            in3 => \N__13782\,
            lcout => \tok.A_stk.tail_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26198\,
            ce => \N__14707\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i48_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13780\,
            in1 => \N__10889\,
            in2 => \N__10769\,
            in3 => \N__14526\,
            lcout => \tok.A_stk.tail_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26198\,
            ce => \N__14707\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i64_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14523\,
            in1 => \N__10880\,
            in2 => \N__10753\,
            in3 => \N__13783\,
            lcout => \tok.A_stk.tail_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26198\,
            ce => \N__14707\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i80_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13781\,
            in1 => \N__10888\,
            in2 => \N__11143\,
            in3 => \N__14527\,
            lcout => \tok.A_stk.tail_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26198\,
            ce => \N__14707\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i96_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14524\,
            in1 => \N__10879\,
            in2 => \N__11126\,
            in3 => \N__13784\,
            lcout => tail_96,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26198\,
            ce => \N__14707\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i0_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10867\,
            in1 => \N__15741\,
            in2 => \_gnd_net_\,
            in3 => \N__26942\,
            lcout => \tok.S_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26198\,
            ce => \N__14707\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i110_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10852\,
            in1 => \N__13840\,
            in2 => \N__11608\,
            in3 => \N__14458\,
            lcout => tail_110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__14713\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i94_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14456\,
            in1 => \N__10840\,
            in2 => \N__11629\,
            in3 => \N__13839\,
            lcout => \tok.A_stk.tail_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__14713\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i78_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10831\,
            in1 => \N__13842\,
            in2 => \N__10856\,
            in3 => \N__14460\,
            lcout => \tok.A_stk.tail_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__14713\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i62_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14455\,
            in1 => \N__10841\,
            in2 => \N__10822\,
            in3 => \N__13838\,
            lcout => \tok.A_stk.tail_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__14713\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i46_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10832\,
            in1 => \N__13841\,
            in2 => \N__10969\,
            in3 => \N__14459\,
            lcout => \tok.A_stk.tail_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__14713\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i30_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14454\,
            in1 => \N__10955\,
            in2 => \N__10823\,
            in3 => \N__13837\,
            lcout => \tok.A_stk.tail_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__14713\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i14_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__13836\,
            in1 => \N__14457\,
            in2 => \N__10970\,
            in3 => \N__20456\,
            lcout => \tok.A_stk.tail_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__14713\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i14_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10954\,
            in1 => \N__15743\,
            in2 => \_gnd_net_\,
            in3 => \N__24003\,
            lcout => \tok.S_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__14713\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i104_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10942\,
            in1 => \N__13755\,
            in2 => \N__11063\,
            in3 => \N__14428\,
            lcout => tail_104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => \N__14737\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i88_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14426\,
            in1 => \N__11074\,
            in2 => \N__13888\,
            in3 => \N__10933\,
            lcout => \tok.A_stk.tail_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => \N__14737\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i72_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10943\,
            in1 => \N__13757\,
            in2 => \N__10924\,
            in3 => \N__14430\,
            lcout => \tok.A_stk.tail_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => \N__14737\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i56_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14425\,
            in1 => \N__10906\,
            in2 => \N__13887\,
            in3 => \N__10934\,
            lcout => \tok.A_stk.tail_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => \N__14737\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i40_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10897\,
            in1 => \N__13756\,
            in2 => \N__10925\,
            in3 => \N__14429\,
            lcout => \tok.A_stk.tail_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => \N__14737\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i24_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14424\,
            in1 => \N__10907\,
            in2 => \N__13886\,
            in3 => \N__11156\,
            lcout => \tok.A_stk.tail_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => \N__14737\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i8_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10898\,
            in1 => \N__14427\,
            in2 => \N__19554\,
            in3 => \N__13767\,
            lcout => \tok.A_stk.tail_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => \N__14737\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i8_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11155\,
            in1 => \N__15719\,
            in2 => \_gnd_net_\,
            in3 => \N__24854\,
            lcout => \tok.S_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => \N__14737\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i112_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__11122\,
            in1 => \N__13745\,
            in2 => \N__14528\,
            in3 => \N__11144\,
            lcout => tail_112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i122_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__14445\,
            in1 => \N__11249\,
            in2 => \N__13885\,
            in3 => \N__10984\,
            lcout => tail_122,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i121_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__11089\,
            in1 => \N__13748\,
            in2 => \N__14529\,
            in3 => \N__11108\,
            lcout => tail_121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i120_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__14444\,
            in1 => \N__11075\,
            in2 => \N__13884\,
            in3 => \N__11059\,
            lcout => tail_120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i119_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__11014\,
            in1 => \N__13747\,
            in2 => \N__11045\,
            in3 => \N__14447\,
            lcout => tail_119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2573_2_lut_3_lut_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20752\,
            in1 => \N__29304\,
            in2 => \_gnd_net_\,
            in3 => \N__23900\,
            lcout => \tok.table_wr_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i118_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__11827\,
            in1 => \N__13746\,
            in2 => \N__11813\,
            in3 => \N__14446\,
            lcout => tail_118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i106_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__11227\,
            in1 => \N__13768\,
            in2 => \N__10988\,
            in3 => \N__14421\,
            lcout => tail_106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26214\,
            ce => \N__14738\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i90_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14419\,
            in1 => \N__11218\,
            in2 => \N__11248\,
            in3 => \N__13891\,
            lcout => \tok.A_stk.tail_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26214\,
            ce => \N__14738\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i74_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__11209\,
            in1 => \N__13770\,
            in2 => \N__11231\,
            in3 => \N__14423\,
            lcout => \tok.A_stk.tail_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26214\,
            ce => \N__14738\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i58_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14418\,
            in1 => \N__11219\,
            in2 => \N__11200\,
            in3 => \N__13890\,
            lcout => \tok.A_stk.tail_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26214\,
            ce => \N__14738\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i42_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11210\,
            in1 => \N__13769\,
            in2 => \N__11186\,
            in3 => \N__14422\,
            lcout => \tok.A_stk.tail_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26214\,
            ce => \N__14738\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i26_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14417\,
            in1 => \N__11174\,
            in2 => \N__11201\,
            in3 => \N__13889\,
            lcout => \tok.A_stk.tail_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26214\,
            ce => \N__14738\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i10_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11185\,
            in1 => \N__14420\,
            in2 => \N__20948\,
            in3 => \N__13771\,
            lcout => \tok.A_stk.tail_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26214\,
            ce => \N__14738\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i10_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21068\,
            in1 => \N__11173\,
            in2 => \_gnd_net_\,
            in3 => \N__15745\,
            lcout => \tok.S_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26214\,
            ce => \N__14738\,
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_7_i2_2_lut_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21719\,
            in2 => \_gnd_net_\,
            in3 => \N__24495\,
            lcout => \tok.n2_adj_763\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_107_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111111011"
        )
    port map (
            in0 => \N__13031\,
            in1 => \N__26615\,
            in2 => \N__19790\,
            in3 => \N__17923\,
            lcout => OPEN,
            ltout => \tok.n13_adj_765_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_109_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__19673\,
            in1 => \N__11165\,
            in2 => \N__11159\,
            in3 => \N__29465\,
            lcout => OPEN,
            ltout => \tok.n18_adj_767_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_111_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__24074\,
            in1 => \N__14783\,
            in2 => \N__11294\,
            in3 => \N__20313\,
            lcout => OPEN,
            ltout => \tok.n20_adj_770_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_114_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__11480\,
            in1 => \N__17489\,
            in2 => \N__11291\,
            in3 => \N__11981\,
            lcout => \tok.A_15_N_113_7\,
            ltout => \tok.A_15_N_113_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A__15__I_16_i8_3_lut_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__19761\,
            in1 => \_gnd_net_\,
            in2 => \N__11288\,
            in3 => \N__17750\,
            lcout => \tok.A_15_N_84_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i8_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19674\,
            in1 => \N__17390\,
            in2 => \_gnd_net_\,
            in3 => \N__11279\,
            lcout => \tok.A_low_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26220\,
            ce => \N__17279\,
            sr => \N__19144\
        );

    \tok.i2_4_lut_adj_94_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__19757\,
            in1 => \N__20312\,
            in2 => \N__27074\,
            in3 => \N__17924\,
            lcout => \tok.n13_adj_748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i2_4_lut_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__11272\,
            in1 => \N__12153\,
            in2 => \N__11264\,
            in3 => \N__12129\,
            lcout => \tok.uart_tx_busy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sentbits_146__i3_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12131\,
            in1 => \N__11263\,
            in2 => \N__12158\,
            in3 => \N__11273\,
            lcout => \tok.uart.sentbits_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26228\,
            ce => \N__12110\,
            sr => \N__12092\
        );

    \tok.uart.sentbits_146__i2_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__11262\,
            in1 => \N__12154\,
            in2 => \_gnd_net_\,
            in3 => \N__12130\,
            lcout => \tok.uart.sentbits_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26228\,
            ce => \N__12110\,
            sr => \N__12092\
        );

    \tok.uart.i3_4_lut_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11357\,
            in1 => \N__11488\,
            in2 => \N__11449\,
            in3 => \N__11420\,
            lcout => OPEN,
            ltout => \tok.uart.n3994_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_3_lut_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14576\,
            in2 => \N__11528\,
            in3 => \N__11561\,
            lcout => \rx_data_7__N_511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i4355_2_lut_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11358\,
            in1 => \_gnd_net_\,
            in2 => \N__11450\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \tok.uart.n4506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rxrst_I_0_4_lut_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110011"
        )
    port map (
            in0 => \N__11489\,
            in1 => \N__11525\,
            in2 => \N__11510\,
            in3 => \N__11495\,
            lcout => \tok.uart.rxclkcounter_6__N_477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_adj_29_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__11324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11421\,
            lcout => \tok.uart.n4438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i2_2_lut_3_lut_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__11468\,
            in1 => \N__11399\,
            in2 => \_gnd_net_\,
            in3 => \N__11379\,
            lcout => \tok.uart.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_adj_110_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__16597\,
            in1 => \N__12314\,
            in2 => \_gnd_net_\,
            in3 => \N__27232\,
            lcout => \tok.n16_adj_769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i24_4_lut_4_lut_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100000"
        )
    port map (
            in0 => \N__11469\,
            in1 => \N__11447\,
            in2 => \N__11323\,
            in3 => \N__11422\,
            lcout => OPEN,
            ltout => \tok.uart.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_3_lut_4_lut_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11400\,
            in1 => \N__11380\,
            in2 => \N__11363\,
            in3 => \N__11359\,
            lcout => \bytephase_5__N_510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i9_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11316\,
            in1 => \N__11559\,
            in2 => \_gnd_net_\,
            in3 => \N__16928\,
            lcout => capture_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i4_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22138\,
            in1 => \N__21207\,
            in2 => \_gnd_net_\,
            in3 => \N__16926\,
            lcout => capture_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i5_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16927\,
            in1 => \N__12260\,
            in2 => \_gnd_net_\,
            in3 => \N__22137\,
            lcout => capture_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4607_4_lut_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__14987\,
            in1 => \N__21173\,
            in2 => \N__21089\,
            in3 => \N__29458\,
            lcout => \tok.n4680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_3_lut_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22589\,
            in1 => \N__26617\,
            in2 => \_gnd_net_\,
            in3 => \N__17922\,
            lcout => OPEN,
            ltout => \tok.n4508_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_41_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__13193\,
            in1 => \N__17516\,
            in2 => \N__11540\,
            in3 => \N__11585\,
            lcout => OPEN,
            ltout => \tok.n16_adj_660_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i10_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__17380\,
            in1 => \N__11537\,
            in2 => \N__11531\,
            in3 => \N__21181\,
            lcout => \tok.n59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26239\,
            ce => \N__17275\,
            sr => \N__19135\
        );

    \tok.A_i13_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001110101010"
        )
    port map (
            in0 => \N__20753\,
            in1 => \N__17518\,
            in2 => \N__11570\,
            in3 => \N__17381\,
            lcout => \tok.n56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26239\,
            ce => \N__17275\,
            sr => \N__19135\
        );

    \tok.A_i15_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110001011100"
        )
    port map (
            in0 => \N__17517\,
            in1 => \N__20495\,
            in2 => \N__17389\,
            in3 => \N__15356\,
            lcout => \tok.n54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26239\,
            ce => \N__17275\,
            sr => \N__19135\
        );

    \tok.i1_4_lut_adj_77_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100000101"
        )
    port map (
            in0 => \N__26616\,
            in1 => \N__22588\,
            in2 => \N__23982\,
            in3 => \N__24736\,
            lcout => \tok.n12_adj_723\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24737\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27445\,
            lcout => \tok.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i15_1_lut_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23952\,
            lcout => \tok.n288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_101_i11_2_lut_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22719\,
            in2 => \_gnd_net_\,
            in3 => \N__28271\,
            lcout => OPEN,
            ltout => \tok.n206_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_49_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101010000"
        )
    port map (
            in0 => \N__24497\,
            in1 => \N__29459\,
            in2 => \N__11579\,
            in3 => \N__20958\,
            lcout => \tok.n16_adj_673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i13_1_lut_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22932\,
            lcout => \tok.n290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_101_i13_2_lut_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__22718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24846\,
            lcout => OPEN,
            ltout => \tok.n204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_63_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__29460\,
            in1 => \N__20751\,
            in2 => \N__11576\,
            in3 => \N__24496\,
            lcout => OPEN,
            ltout => \tok.n16_adj_699_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4676_4_lut_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__22907\,
            in1 => \N__12410\,
            in2 => \N__11573\,
            in3 => \N__17828\,
            lcout => \tok.n4667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i124_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__12346\,
            in1 => \N__13817\,
            in2 => \N__12365\,
            in3 => \N__14513\,
            lcout => tail_124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i18_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11684\,
            in1 => \N__13703\,
            in2 => \N__11645\,
            in3 => \N__14488\,
            lcout => \tok.A_stk.tail_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26206\,
            ce => \N__14703\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i34_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14484\,
            in1 => \N__11692\,
            in2 => \N__13873\,
            in3 => \N__11674\,
            lcout => \tok.A_stk.tail_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26206\,
            ce => \N__14703\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i2_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11693\,
            in1 => \N__14487\,
            in2 => \N__20028\,
            in3 => \N__13715\,
            lcout => \tok.A_stk.tail_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26206\,
            ce => \N__14703\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i50_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14485\,
            in1 => \N__11683\,
            in2 => \N__13874\,
            in3 => \N__11663\,
            lcout => \tok.A_stk.tail_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26206\,
            ce => \N__14703\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i66_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11654\,
            in1 => \N__13704\,
            in2 => \N__11675\,
            in3 => \N__14489\,
            lcout => \tok.A_stk.tail_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26206\,
            ce => \N__14703\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i82_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14486\,
            in1 => \N__11755\,
            in2 => \N__13875\,
            in3 => \N__11662\,
            lcout => \tok.A_stk.tail_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26206\,
            ce => \N__14703\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i98_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__11653\,
            in1 => \N__13705\,
            in2 => \N__11744\,
            in3 => \N__14490\,
            lcout => tail_98,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26206\,
            ce => \N__14703\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i2_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11641\,
            in1 => \N__15720\,
            in2 => \_gnd_net_\,
            in3 => \N__21987\,
            lcout => \tok.S_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26206\,
            ce => \N__14703\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i126_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__11630\,
            in1 => \N__13860\,
            in2 => \N__11609\,
            in3 => \N__14338\,
            lcout => tail_126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i125_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__14335\,
            in1 => \N__11717\,
            in2 => \N__13928\,
            in3 => \N__11729\,
            lcout => tail_125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i117_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__14334\,
            in1 => \N__12725\,
            in2 => \N__13927\,
            in3 => \N__12739\,
            lcout => tail_117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i116_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__12826\,
            in1 => \N__13859\,
            in2 => \N__12812\,
            in3 => \N__14337\,
            lcout => tail_116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i2_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16708\,
            in1 => \N__22121\,
            in2 => \_gnd_net_\,
            in3 => \N__17200\,
            lcout => uart_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i114_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__11743\,
            in1 => \N__13858\,
            in2 => \N__11759\,
            in3 => \N__14336\,
            lcout => tail_114,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i115_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__14333\,
            in1 => \N__12703\,
            in2 => \N__13926\,
            in3 => \N__12542\,
            lcout => tail_115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i109_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__11701\,
            in1 => \N__11728\,
            in2 => \N__13922\,
            in3 => \N__14519\,
            lcout => tail_109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26215\,
            ce => \N__14727\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i93_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14517\,
            in1 => \N__11716\,
            in2 => \N__13925\,
            in3 => \N__11881\,
            lcout => \tok.A_stk.tail_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26215\,
            ce => \N__14727\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i77_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__11872\,
            in1 => \N__13847\,
            in2 => \N__11705\,
            in3 => \N__14521\,
            lcout => \tok.A_stk.tail_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26215\,
            ce => \N__14727\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i61_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14516\,
            in1 => \N__11863\,
            in2 => \N__13924\,
            in3 => \N__11882\,
            lcout => \tok.A_stk.tail_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26215\,
            ce => \N__14727\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i45_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11873\,
            in1 => \N__13846\,
            in2 => \N__11855\,
            in3 => \N__14520\,
            lcout => \tok.A_stk.tail_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26215\,
            ce => \N__14727\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i29_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14515\,
            in1 => \N__11843\,
            in2 => \N__13923\,
            in3 => \N__11864\,
            lcout => \tok.A_stk.tail_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26215\,
            ce => \N__14727\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i13_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11854\,
            in1 => \N__14518\,
            in2 => \N__20564\,
            in3 => \N__13857\,
            lcout => \tok.A_stk.tail_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26215\,
            ce => \N__14727\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i13_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11842\,
            in1 => \N__15682\,
            in2 => \_gnd_net_\,
            in3 => \N__20680\,
            lcout => \tok.S_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26215\,
            ce => \N__14727\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i102_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__11788\,
            in1 => \N__13801\,
            in2 => \N__11831\,
            in3 => \N__14510\,
            lcout => tail_102,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26223\,
            ce => \N__14708\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i86_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14508\,
            in1 => \N__11779\,
            in2 => \N__11809\,
            in3 => \N__13872\,
            lcout => \tok.A_stk.tail_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26223\,
            ce => \N__14708\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i70_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11789\,
            in1 => \N__13803\,
            in2 => \N__11771\,
            in3 => \N__14512\,
            lcout => \tok.A_stk.tail_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26223\,
            ce => \N__14708\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i54_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14507\,
            in1 => \N__11780\,
            in2 => \N__11968\,
            in3 => \N__13871\,
            lcout => \tok.A_stk.tail_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26223\,
            ce => \N__14708\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i38_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11770\,
            in1 => \N__13802\,
            in2 => \N__11953\,
            in3 => \N__14511\,
            lcout => \tok.A_stk.tail_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26223\,
            ce => \N__14708\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i22_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14506\,
            in1 => \N__11939\,
            in2 => \N__11969\,
            in3 => \N__13870\,
            lcout => \tok.A_stk.tail_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26223\,
            ce => \N__14708\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i6_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__21269\,
            in1 => \N__14509\,
            in2 => \N__11954\,
            in3 => \N__13800\,
            lcout => \tok.A_stk.tail_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26223\,
            ce => \N__14708\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i6_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15732\,
            in1 => \N__11938\,
            in2 => \_gnd_net_\,
            in3 => \N__28255\,
            lcout => \tok.S_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26223\,
            ce => \N__14708\,
            sr => \_gnd_net_\
        );

    \tok.i12_4_lut_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12026\,
            in1 => \N__12074\,
            in2 => \N__12041\,
            in3 => \N__12062\,
            lcout => \tok.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_198_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__11926\,
            in1 => \N__11917\,
            in2 => \N__22403\,
            in3 => \N__21840\,
            lcout => OPEN,
            ltout => \tok.n20_adj_803_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_136_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__24835\,
            in1 => \N__11908\,
            in2 => \N__11930\,
            in3 => \N__12953\,
            lcout => \tok.n26_adj_805\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_80_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__11927\,
            in1 => \N__11918\,
            in2 => \N__11909\,
            in3 => \N__12967\,
            lcout => \tok.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_86_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15094\,
            in1 => \N__15043\,
            in2 => \N__15121\,
            in3 => \N__15067\,
            lcout => OPEN,
            ltout => \tok.n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i15_4_lut_adj_178_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12947\,
            in1 => \N__11897\,
            in2 => \N__11891\,
            in3 => \N__11888\,
            lcout => \tok.found_slot_N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_51_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__12073\,
            in1 => \N__12061\,
            in2 => \N__24009\,
            in3 => \N__21429\,
            lcout => \tok.n23_adj_677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i12_1_lut_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2574_2_lut_3_lut_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20842\,
            in1 => \N__29265\,
            in2 => \_gnd_net_\,
            in3 => \N__23878\,
            lcout => \tok.table_wr_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_4_lut_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__12037\,
            in1 => \N__12025\,
            in2 => \N__20311\,
            in3 => \N__22636\,
            lcout => \tok.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1512_3_lut_4_lut_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__18890\,
            in1 => \N__29260\,
            in2 => \N__19691\,
            in3 => \N__23875\,
            lcout => \tok.table_wr_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i8_1_lut_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19774\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1623_3_lut_4_lut_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__24375\,
            in1 => \N__29261\,
            in2 => \N__25307\,
            in3 => \N__23876\,
            lcout => \tok.table_wr_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1734_3_lut_4_lut_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__23877\,
            in1 => \N__18650\,
            in2 => \N__29291\,
            in3 => \N__20154\,
            lcout => \tok.table_wr_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_112_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111000"
        )
    port map (
            in0 => \N__21977\,
            in1 => \N__24726\,
            in2 => \N__19592\,
            in3 => \N__28834\,
            lcout => \tok.n15_adj_771\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i3_1_lut_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21976\,
            lcout => \tok.n300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i4707_2_lut_3_lut_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__19344\,
            in1 => \N__12239\,
            in2 => \_gnd_net_\,
            in3 => \N__16423\,
            lcout => \tok.uart.n1083\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__28835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16079\,
            lcout => OPEN,
            ltout => \tok.uart.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i4698_4_lut_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19343\,
            in1 => \N__28014\,
            in2 => \N__12164\,
            in3 => \N__30441\,
            lcout => n23,
            ltout => \n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_3_lut_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__12240\,
            in1 => \_gnd_net_\,
            in2 => \N__12161\,
            in3 => \N__19345\,
            lcout => \tok.uart.n978\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sentbits_146__i0_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12151\,
            lcout => \tok.uart.sentbits_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26240\,
            ce => \N__12109\,
            sr => \N__12088\
        );

    \tok.uart.sentbits_146__i1_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12128\,
            lcout => \tok.uart.sentbits_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26240\,
            ce => \N__12109\,
            sr => \N__12088\
        );

    \tok.i5_4_lut_adj_203_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__20953\,
            in1 => \N__22969\,
            in2 => \N__20761\,
            in3 => \N__21047\,
            lcout => \tok.n21_adj_857\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i5_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12256\,
            in1 => \N__22101\,
            in2 => \_gnd_net_\,
            in3 => \N__15322\,
            lcout => uart_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i3_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16701\,
            in1 => \N__16942\,
            in2 => \_gnd_net_\,
            in3 => \N__21214\,
            lcout => capture_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_4_lut_adj_200_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__21169\,
            in1 => \N__20280\,
            in2 => \N__20400\,
            in3 => \N__22631\,
            lcout => \tok.n24_adj_854\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i7_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12270\,
            in1 => \N__16944\,
            in2 => \_gnd_net_\,
            in3 => \N__14929\,
            lcout => capture_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i6_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21340\,
            in1 => \N__12272\,
            in2 => \_gnd_net_\,
            in3 => \N__22102\,
            lcout => uart_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i6_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12271\,
            in1 => \N__16943\,
            in2 => \_gnd_net_\,
            in3 => \N__12255\,
            lcout => capture_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i2_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__12232\,
            in1 => \N__13300\,
            in2 => \N__16268\,
            in3 => \N__16427\,
            lcout => sender_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_2_lut_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17088\,
            in1 => \N__13139\,
            in2 => \N__29571\,
            in3 => \N__12185\,
            lcout => \tok.n6_adj_684\,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \tok.n3910\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_3_lut_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17643\,
            in1 => \N__14963\,
            in2 => \N__20170\,
            in3 => \N__12182\,
            lcout => \tok.n10_adj_786\,
            ltout => OPEN,
            carryin => \tok.n3910\,
            carryout => \tok.n3911\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_4_lut_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17086\,
            in1 => \N__12179\,
            in2 => \N__20064\,
            in3 => \N__12170\,
            lcout => \tok.n6_adj_667\,
            ltout => OPEN,
            carryin => \tok.n3911\,
            carryout => \tok.n3912\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_5_lut_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17642\,
            in1 => \N__15419\,
            in2 => \N__21550\,
            in3 => \N__12167\,
            lcout => \tok.n9_adj_836\,
            ltout => OPEN,
            carryin => \tok.n3912\,
            carryout => \tok.n3913\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_6_lut_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17644\,
            in1 => \N__24367\,
            in2 => \N__13220\,
            in3 => \N__12332\,
            lcout => \tok.n3_adj_826\,
            ltout => OPEN,
            carryin => \tok.n3913\,
            carryout => \tok.n3914\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_7_lut_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17090\,
            in1 => \N__15452\,
            in2 => \N__19946\,
            in3 => \N__12329\,
            lcout => \tok.n6_adj_814\,
            ltout => OPEN,
            carryin => \tok.n3914\,
            carryout => \tok.n3915\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_8_lut_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17087\,
            in1 => \N__21299\,
            in2 => \N__22739\,
            in3 => \N__12326\,
            lcout => \tok.n6_adj_780\,
            ltout => OPEN,
            carryin => \tok.n3915\,
            carryout => \tok.n3916\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_9_lut_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17089\,
            in1 => \N__12323\,
            in2 => \N__19689\,
            in3 => \N__12302\,
            lcout => \tok.n6_adj_768\,
            ltout => OPEN,
            carryin => \tok.n3916\,
            carryout => \tok.n3917\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_10_lut_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17109\,
            in1 => \N__19563\,
            in2 => \N__13247\,
            in3 => \N__12299\,
            lcout => \tok.n6_adj_653\,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \tok.n3918\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_11_lut_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17645\,
            in1 => \N__21180\,
            in2 => \N__14873\,
            in3 => \N__12296\,
            lcout => \tok.n13_adj_657\,
            ltout => OPEN,
            carryin => \tok.n3918\,
            carryout => \tok.n3919\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_12_lut_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17111\,
            in1 => \N__12377\,
            in2 => \N__20966\,
            in3 => \N__12293\,
            lcout => \tok.n6_adj_676\,
            ltout => OPEN,
            carryin => \tok.n3919\,
            carryout => \tok.n3920\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_13_lut_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17113\,
            in1 => \N__20867\,
            in2 => \N__12290\,
            in3 => \N__12275\,
            lcout => \tok.n6_adj_692\,
            ltout => OPEN,
            carryin => \tok.n3920\,
            carryout => \tok.n3921\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_14_lut_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17110\,
            in1 => \N__20762\,
            in2 => \N__12422\,
            in3 => \N__12401\,
            lcout => \tok.n6_adj_701\,
            ltout => OPEN,
            carryin => \tok.n3921\,
            carryout => \tok.n3922\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_15_lut_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17112\,
            in1 => \N__20563\,
            in2 => \N__13211\,
            in3 => \N__12398\,
            lcout => \tok.n6_adj_711\,
            ltout => OPEN,
            carryin => \tok.n3922\,
            carryout => \tok.n3923\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_16_lut_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17108\,
            in1 => \N__20505\,
            in2 => \N__12395\,
            in3 => \N__12383\,
            lcout => \tok.n6_adj_731\,
            ltout => OPEN,
            carryin => \tok.n3923\,
            carryout => \tok.n3924\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_16_THRU_CRY_0_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21610\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \tok.n3924\,
            carryout => \tok.n3924_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_17_lut_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__12371\,
            in1 => \N__20401\,
            in2 => \N__17117\,
            in3 => \N__12380\,
            lcout => \tok.n6_adj_753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i11_1_lut_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21059\,
            lcout => \tok.n292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i16_1_lut_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20305\,
            lcout => \tok.n287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i108_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14410\,
            in1 => \N__12520\,
            in2 => \N__12364\,
            in3 => \N__13504\,
            lcout => tail_108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26207\,
            ce => \N__14681\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i92_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13502\,
            in1 => \N__12511\,
            in2 => \N__12347\,
            in3 => \N__14416\,
            lcout => \tok.A_stk.tail_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26207\,
            ce => \N__14681\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i76_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14413\,
            in1 => \N__12521\,
            in2 => \N__12503\,
            in3 => \N__13506\,
            lcout => \tok.A_stk.tail_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26207\,
            ce => \N__14681\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i60_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13501\,
            in1 => \N__12512\,
            in2 => \N__12484\,
            in3 => \N__14415\,
            lcout => \tok.A_stk.tail_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26207\,
            ce => \N__14681\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i44_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14412\,
            in1 => \N__12499\,
            in2 => \N__12469\,
            in3 => \N__13505\,
            lcout => \tok.A_stk.tail_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26207\,
            ce => \N__14681\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i28_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13500\,
            in1 => \N__12455\,
            in2 => \N__12485\,
            in3 => \N__14414\,
            lcout => \tok.A_stk.tail_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26207\,
            ce => \N__14681\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i12_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__14411\,
            in1 => \N__13503\,
            in2 => \N__12470\,
            in3 => \N__20723\,
            lcout => \tok.A_stk.tail_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26207\,
            ce => \N__14681\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i12_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12454\,
            in1 => \N__15739\,
            in2 => \_gnd_net_\,
            in3 => \N__23006\,
            lcout => \tok.S_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26207\,
            ce => \N__14681\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i17_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__12431\,
            in1 => \N__12551\,
            in2 => \N__13876\,
            in3 => \N__14242\,
            lcout => \tok.A_stk.tail_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26211\,
            ce => \N__14664\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i1_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14239\,
            in1 => \N__12442\,
            in2 => \N__13723\,
            in3 => \N__20113\,
            lcout => \tok.A_stk.tail_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26211\,
            ce => \N__14664\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i33_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__12580\,
            in1 => \N__13524\,
            in2 => \N__12443\,
            in3 => \N__14243\,
            lcout => \tok.A_stk.tail_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26211\,
            ce => \N__14664\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i49_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14240\,
            in1 => \N__12430\,
            in2 => \N__13724\,
            in3 => \N__12569\,
            lcout => \tok.A_stk.tail_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26211\,
            ce => \N__14664\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i65_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__12560\,
            in1 => \N__13525\,
            in2 => \N__12581\,
            in3 => \N__14244\,
            lcout => \tok.A_stk.tail_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26211\,
            ce => \N__14664\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i81_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14241\,
            in1 => \N__13960\,
            in2 => \N__13725\,
            in3 => \N__12568\,
            lcout => \tok.A_stk.tail_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26211\,
            ce => \N__14664\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i97_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__12559\,
            in1 => \N__13526\,
            in2 => \N__13949\,
            in3 => \N__14245\,
            lcout => tail_97,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26211\,
            ce => \N__14664\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i1_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12550\,
            in1 => \N__15740\,
            in2 => \_gnd_net_\,
            in3 => \N__24188\,
            lcout => \tok.S_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26211\,
            ce => \N__14664\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i99_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14235\,
            in1 => \N__12541\,
            in2 => \N__13729\,
            in3 => \N__12688\,
            lcout => tail_99,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26216\,
            ce => \N__14682\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i35_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__12530\,
            in1 => \N__13537\,
            in2 => \N__12653\,
            in3 => \N__14237\,
            lcout => \tok.A_stk.tail_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26216\,
            ce => \N__14682\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i67_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14233\,
            in1 => \N__12529\,
            in2 => \N__13727\,
            in3 => \N__12689\,
            lcout => \tok.A_stk.tail_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26216\,
            ce => \N__14682\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i3_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12667\,
            in1 => \N__15724\,
            in2 => \_gnd_net_\,
            in3 => \N__21851\,
            lcout => \tok.S_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26216\,
            ce => \N__14682\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i51_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14232\,
            in1 => \N__12679\,
            in2 => \N__13726\,
            in3 => \N__12713\,
            lcout => \tok.A_stk.tail_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26216\,
            ce => \N__14682\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i101_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__12634\,
            in1 => \N__13536\,
            in2 => \N__12740\,
            in3 => \N__14236\,
            lcout => tail_101,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26216\,
            ce => \N__14682\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i85_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14234\,
            in1 => \N__12724\,
            in2 => \N__13728\,
            in3 => \N__12622\,
            lcout => \tok.A_stk.tail_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26216\,
            ce => \N__14682\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i83_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__12712\,
            in1 => \N__13538\,
            in2 => \N__12704\,
            in3 => \N__14238\,
            lcout => \tok.A_stk.tail_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26216\,
            ce => \N__14682\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i3_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__14247\,
            in1 => \N__13641\,
            in2 => \N__12652\,
            in3 => \N__21491\,
            lcout => \tok.A_stk.tail_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26224\,
            ce => \N__14712\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i19_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13638\,
            in1 => \N__12680\,
            in2 => \N__12668\,
            in3 => \N__14250\,
            lcout => \tok.A_stk.tail_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26224\,
            ce => \N__14712\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i69_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14249\,
            in1 => \N__12635\,
            in2 => \N__12607\,
            in3 => \N__13644\,
            lcout => \tok.A_stk.tail_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26224\,
            ce => \N__14712\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i53_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13640\,
            in1 => \N__12593\,
            in2 => \N__12623\,
            in3 => \N__14252\,
            lcout => \tok.A_stk.tail_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26224\,
            ce => \N__14712\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i37_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14246\,
            in1 => \N__12847\,
            in2 => \N__12608\,
            in3 => \N__13643\,
            lcout => \tok.A_stk.tail_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26224\,
            ce => \N__14712\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i21_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13639\,
            in1 => \N__12592\,
            in2 => \N__12839\,
            in3 => \N__14251\,
            lcout => \tok.A_stk.tail_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26224\,
            ce => \N__14712\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i5_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__14248\,
            in1 => \N__13642\,
            in2 => \N__19919\,
            in3 => \N__12848\,
            lcout => \tok.A_stk.tail_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26224\,
            ce => \N__14712\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i5_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12835\,
            in1 => \N__15681\,
            in2 => \_gnd_net_\,
            in3 => \N__22402\,
            lcout => \tok.S_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26224\,
            ce => \N__14712\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i100_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__12790\,
            in1 => \N__12827\,
            in2 => \N__13905\,
            in3 => \N__14385\,
            lcout => tail_100,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26229\,
            ce => \N__14722\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i84_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14383\,
            in1 => \N__12805\,
            in2 => \N__12781\,
            in3 => \N__13815\,
            lcout => \tok.A_stk.tail_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26229\,
            ce => \N__14722\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i68_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__12791\,
            in1 => \N__14387\,
            in2 => \N__13907\,
            in3 => \N__12766\,
            lcout => \tok.A_stk.tail_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26229\,
            ce => \N__14722\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i52_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14382\,
            in1 => \N__12757\,
            in2 => \N__12782\,
            in3 => \N__13814\,
            lcout => \tok.A_stk.tail_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26229\,
            ce => \N__14722\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i36_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__12748\,
            in1 => \N__14386\,
            in2 => \N__13906\,
            in3 => \N__12767\,
            lcout => \tok.A_stk.tail_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26229\,
            ce => \N__14722\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i20_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14381\,
            in1 => \N__12758\,
            in2 => \N__13013\,
            in3 => \N__13813\,
            lcout => \tok.A_stk.tail_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26229\,
            ce => \N__14722\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i4_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__12749\,
            in1 => \N__14384\,
            in2 => \N__24376\,
            in3 => \N__13645\,
            lcout => \tok.A_stk.tail_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26229\,
            ce => \N__14722\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i4_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13009\,
            in1 => \N__15731\,
            in2 => \_gnd_net_\,
            in3 => \N__27434\,
            lcout => \tok.S_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26229\,
            ce => \N__14722\,
            sr => \_gnd_net_\
        );

    \tok.i14_4_lut_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12857\,
            in1 => \N__12902\,
            in2 => \N__13001\,
            in3 => \N__12992\,
            lcout => OPEN,
            ltout => \tok.n30_adj_824_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4597_4_lut_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12986\,
            in1 => \N__15080\,
            in2 => \N__12980\,
            in3 => \N__15029\,
            lcout => OPEN,
            ltout => \tok.n4642_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_190_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__12977\,
            in1 => \N__14855\,
            in2 => \N__12971\,
            in3 => \N__22519\,
            lcout => \tok.found_slot\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.key_rd_15__I_0_241_i14_2_lut_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12968\,
            in2 => \_gnd_net_\,
            in3 => \N__20677\,
            lcout => \tok.n14_adj_804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i11_4_lut_adj_85_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12919\,
            in1 => \N__12877\,
            in2 => \N__12941\,
            in3 => \N__12895\,
            lcout => \tok.n27_adj_734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_70_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__12940\,
            in1 => \N__21034\,
            in2 => \N__12923\,
            in3 => \N__22979\,
            lcout => \tok.n21_adj_714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_44_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__12896\,
            in1 => \N__12881\,
            in2 => \N__19812\,
            in3 => \N__21967\,
            lcout => \tok.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_2_lut_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29078\,
            in1 => \N__29548\,
            in2 => \_gnd_net_\,
            in3 => \N__12851\,
            lcout => \tok.n10_adj_679\,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \tok.n3940\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_3_lut_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23746\,
            in1 => \N__20150\,
            in2 => \_gnd_net_\,
            in3 => \N__13049\,
            lcout => \tok.n28_adj_821\,
            ltout => OPEN,
            carryin => \tok.n3940\,
            carryout => \tok.n3941\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_4_lut_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29077\,
            in1 => \N__20035\,
            in2 => \_gnd_net_\,
            in3 => \N__13046\,
            lcout => \tok.n10_adj_818\,
            ltout => OPEN,
            carryin => \tok.n3941\,
            carryout => \tok.n3942\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_5_lut_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23745\,
            in1 => \_gnd_net_\,
            in2 => \N__21540\,
            in3 => \N__13043\,
            lcout => \tok.n6_adj_812\,
            ltout => OPEN,
            carryin => \tok.n3942\,
            carryout => \tok.n3943\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_6_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23744\,
            in1 => \N__24366\,
            in2 => \_gnd_net_\,
            in3 => \N__13040\,
            lcout => \tok.n9_adj_807\,
            ltout => OPEN,
            carryin => \tok.n3943\,
            carryout => \tok.n3944\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_7_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29080\,
            in1 => \N__19906\,
            in2 => \_gnd_net_\,
            in3 => \N__13037\,
            lcout => \tok.n10_adj_806\,
            ltout => OPEN,
            carryin => \tok.n3944\,
            carryout => \tok.n3945\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_8_lut_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29079\,
            in1 => \N__21298\,
            in2 => \_gnd_net_\,
            in3 => \N__13034\,
            lcout => \tok.n10_adj_783\,
            ltout => OPEN,
            carryin => \tok.n3945\,
            carryout => \tok.n3946\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_9_lut_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29081\,
            in1 => \N__19679\,
            in2 => \_gnd_net_\,
            in3 => \N__13022\,
            lcout => \tok.n10_adj_764\,
            ltout => OPEN,
            carryin => \tok.n3946\,
            carryout => \tok.n3947\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_10_lut_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29103\,
            in1 => \N__19549\,
            in2 => \_gnd_net_\,
            in3 => \N__13019\,
            lcout => \tok.n10_adj_652\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \tok.n3948\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_11_lut_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23750\,
            in1 => \N__21168\,
            in2 => \_gnd_net_\,
            in3 => \N__13016\,
            lcout => \tok.n10_adj_656\,
            ltout => OPEN,
            carryin => \tok.n3948\,
            carryout => \tok.n3949\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_12_lut_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29105\,
            in1 => \N__20952\,
            in2 => \_gnd_net_\,
            in3 => \N__13097\,
            lcout => \tok.n10_adj_671\,
            ltout => OPEN,
            carryin => \tok.n3949\,
            carryout => \tok.n3950\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_13_lut_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29108\,
            in1 => \N__20853\,
            in2 => \_gnd_net_\,
            in3 => \N__13094\,
            lcout => \tok.n4674\,
            ltout => OPEN,
            carryin => \tok.n3950\,
            carryout => \tok.n3951\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_14_lut_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29102\,
            in1 => \N__20732\,
            in2 => \_gnd_net_\,
            in3 => \N__13091\,
            lcout => \tok.n10_adj_697\,
            ltout => OPEN,
            carryin => \tok.n3951\,
            carryout => \tok.n3952\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_15_lut_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29107\,
            in1 => \N__20587\,
            in2 => \_gnd_net_\,
            in3 => \N__13088\,
            lcout => \tok.n10_adj_705\,
            ltout => OPEN,
            carryin => \tok.n3952\,
            carryout => \tok.n3953\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_16_lut_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29104\,
            in1 => \N__20506\,
            in2 => \_gnd_net_\,
            in3 => \N__13085\,
            lcout => \tok.n4661\,
            ltout => OPEN,
            carryin => \tok.n3953\,
            carryout => \tok.n3954\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_17_lut_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__20395\,
            in1 => \N__29106\,
            in2 => \_gnd_net_\,
            in3 => \N__13082\,
            lcout => \tok.n4656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_15_i2_3_lut_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__22717\,
            in1 => \N__21402\,
            in2 => \_gnd_net_\,
            in3 => \N__24494\,
            lcout => OPEN,
            ltout => \tok.n2_adj_739_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_89_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__21403\,
            in1 => \N__28348\,
            in2 => \N__13079\,
            in3 => \N__26810\,
            lcout => OPEN,
            ltout => \tok.n14_adj_741_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_96_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13076\,
            in1 => \N__15254\,
            in2 => \N__13064\,
            in3 => \N__13061\,
            lcout => OPEN,
            ltout => \tok.n20_adj_754_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4673_4_lut_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13181\,
            in1 => \N__13145\,
            in2 => \N__13175\,
            in3 => \N__13172\,
            lcout => \tok.n4653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_15_i9_2_lut_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20394\,
            in2 => \_gnd_net_\,
            in3 => \N__29461\,
            lcout => \tok.n9_adj_749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_adj_95_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__13163\,
            in1 => \N__20213\,
            in2 => \_gnd_net_\,
            in3 => \N__27245\,
            lcout => \tok.n16_adj_751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_inv_0_i1_1_lut_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26899\,
            lcout => \tok.n17_adj_774\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_65_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101111"
        )
    port map (
            in0 => \N__13133\,
            in1 => \N__22632\,
            in2 => \N__28349\,
            in3 => \N__26811\,
            lcout => \tok.n16_adj_706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_57_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100010001"
        )
    port map (
            in0 => \N__21400\,
            in1 => \N__26598\,
            in2 => \N__28270\,
            in3 => \N__24727\,
            lcout => \tok.n12_adj_687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_58_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__21841\,
            in1 => \N__21401\,
            in2 => \N__27072\,
            in3 => \N__17921\,
            lcout => OPEN,
            ltout => \tok.n13_adj_688_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_59_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13124\,
            in1 => \N__13310\,
            in2 => \N__13118\,
            in3 => \N__13115\,
            lcout => OPEN,
            ltout => \tok.n20_adj_693_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4672_4_lut_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17978\,
            in1 => \N__13109\,
            in2 => \N__13100\,
            in3 => \N__15134\,
            lcout => \tok.n4671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_adj_177_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__25792\,
            in1 => \N__13256\,
            in2 => \_gnd_net_\,
            in3 => \N__27242\,
            lcout => \tok.n16_adj_845\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i9_1_lut_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1660_3_lut_4_lut_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__23893\,
            in1 => \N__21539\,
            in2 => \N__23627\,
            in3 => \N__29305\,
            lcout => \tok.table_wr_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i5_1_lut_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27427\,
            lcout => \tok.n298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i14_1_lut_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20652\,
            lcout => \tok.n289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_adj_145_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__13202\,
            in1 => \N__23428\,
            in2 => \_gnd_net_\,
            in3 => \N__27243\,
            lcout => \tok.n16_adj_820\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__22701\,
            in1 => \N__22375\,
            in2 => \_gnd_net_\,
            in3 => \N__24493\,
            lcout => OPEN,
            ltout => \tok.n34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__22376\,
            in1 => \N__28344\,
            in2 => \N__13196\,
            in3 => \N__26816\,
            lcout => \tok.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_11_i2_3_lut_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__19806\,
            in1 => \_gnd_net_\,
            in2 => \N__22716\,
            in3 => \N__24492\,
            lcout => OPEN,
            ltout => \tok.n2_adj_685_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_56_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111101"
        )
    port map (
            in0 => \N__28337\,
            in1 => \N__19807\,
            in2 => \N__13313\,
            in3 => \N__26815\,
            lcout => \tok.n14_adj_686\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i1_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13304\,
            lcout => tx_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26263\,
            ce => \N__16386\,
            sr => \N__16465\
        );

    \tok.reset_I_0_1_lut_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13280\,
            lcout => \tok.reset_N_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i111_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__14005\,
            in1 => \N__13511\,
            in2 => \N__13985\,
            in3 => \N__14407\,
            lcout => tail_111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26212\,
            ce => \N__14680\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i15_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20310\,
            in1 => \N__15712\,
            in2 => \_gnd_net_\,
            in3 => \N__14026\,
            lcout => \tok.S_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26212\,
            ce => \N__14680\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i79_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__13273\,
            in1 => \N__13513\,
            in2 => \N__14009\,
            in3 => \N__14409\,
            lcout => \tok.A_stk.tail_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26212\,
            ce => \N__14680\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i63_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14404\,
            in1 => \N__13264\,
            in2 => \N__13721\,
            in3 => \N__14018\,
            lcout => \tok.A_stk.tail_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26212\,
            ce => \N__14680\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i47_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__13274\,
            in1 => \N__13512\,
            in2 => \N__14039\,
            in3 => \N__14408\,
            lcout => \tok.A_stk.tail_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26212\,
            ce => \N__14680\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i31_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14403\,
            in1 => \N__14027\,
            in2 => \N__13720\,
            in3 => \N__13265\,
            lcout => \tok.A_stk.tail_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26212\,
            ce => \N__14680\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i15_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__14038\,
            in1 => \N__14406\,
            in2 => \N__20369\,
            in3 => \N__13523\,
            lcout => \tok.A_stk.tail_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26212\,
            ce => \N__14680\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i95_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14405\,
            in1 => \N__13996\,
            in2 => \N__13722\,
            in3 => \N__14017\,
            lcout => \tok.A_stk.tail_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26212\,
            ce => \N__14680\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i127_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__14135\,
            in1 => \N__13981\,
            in2 => \N__13719\,
            in3 => \N__13997\,
            lcout => tail_127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_189_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__22520\,
            in1 => \N__15941\,
            in2 => \_gnd_net_\,
            in3 => \N__28832\,
            lcout => \tok.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i58_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__15478\,
            in1 => \N__25598\,
            in2 => \N__16580\,
            in3 => \N__25422\,
            lcout => \tok.tail_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i57_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__25420\,
            in1 => \N__15491\,
            in2 => \N__25660\,
            in3 => \N__15512\,
            lcout => \tok.tail_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i56_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__18493\,
            in1 => \N__25597\,
            in2 => \N__18470\,
            in3 => \N__25421\,
            lcout => \tok.tail_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i113_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__13945\,
            in1 => \N__13507\,
            in2 => \N__13964\,
            in3 => \N__14136\,
            lcout => tail_113,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_4_lut_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__28833\,
            in1 => \N__15597\,
            in2 => \N__16631\,
            in3 => \N__28691\,
            lcout => n29,
            ltout => \n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.i567_2_lut_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14741\,
            in3 => \N__14134\,
            lcout => \tok.A_stk.rd_15__N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_103_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__23110\,
            in1 => \N__30448\,
            in2 => \N__15224\,
            in3 => \N__30163\,
            lcout => OPEN,
            ltout => \tok.n83_adj_735_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4602_2_lut_3_lut_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29029\,
            in2 => \N__14588\,
            in3 => \N__29869\,
            lcout => \tok.n4649\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_155_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111101111111"
        )
    port map (
            in0 => \N__29868\,
            in1 => \N__30447\,
            in2 => \N__28544\,
            in3 => \N__30162\,
            lcout => OPEN,
            ltout => \tok.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_69_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__14582\,
            in1 => \N__14557\,
            in2 => \N__14585\,
            in3 => \N__29028\,
            lcout => \tok.n2503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4364_2_lut_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__28015\,
            in1 => \N__28689\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n4516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i0_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17180\,
            in1 => \N__14572\,
            in2 => \_gnd_net_\,
            in3 => \N__16960\,
            lcout => capture_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26225\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__28517\,
            in1 => \N__28690\,
            in2 => \N__30452\,
            in3 => \N__30164\,
            lcout => OPEN,
            ltout => \tok.n4_adj_654_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_173_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14558\,
            in1 => \N__28016\,
            in2 => \N__14546\,
            in3 => \N__29030\,
            lcout => n786,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_72_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__16801\,
            in1 => \N__30146\,
            in2 => \N__17563\,
            in3 => \N__30417\,
            lcout => OPEN,
            ltout => \tok.n83_adj_716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4631_2_lut_3_lut_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__29854\,
            in1 => \_gnd_net_\,
            in2 => \N__14804\,
            in3 => \N__28999\,
            lcout => \tok.n4690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_2_lut_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30145\,
            in2 => \_gnd_net_\,
            in3 => \N__29853\,
            lcout => OPEN,
            ltout => \tok.n12_adj_740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_134_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30416\,
            in1 => \N__14795\,
            in2 => \N__14801\,
            in3 => \N__15599\,
            lcout => OPEN,
            ltout => \tok.n12_adj_801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_153_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__28523\,
            in1 => \N__28822\,
            in2 => \N__14798\,
            in3 => \N__27999\,
            lcout => \tok.n240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i226_2_lut_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28678\,
            in2 => \_gnd_net_\,
            in3 => \N__28998\,
            lcout => \tok.n284\,
            ltout => \tok.n284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_99_i8_3_lut_4_lut_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001101"
        )
    port map (
            in0 => \N__28524\,
            in1 => \N__21846\,
            in2 => \N__14789\,
            in3 => \N__28821\,
            lcout => OPEN,
            ltout => \tok.n182_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_108_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__14899\,
            in1 => \N__27067\,
            in2 => \N__14786\,
            in3 => \N__26812\,
            lcout => \tok.n12_adj_766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i14_4_lut_adj_208_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16088\,
            in1 => \N__16058\,
            in2 => \N__14771\,
            in3 => \N__14756\,
            lcout => OPEN,
            ltout => \tok.n30_adj_862_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_210_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14942\,
            in2 => \N__14744\,
            in3 => \N__26486\,
            lcout => \tok.n4051\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_207_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__28253\,
            in1 => \N__29549\,
            in2 => \N__21303\,
            in3 => \N__26928\,
            lcout => \tok.n17_adj_861\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_206_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__20679\,
            in1 => \N__19555\,
            in2 => \N__20583\,
            in3 => \N__24794\,
            lcout => OPEN,
            ltout => \tok.n19_adj_860_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i13_4_lut_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15431\,
            in1 => \N__16094\,
            in2 => \N__14951\,
            in3 => \N__14948\,
            lcout => \tok.n29_adj_864\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i7_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__14936\,
            in1 => \N__22114\,
            in2 => \N__14903\,
            in3 => \_gnd_net_\,
            lcout => uart_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2575_2_lut_3_lut_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__29281\,
            in1 => \N__20947\,
            in2 => \_gnd_net_\,
            in3 => \N__23871\,
            lcout => \tok.table_wr_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i10_1_lut_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22650\,
            lcout => \tok.n293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2580_3_lut_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__29279\,
            in1 => \N__23869\,
            in2 => \_gnd_net_\,
            in3 => \N__26416\,
            lcout => \tok.n2634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_4_lut_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__26417\,
            in1 => \N__19371\,
            in2 => \N__23894\,
            in3 => \N__29282\,
            lcout => \tok.write_slot\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1586_3_lut_4_lut_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__29280\,
            in1 => \N__23383\,
            in2 => \N__19950\,
            in3 => \N__23870\,
            lcout => \tok.table_wr_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_97_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__24131\,
            in1 => \N__15122\,
            in2 => \N__15101\,
            in3 => \N__27435\,
            lcout => \tok.n18_adj_756\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_3_lut_4_lut_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__29283\,
            in1 => \N__22112\,
            in2 => \N__19313\,
            in3 => \N__27806\,
            lcout => \tok.uart.n922\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4599_4_lut_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__15074\,
            in1 => \N__28259\,
            in2 => \N__15053\,
            in3 => \N__26929\,
            lcout => \tok.n4645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_39_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__15020\,
            in1 => \N__15008\,
            in2 => \N__24149\,
            in3 => \N__27804\,
            lcout => OPEN,
            ltout => \tok.n30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_40_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__15002\,
            in1 => \N__29258\,
            in2 => \N__14990\,
            in3 => \N__27244\,
            lcout => \tok.n12_adj_659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.valid_54_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__29259\,
            in1 => \N__19299\,
            in2 => \_gnd_net_\,
            in3 => \N__27805\,
            lcout => \tok.uart_rx_valid\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26245\,
            ce => \N__14972\,
            sr => \_gnd_net_\
        );

    \tok.inv_106_i2_1_lut_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24118\,
            lcout => \tok.n301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_99_i6_3_lut_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011010"
        )
    port map (
            in0 => \N__29027\,
            in1 => \_gnd_net_\,
            in2 => \N__28700\,
            in3 => \N__24140\,
            lcout => \tok.n184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_142_i15_2_lut_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28692\,
            in2 => \_gnd_net_\,
            in3 => \N__29025\,
            lcout => OPEN,
            ltout => \tok.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i3_4_lut_adj_27_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30135\,
            in1 => \N__29848\,
            in2 => \N__15236\,
            in3 => \N__28528\,
            lcout => \tok.n880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_99_i7_3_lut_4_lut_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110101"
        )
    port map (
            in0 => \N__28529\,
            in1 => \N__28693\,
            in2 => \N__21971\,
            in3 => \N__29026\,
            lcout => \tok.n183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_117_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__21866\,
            in1 => \N__24473\,
            in2 => \N__15233\,
            in3 => \N__26790\,
            lcout => OPEN,
            ltout => \tok.n16_adj_778_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_4_lut_adj_119_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__15220\,
            in1 => \N__27209\,
            in2 => \N__15194\,
            in3 => \N__15191\,
            lcout => \tok.n20_adj_781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_0_i1_2_lut_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26789\,
            in2 => \_gnd_net_\,
            in3 => \N__30148\,
            lcout => \tok.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4624_4_lut_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__20588\,
            in1 => \N__27211\,
            in2 => \N__15179\,
            in3 => \N__29411\,
            lcout => \tok.n4664\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_adj_46_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__27208\,
            in1 => \N__20882\,
            in2 => \_gnd_net_\,
            in3 => \N__15167\,
            lcout => OPEN,
            ltout => \tok.n14_adj_669_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_48_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__27063\,
            in1 => \N__15155\,
            in2 => \N__15149\,
            in3 => \N__21957\,
            lcout => \tok.n18_adj_672\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__15146\,
            in1 => \N__27210\,
            in2 => \_gnd_net_\,
            in3 => \N__20774\,
            lcout => \tok.n16_adj_691\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i9_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__17499\,
            in1 => \N__17370\,
            in2 => \N__19571\,
            in3 => \N__17936\,
            lcout => \tok.n60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26255\,
            ce => \N__17252\,
            sr => \N__19118\
        );

    \tok.A_i16_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__20368\,
            in1 => \N__17500\,
            in2 => \N__17385\,
            in3 => \N__15305\,
            lcout => \tok.n53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26255\,
            ce => \N__17252\,
            sr => \N__19118\
        );

    \tok.A_i12_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__17498\,
            in1 => \N__17369\,
            in2 => \N__20868\,
            in3 => \N__15299\,
            lcout => \tok.n57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26255\,
            ce => \N__17252\,
            sr => \N__19118\
        );

    \tok.i9_4_lut_adj_50_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__24729\,
            in1 => \N__15242\,
            in2 => \N__15293\,
            in3 => \N__22373\,
            lcout => OPEN,
            ltout => \tok.n20_adj_674_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4674_4_lut_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__15248\,
            in1 => \N__15284\,
            in2 => \N__15272\,
            in3 => \N__15269\,
            lcout => OPEN,
            ltout => \tok.n4676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i11_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011101110"
        )
    port map (
            in0 => \N__17368\,
            in1 => \N__20954\,
            in2 => \N__15257\,
            in3 => \N__17501\,
            lcout => \tok.n58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26255\,
            ce => \N__17252\,
            sr => \N__19118\
        );

    \tok.i1_4_lut_adj_91_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000011"
        )
    port map (
            in0 => \N__21032\,
            in1 => \N__26622\,
            in2 => \N__20287\,
            in3 => \N__24728\,
            lcout => \tok.n12_adj_744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4371_2_lut_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26623\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21033\,
            lcout => \tok.n4524\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_47_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__26804\,
            in1 => \N__21031\,
            in2 => \N__28148\,
            in3 => \N__17908\,
            lcout => \tok.n12_adj_670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_14_i2_3_lut_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__21029\,
            in1 => \N__22720\,
            in2 => \_gnd_net_\,
            in3 => \N__24485\,
            lcout => OPEN,
            ltout => \tok.n2_adj_720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_76_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110001"
        )
    port map (
            in0 => \N__26803\,
            in1 => \N__28325\,
            in2 => \N__15404\,
            in3 => \N__21030\,
            lcout => \tok.n14_adj_722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_79_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__23984\,
            in1 => \N__28264\,
            in2 => \N__27071\,
            in3 => \N__17909\,
            lcout => OPEN,
            ltout => \tok.n13_adj_726_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_83_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15401\,
            in1 => \N__15395\,
            in2 => \N__15383\,
            in3 => \N__15380\,
            lcout => OPEN,
            ltout => \tok.n20_adj_732_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4671_4_lut_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15371\,
            in1 => \N__17132\,
            in2 => \N__15359\,
            in3 => \N__15347\,
            lcout => \tok.n4658\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_14_i9_2_lut_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__20509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29440\,
            lcout => \tok.n9_adj_728\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_142_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__15341\,
            in1 => \N__27057\,
            in2 => \N__15329\,
            in3 => \N__26813\,
            lcout => OPEN,
            ltout => \tok.n12_adj_815_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_146_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__24073\,
            in1 => \N__20641\,
            in2 => \N__15308\,
            in3 => \N__16292\,
            lcout => OPEN,
            ltout => \tok.n20_adj_822_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_151_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__15467\,
            in1 => \N__17497\,
            in2 => \N__15458\,
            in3 => \N__16286\,
            lcout => \tok.A_15_N_113_5\,
            ltout => \tok.A_15_N_113_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A__15__I_16_i6_3_lut_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22334\,
            in2 => \N__15455\,
            in3 => \N__17749\,
            lcout => \tok.A_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__24491\,
            in1 => \N__19570\,
            in2 => \N__15440\,
            in3 => \N__29445\,
            lcout => \tok.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i6_1_lut_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22333\,
            lcout => \tok.n297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_101_i9_2_lut_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22721\,
            in2 => \_gnd_net_\,
            in3 => \N__27428\,
            lcout => \tok.n208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_204_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__21832\,
            in1 => \N__21538\,
            in2 => \N__19949\,
            in3 => \N__22332\,
            lcout => \tok.n20_adj_858\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i4_1_lut_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21831\,
            lcout => \tok.n299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_30_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__22528\,
            in1 => \N__19817\,
            in2 => \N__22277\,
            in3 => \N__17999\,
            lcout => OPEN,
            ltout => \tok.n27_adj_644_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i7_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__19280\,
            in1 => \N__18037\,
            in2 => \N__15407\,
            in3 => \N__18974\,
            lcout => \tok.n39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26266\,
            ce => 'H',
            sr => \N__19096\
        );

    \tok.idx_i5_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111001101010000"
        )
    port map (
            in0 => \N__18973\,
            in1 => \N__19279\,
            in2 => \N__18114\,
            in3 => \N__22190\,
            lcout => \tok.n44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26266\,
            ce => 'H',
            sr => \N__19096\
        );

    \tok.C_stk.tail_i0_i9_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15545\,
            in1 => \N__16822\,
            in2 => \_gnd_net_\,
            in3 => \N__25588\,
            lcout => \tok.tail_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26218\,
            ce => \N__25426\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i1_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25581\,
            in1 => \N__15554\,
            in2 => \_gnd_net_\,
            in3 => \N__16805\,
            lcout => \tok.C_stk.tail_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26218\,
            ce => \N__25426\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i17_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__15553\,
            in1 => \_gnd_net_\,
            in2 => \N__15536\,
            in3 => \N__25585\,
            lcout => \tok.C_stk.tail_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26218\,
            ce => \N__25426\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i25_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25582\,
            in1 => \N__15544\,
            in2 => \_gnd_net_\,
            in3 => \N__15521\,
            lcout => \tok.tail_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26218\,
            ce => \N__25426\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i33_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15532\,
            in1 => \N__15500\,
            in2 => \_gnd_net_\,
            in3 => \N__25586\,
            lcout => \tok.C_stk.tail_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26218\,
            ce => \N__25426\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i41_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25583\,
            in1 => \N__15490\,
            in2 => \_gnd_net_\,
            in3 => \N__15520\,
            lcout => \tok.tail_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26218\,
            ce => \N__25426\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i49_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15511\,
            in1 => \N__15499\,
            in2 => \_gnd_net_\,
            in3 => \N__25587\,
            lcout => \tok.tail_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26218\,
            ce => \N__25426\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i50_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__25584\,
            in1 => \N__15479\,
            in2 => \N__16550\,
            in3 => \_gnd_net_\,
            lcout => \tok.tail_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26218\,
            ce => \N__25426\,
            sr => \_gnd_net_\
        );

    \tok.i2559_2_lut_4_lut_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16616\,
            in1 => \N__15598\,
            in2 => \N__16685\,
            in3 => \N__15578\,
            lcout => \tok.C_stk_delta_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_135_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16049\,
            in2 => \_gnd_net_\,
            in3 => \N__15817\,
            lcout => \tok.n875\,
            ltout => \tok.n875_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2510_2_lut_3_lut_4_lut_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22521\,
            in1 => \N__15784\,
            in2 => \N__15602\,
            in3 => \N__15895\,
            lcout => \tok.n2562\,
            ltout => \tok.n2562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i568_2_lut_4_lut_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101010101"
        )
    port map (
            in0 => \N__15577\,
            in1 => \N__16680\,
            in2 => \N__15569\,
            in3 => \N__16615\,
            lcout => \tok.rd_7__N_374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4325_2_lut_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__15818\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15897\,
            lcout => OPEN,
            ltout => \tok.n4474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_115_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__15786\,
            in1 => \N__16681\,
            in2 => \N__15566\,
            in3 => \N__16050\,
            lcout => \tok.n802\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_142_i20_2_lut_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15785\,
            in2 => \_gnd_net_\,
            in3 => \N__15896\,
            lcout => OPEN,
            ltout => \tok.n20_adj_772_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_113_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__15563\,
            in1 => \N__28829\,
            in2 => \N__15557\,
            in3 => \N__28017\,
            lcout => \tok.n4446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_i3_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011110101000010"
        )
    port map (
            in0 => \N__15911\,
            in1 => \N__15860\,
            in2 => \N__15899\,
            in3 => \N__15788\,
            lcout => \tok.n61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26230\,
            ce => 'H',
            sr => \N__19131\
        );

    \tok.depth_i1_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001011011110000"
        )
    port map (
            in0 => \N__16048\,
            in1 => \N__15943\,
            in2 => \N__15823\,
            in3 => \N__16008\,
            lcout => \tok.n63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26230\,
            ce => 'H',
            sr => \N__19131\
        );

    \tok.i2_4_lut_4_lut_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011011110000"
        )
    port map (
            in0 => \N__15942\,
            in1 => \N__16047\,
            in2 => \N__15824\,
            in3 => \N__16002\,
            lcout => \tok.depth_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_4_lut_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15813\,
            in1 => \N__15783\,
            in2 => \N__16052\,
            in3 => \N__15889\,
            lcout => \tok.A_stk_delta_1__N_4\,
            ltout => \tok.A_stk_delta_1__N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__15819\,
            in1 => \N__16046\,
            in2 => \N__15791\,
            in3 => \N__16001\,
            lcout => \tok.n4_adj_809\,
            ltout => \tok.n4_adj_809_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_196_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101101010"
        )
    port map (
            in0 => \N__15787\,
            in1 => \N__15890\,
            in2 => \N__15761\,
            in3 => \N__15909\,
            lcout => OPEN,
            ltout => \tok.depth_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_197_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15758\,
            in3 => \N__15755\,
            lcout => \tok.n6_adj_853\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_i2_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15859\,
            in1 => \N__15894\,
            in2 => \_gnd_net_\,
            in3 => \N__15910\,
            lcout => \tok.n62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26230\,
            ce => 'H',
            sr => \N__19131\
        );

    \tok.i4353_2_lut_3_lut_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__22492\,
            in1 => \N__28812\,
            in2 => \_gnd_net_\,
            in3 => \N__28512\,
            lcout => \tok.n4504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4400_2_lut_4_lut_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28513\,
            in1 => \N__22493\,
            in2 => \N__28831\,
            in3 => \N__15940\,
            lcout => OPEN,
            ltout => \tok.n4554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_164_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27993\,
            in1 => \N__27311\,
            in2 => \N__15749\,
            in3 => \N__15962\,
            lcout => \tok.n237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_161_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28662\,
            in2 => \_gnd_net_\,
            in3 => \N__28972\,
            lcout => \tok.n6_adj_832\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_194_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000010"
        )
    port map (
            in0 => \N__27992\,
            in1 => \N__30394\,
            in2 => \N__15944\,
            in3 => \N__30137\,
            lcout => OPEN,
            ltout => \tok.n4432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_195_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15961\,
            in1 => \N__15953\,
            in2 => \N__15947\,
            in3 => \N__29852\,
            lcout => \tok.n1_adj_802\,
            ltout => \tok.n1_adj_802_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2578_2_lut_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__15939\,
            in1 => \_gnd_net_\,
            in2 => \N__15914\,
            in3 => \_gnd_net_\,
            lcout => \tok.n189\,
            ltout => \tok.n189_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_192_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__15898\,
            in1 => \_gnd_net_\,
            in2 => \N__15863\,
            in3 => \N__15858\,
            lcout => \tok.depth_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i11_4_lut_adj_128_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22996\,
            in1 => \N__21937\,
            in2 => \N__19825\,
            in3 => \N__21054\,
            lcout => OPEN,
            ltout => \tok.n27_adj_793_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i15_4_lut_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15836\,
            in1 => \N__15830\,
            in2 => \N__15845\,
            in3 => \N__15842\,
            lcout => \tok.tc__7__N_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_129_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24129\,
            in1 => \N__28254\,
            in2 => \N__27446\,
            in3 => \N__26927\,
            lcout => \tok.n25_adj_794\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_127_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22366\,
            in1 => \N__21839\,
            in2 => \N__24847\,
            in3 => \N__20678\,
            lcout => \tok.n26_adj_792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i12_4_lut_adj_126_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24013\,
            in1 => \N__22655\,
            in2 => \N__20309\,
            in3 => \N__21428\,
            lcout => \tok.n28_adj_791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_205_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__20143\,
            in1 => \N__27433\,
            in2 => \N__24368\,
            in3 => \N__24130\,
            lcout => \tok.n18_adj_859\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_201_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__20042\,
            in1 => \N__19813\,
            in2 => \N__19660\,
            in3 => \N__21938\,
            lcout => \tok.n22_adj_855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i3_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17344\,
            in1 => \N__20043\,
            in2 => \_gnd_net_\,
            in3 => \N__16856\,
            lcout => \tok.A_low_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26246\,
            ce => \N__17268\,
            sr => \N__19142\
        );

    \tok.i2_3_lut_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__16075\,
            in1 => \N__16520\,
            in2 => \_gnd_net_\,
            in3 => \N__30411\,
            lcout => \tok.n23\,
            ltout => \tok.n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i2_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20155\,
            in2 => \N__16061\,
            in3 => \N__16127\,
            lcout => \tok.A_low_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26246\,
            ce => \N__17268\,
            sr => \N__19142\
        );

    \tok.i7_4_lut_adj_202_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__20857\,
            in1 => \N__24008\,
            in2 => \N__20508\,
            in3 => \N__21410\,
            lcout => \tok.n23_adj_856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_i0_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__16010\,
            in1 => \_gnd_net_\,
            in2 => \N__16051\,
            in3 => \_gnd_net_\,
            lcout => \tok.n64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26250\,
            ce => 'H',
            sr => \N__19114\
        );

    \tok.i1_2_lut_adj_193_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16039\,
            in2 => \_gnd_net_\,
            in3 => \N__16009\,
            lcout => OPEN,
            ltout => \tok.depth_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_199_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22503\,
            in1 => \N__15983\,
            in2 => \N__15974\,
            in3 => \N__15971\,
            lcout => \tok.A__15__N_129\,
            ltout => \tok.A__15__N_129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A__15__I_16_i3_3_lut_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21942\,
            in2 => \N__16112\,
            in3 => \N__16855\,
            lcout => \tok.A_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_214_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__21823\,
            in1 => \N__22237\,
            in2 => \N__22522\,
            in3 => \N__18236\,
            lcout => \tok.n27_adj_866\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.search_clk_198_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22239\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.search_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26250\,
            ce => 'H',
            sr => \N__19114\
        );

    \tok.i50_4_lut_adj_216_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__22507\,
            in1 => \N__22238\,
            in2 => \N__18155\,
            in3 => \N__27429\,
            lcout => OPEN,
            ltout => \tok.n27_adj_867_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i4_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__19260\,
            in1 => \N__18174\,
            in2 => \N__16109\,
            in3 => \N__18954\,
            lcout => \tok.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26250\,
            ce => 'H',
            sr => \N__19114\
        );

    \tok.i4390_2_lut_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__30150\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24705\,
            lcout => \tok.n4544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_2_lut_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__21685\,
            in1 => \N__22181\,
            in2 => \_gnd_net_\,
            in3 => \N__30149\,
            lcout => \tok.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_52_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111011"
        )
    port map (
            in0 => \N__26925\,
            in1 => \N__26604\,
            in2 => \N__16106\,
            in3 => \N__17904\,
            lcout => OPEN,
            ltout => \tok.n14_adj_678_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_54_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011111111"
        )
    port map (
            in0 => \N__17155\,
            in1 => \N__27062\,
            in2 => \N__16097\,
            in3 => \N__17509\,
            lcout => OPEN,
            ltout => \tok.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18929\,
            in1 => \N__16169\,
            in2 => \N__16163\,
            in3 => \N__29342\,
            lcout => OPEN,
            ltout => \tok.n22_adj_683_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i11_4_lut_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__16160\,
            in1 => \N__24200\,
            in2 => \N__16148\,
            in3 => \N__16145\,
            lcout => \tok.A_15_N_113_0\,
            ltout => \tok.A_15_N_113_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A__15__I_16_i1_3_lut_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26926\,
            in1 => \_gnd_net_\,
            in2 => \N__16139\,
            in3 => \N__17715\,
            lcout => \tok.A_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_171_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__21449\,
            in1 => \N__24242\,
            in2 => \N__17520\,
            in3 => \N__16136\,
            lcout => \tok.A_15_N_113_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i44_3_lut_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21795\,
            in1 => \N__26618\,
            in2 => \_gnd_net_\,
            in3 => \N__17890\,
            lcout => \tok.n4520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_3_lut_adj_187_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__17891\,
            in1 => \_gnd_net_\,
            in2 => \N__26624\,
            in3 => \N__24168\,
            lcout => OPEN,
            ltout => \tok.n46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_188_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__17534\,
            in1 => \N__17508\,
            in2 => \N__16130\,
            in3 => \N__17573\,
            lcout => \tok.A_15_N_113_1\,
            ltout => \tok.A_15_N_113_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A__15__I_16_i2_3_lut_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17738\,
            in2 => \N__16118\,
            in3 => \N__24169\,
            lcout => OPEN,
            ltout => \tok.A_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16467\,
            in1 => \_gnd_net_\,
            in2 => \N__16115\,
            in3 => \N__16247\,
            lcout => \tok.uart.sender_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26261\,
            ce => \N__16388\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i3_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16280\,
            in1 => \N__16466\,
            in2 => \_gnd_net_\,
            in3 => \N__16274\,
            lcout => sender_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26261\,
            ce => \N__16388\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i5_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16468\,
            in1 => \N__16397\,
            in2 => \_gnd_net_\,
            in3 => \N__16256\,
            lcout => \tok.uart.sender_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26261\,
            ce => \N__16388\,
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_118_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__26603\,
            in1 => \N__28218\,
            in2 => \_gnd_net_\,
            in3 => \N__17889\,
            lcout => OPEN,
            ltout => \tok.n14_adj_779_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_121_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16241\,
            in1 => \N__19841\,
            in2 => \N__16229\,
            in3 => \N__16226\,
            lcout => OPEN,
            ltout => \tok.n22_adj_784_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_123_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__21233\,
            in1 => \N__17521\,
            in2 => \N__16214\,
            in3 => \N__23909\,
            lcout => \tok.A_15_N_113_6\,
            ltout => \tok.A_15_N_113_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A__15__I_16_i7_3_lut_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28219\,
            in1 => \_gnd_net_\,
            in2 => \N__16211\,
            in3 => \N__17748\,
            lcout => OPEN,
            ltout => \tok.A_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i9_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16472\,
            in1 => \_gnd_net_\,
            in2 => \N__16208\,
            in3 => \N__16205\,
            lcout => \tok.uart.sender_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26264\,
            ce => \N__16387\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i8_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16187\,
            in1 => \N__16471\,
            in2 => \_gnd_net_\,
            in3 => \N__16181\,
            lcout => \tok.uart.sender_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26264\,
            ce => \N__16387\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i7_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16470\,
            in1 => \N__16175\,
            in2 => \_gnd_net_\,
            in3 => \N__17528\,
            lcout => \tok.uart.sender_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26264\,
            ce => \N__16387\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i6_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16478\,
            in1 => \N__16469\,
            in2 => \_gnd_net_\,
            in3 => \N__17684\,
            lcout => \tok.uart.sender_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26264\,
            ce => \N__16387\,
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_66_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001011101"
        )
    port map (
            in0 => \N__26602\,
            in1 => \N__22349\,
            in2 => \N__27073\,
            in3 => \N__20642\,
            lcout => \tok.n14_adj_707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_4_lut_adj_67_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__20643\,
            in1 => \N__16337\,
            in2 => \N__22541\,
            in3 => \N__17881\,
            lcout => OPEN,
            ltout => \tok.n20_adj_708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_68_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__17522\,
            in1 => \N__16325\,
            in2 => \N__16319\,
            in3 => \N__24635\,
            lcout => OPEN,
            ltout => \tok.n22_adj_709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i14_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__17378\,
            in1 => \N__22763\,
            in2 => \N__16316\,
            in3 => \N__20597\,
            lcout => \tok.n55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26267\,
            ce => \N__17267\,
            sr => \N__19066\
        );

    \tok.A_i6_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19948\,
            in1 => \N__17379\,
            in2 => \_gnd_net_\,
            in3 => \N__16313\,
            lcout => \tok.A_low_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26267\,
            ce => \N__17267\,
            sr => \N__19066\
        );

    \tok.i2_4_lut_adj_140_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111111011"
        )
    port map (
            in0 => \N__16307\,
            in1 => \N__26601\,
            in2 => \N__22374\,
            in3 => \N__17880\,
            lcout => OPEN,
            ltout => \tok.n13_adj_813_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_144_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__19947\,
            in1 => \N__22805\,
            in2 => \N__16295\,
            in3 => \N__29444\,
            lcout => \tok.n18_adj_819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_149_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111000"
        )
    port map (
            in0 => \N__26920\,
            in1 => \N__24735\,
            in2 => \N__19862\,
            in3 => \N__28698\,
            lcout => \tok.n15_adj_823\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_43_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__17759\,
            in1 => \N__26921\,
            in2 => \N__22529\,
            in3 => \N__22272\,
            lcout => \tok.n27_adj_664\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_209_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__22527\,
            in1 => \N__18374\,
            in2 => \N__22282\,
            in3 => \N__24185\,
            lcout => OPEN,
            ltout => \tok.n27_adj_863_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i1_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__19276\,
            in1 => \N__18408\,
            in2 => \N__16502\,
            in3 => \N__18970\,
            lcout => \tok.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26269\,
            ce => 'H',
            sr => \N__19086\
        );

    \tok.i50_4_lut_adj_212_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__22273\,
            in1 => \N__22526\,
            in2 => \N__18308\,
            in3 => \N__21972\,
            lcout => OPEN,
            ltout => \tok.n27_adj_865_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i2_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__19277\,
            in1 => \N__18334\,
            in2 => \N__16499\,
            in3 => \N__18971\,
            lcout => \tok.n49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26269\,
            ce => 'H',
            sr => \N__19086\
        );

    \tok.idx_i0_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__18969\,
            in1 => \N__16496\,
            in2 => \N__17796\,
            in3 => \N__19275\,
            lcout => \tok.n52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26269\,
            ce => 'H',
            sr => \N__19086\
        );

    \tok.idx_i3_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__19278\,
            in1 => \N__18972\,
            in2 => \N__18273\,
            in3 => \N__16490\,
            lcout => \tok.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26269\,
            ce => 'H',
            sr => \N__19086\
        );

    \tok.C_stk.tail_i0_i26_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16559\,
            in1 => \N__23323\,
            in2 => \_gnd_net_\,
            in3 => \N__25594\,
            lcout => \tok.tail_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26226\,
            ce => \N__25427\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i34_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__25590\,
            in1 => \N__18535\,
            in2 => \N__16549\,
            in3 => \_gnd_net_\,
            lcout => \tok.C_stk.tail_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26226\,
            ce => \N__25427\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i36_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23344\,
            in1 => \N__16531\,
            in2 => \_gnd_net_\,
            in3 => \N__25596\,
            lcout => \tok.C_stk.tail_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26226\,
            ce => \N__25427\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i42_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25592\,
            in1 => \_gnd_net_\,
            in2 => \N__16576\,
            in3 => \N__16558\,
            lcout => \tok.tail_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26226\,
            ce => \N__25427\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i20_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18523\,
            in1 => \N__16532\,
            in2 => \_gnd_net_\,
            in3 => \N__25593\,
            lcout => \tok.C_stk.tail_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26226\,
            ce => \N__25427\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i32_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25589\,
            in1 => \N__18482\,
            in2 => \_gnd_net_\,
            in3 => \N__23156\,
            lcout => \tok.C_stk.tail_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26226\,
            ce => \N__25427\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i28_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17989\,
            in1 => \N__18512\,
            in2 => \_gnd_net_\,
            in3 => \N__25595\,
            lcout => \tok.tail_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26226\,
            ce => \N__25427\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i40_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25591\,
            in1 => \N__18460\,
            in2 => \_gnd_net_\,
            in3 => \N__23167\,
            lcout => \tok.tail_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26226\,
            ce => \N__25427\,
            sr => \_gnd_net_\
        );

    \tok.i127_4_lut_4_lut_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010000111111"
        )
    port map (
            in0 => \N__30445\,
            in1 => \N__29870\,
            in2 => \N__28555\,
            in3 => \N__30157\,
            lcout => OPEN,
            ltout => \tok.n127_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_116_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111110"
        )
    port map (
            in0 => \N__29871\,
            in1 => \N__25872\,
            in2 => \N__16523\,
            in3 => \N__29032\,
            lcout => OPEN,
            ltout => \tok.n4394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_124_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__16516\,
            in1 => \N__27310\,
            in2 => \N__16505\,
            in3 => \N__28697\,
            lcout => \tok.n86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29872\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30446\,
            lcout => OPEN,
            ltout => \tok.n28_adj_834_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4564_4_lut_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__29033\,
            in1 => \N__28019\,
            in2 => \N__16637\,
            in3 => \N__30159\,
            lcout => OPEN,
            ltout => \tok.n4604_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i49_4_lut_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__17600\,
            in1 => \N__29034\,
            in2 => \N__16634\,
            in3 => \N__28548\,
            lcout => \tok.n34_adj_719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__30444\,
            in1 => \N__18598\,
            in2 => \N__24233\,
            in3 => \N__30158\,
            lcout => \tok.n83_adj_704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_125_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29031\,
            in2 => \_gnd_net_\,
            in3 => \N__30443\,
            lcout => \tok.n101_adj_776\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4567_4_lut_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010000000"
        )
    port map (
            in0 => \N__29866\,
            in1 => \N__29008\,
            in2 => \N__30442\,
            in3 => \N__30154\,
            lcout => OPEN,
            ltout => \tok.n4610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i58_4_lut_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__30155\,
            in1 => \N__16670\,
            in2 => \N__16619\,
            in3 => \N__28530\,
            lcout => \tok.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_131_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010001000"
        )
    port map (
            in0 => \N__30423\,
            in1 => \N__16607\,
            in2 => \N__18744\,
            in3 => \N__30156\,
            lcout => OPEN,
            ltout => \tok.n83_adj_796_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4604_2_lut_3_lut_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__29009\,
            in1 => \_gnd_net_\,
            in2 => \N__16583\,
            in3 => \N__29867\,
            lcout => \tok.n4602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_133_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__25183\,
            in1 => \N__18880\,
            in2 => \N__25259\,
            in3 => \N__18698\,
            lcout => n92_adj_872,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i2_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16975\,
            in1 => \N__16718\,
            in2 => \_gnd_net_\,
            in3 => \N__16964\,
            lcout => capture_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_73_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__28679\,
            in1 => \N__28828\,
            in2 => \_gnd_net_\,
            in3 => \N__28018\,
            lcout => \tok.n847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i59_3_lut_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__29007\,
            in1 => \N__30419\,
            in2 => \_gnd_net_\,
            in3 => \N__29865\,
            lcout => \tok.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.n602_bdd_4_lut_4749_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__18913\,
            in1 => \N__25107\,
            in2 => \N__26358\,
            in3 => \N__18802\,
            lcout => OPEN,
            ltout => \tok.C_stk.n4906_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i6_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__24962\,
            in1 => \N__23098\,
            in2 => \N__16661\,
            in3 => \N__26352\,
            lcout => \tok.c_stk_r_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i4641_4_lut_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__18911\,
            in1 => \N__26684\,
            in2 => \N__23106\,
            in3 => \N__25990\,
            lcout => OPEN,
            ltout => \tok.ram.n4699_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5_4_lut_adj_25_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__23099\,
            in1 => \N__25897\,
            in2 => \N__16658\,
            in3 => \N__29855\,
            lcout => OPEN,
            ltout => \tok.n1_adj_760_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_104_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__16655\,
            in1 => \N__28550\,
            in2 => \N__16643\,
            in3 => \N__30147\,
            lcout => OPEN,
            ltout => \tok.n13_adj_761_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_106_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__25260\,
            in1 => \N__25189\,
            in2 => \N__16640\,
            in3 => \N__18912\,
            lcout => n92_adj_871,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18856\,
            in1 => \N__18840\,
            in2 => \_gnd_net_\,
            in3 => \N__23516\,
            lcout => \tok.tc_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.n602_bdd_4_lut_4719_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001011000"
        )
    port map (
            in0 => \N__26345\,
            in1 => \N__18643\,
            in2 => \N__25112\,
            in3 => \N__18765\,
            lcout => OPEN,
            ltout => \tok.C_stk.n4870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__16829\,
            in1 => \N__16788\,
            in2 => \N__16811\,
            in3 => \N__26346\,
            lcout => \tok.c_stk_r_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i4662_4_lut_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__26696\,
            in1 => \N__18641\,
            in2 => \N__16794\,
            in3 => \N__25983\,
            lcout => OPEN,
            ltout => \tok.ram.n4714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5_4_lut_adj_20_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__29847\,
            in1 => \N__25898\,
            in2 => \N__16808\,
            in3 => \N__16787\,
            lcout => OPEN,
            ltout => \tok.n1_adj_717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i18_4_lut_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__28554\,
            in1 => \N__16766\,
            in2 => \N__16754\,
            in3 => \N__30134\,
            lcout => OPEN,
            ltout => \tok.n5_adj_718_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_74_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__18642\,
            in1 => \N__25261\,
            in2 => \N__16751\,
            in3 => \N__25190\,
            lcout => n92,
            ltout => \n92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_147_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23498\,
            in2 => \N__16748\,
            in3 => \N__18766\,
            lcout => \tok.tc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_182_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__16730\,
            in1 => \N__27275\,
            in2 => \N__22658\,
            in3 => \N__26435\,
            lcout => OPEN,
            ltout => \tok.n6_adj_848_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_183_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__17008\,
            in1 => \N__17027\,
            in2 => \N__17015\,
            in3 => \N__27794\,
            lcout => OPEN,
            ltout => \tok.n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_184_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__29247\,
            in1 => \N__30410\,
            in2 => \N__17012\,
            in3 => \N__24269\,
            lcout => \tok.n10_adj_849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__17009\,
            in1 => \_gnd_net_\,
            in2 => \N__16985\,
            in3 => \N__22113\,
            lcout => uart_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1549_3_lut_4_lut_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__23867\,
            in1 => \N__18917\,
            in2 => \N__29284\,
            in3 => \N__21320\,
            lcout => \tok.table_wr_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17172\,
            in1 => \N__16981\,
            in2 => \_gnd_net_\,
            in3 => \N__16953\,
            lcout => capture_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1697_3_lut_4_lut_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__20059\,
            in1 => \N__29251\,
            in2 => \N__26036\,
            in3 => \N__23868\,
            lcout => \tok.table_wr_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_176_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__22016\,
            in1 => \N__29394\,
            in2 => \N__20069\,
            in3 => \N__17660\,
            lcout => OPEN,
            ltout => \tok.n18_adj_844_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_180_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__24067\,
            in1 => \N__17186\,
            in2 => \N__16874\,
            in3 => \N__21060\,
            lcout => OPEN,
            ltout => \tok.n20_adj_846_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_181_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__16871\,
            in1 => \N__17488\,
            in2 => \N__16859\,
            in3 => \N__17216\,
            lcout => \tok.A_15_N_113_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_3_lut_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__29850\,
            in1 => \_gnd_net_\,
            in2 => \N__19970\,
            in3 => \N__24712\,
            lcout => \tok.n15_adj_847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_175_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101010000"
        )
    port map (
            in0 => \N__27046\,
            in1 => \N__26791\,
            in2 => \N__17210\,
            in3 => \N__29849\,
            lcout => \tok.n12_adj_843\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i0_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17173\,
            in1 => \N__22122\,
            in2 => \_gnd_net_\,
            in3 => \N__17156\,
            lcout => uart_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_adj_82_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__27217\,
            in1 => \N__17144\,
            in2 => \_gnd_net_\,
            in3 => \N__20411\,
            lcout => \tok.n16_adj_730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_155_i16_2_lut_3_lut_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__28075\,
            in1 => \N__29221\,
            in2 => \_gnd_net_\,
            in3 => \N__28117\,
            lcout => \tok.n400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2649_3_lut_4_lut_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__27216\,
            in1 => \N__17036\,
            in2 => \N__29267\,
            in3 => \N__23865\,
            lcout => \tok.n2724\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1771_3_lut_4_lut_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__23866\,
            in1 => \N__18677\,
            in2 => \N__29576\,
            in3 => \N__29226\,
            lcout => \tok.table_wr_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2562_3_lut_4_lut_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110110000"
        )
    port map (
            in0 => \N__24622\,
            in1 => \N__28076\,
            in2 => \N__29266\,
            in3 => \N__26410\,
            lcout => \tok.n2614\,
            ltout => \tok.n2614_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2564_3_lut_4_lut_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__28130\,
            in1 => \N__29222\,
            in2 => \N__17030\,
            in3 => \N__28118\,
            lcout => \tok.n2616\,
            ltout => \tok.n2616_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_186_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__20162\,
            in1 => \N__22028\,
            in2 => \N__17585\,
            in3 => \N__17582\,
            lcout => \tok.n12_adj_851\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_185_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__17564\,
            in1 => \N__20078\,
            in2 => \_gnd_net_\,
            in3 => \N__27215\,
            lcout => \tok.n8_adj_850\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A__15__I_16_i5_3_lut_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27392\,
            in1 => \N__17736\,
            in2 => \_gnd_net_\,
            in3 => \N__17411\,
            lcout => \tok.A_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_163_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__23018\,
            in1 => \N__24278\,
            in2 => \N__17519\,
            in3 => \N__17606\,
            lcout => \tok.A_15_N_113_4\,
            ltout => \tok.A_15_N_113_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i5_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__17348\,
            in1 => \_gnd_net_\,
            in2 => \N__17405\,
            in3 => \N__24394\,
            lcout => \tok.A_low_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26265\,
            ce => \N__17239\,
            sr => \N__19130\
        );

    \tok.i4681_2_lut_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__17737\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17346\,
            lcout => \tok.n950\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17347\,
            in1 => \N__29572\,
            in2 => \_gnd_net_\,
            in3 => \N__17402\,
            lcout => \tok.A_low_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26265\,
            ce => \N__17239\,
            sr => \N__19130\
        );

    \tok.A_i7_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21323\,
            in1 => \N__17349\,
            in2 => \_gnd_net_\,
            in3 => \N__17396\,
            lcout => \tok.A_low_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26265\,
            ce => \N__17239\,
            sr => \N__19130\
        );

    \tok.A_i4_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__17693\,
            in1 => \_gnd_net_\,
            in2 => \N__17374\,
            in3 => \N__21546\,
            lcout => \tok.A_low_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26265\,
            ce => \N__17239\,
            sr => \N__19130\
        );

    \tok.A__15__I_16_i4_3_lut_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17735\,
            in1 => \N__17692\,
            in2 => \_gnd_net_\,
            in3 => \N__21796\,
            lcout => \tok.A_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4375_4_lut_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27228\,
            in1 => \N__26485\,
            in2 => \N__26597\,
            in3 => \N__24268\,
            lcout => OPEN,
            ltout => \tok.n4528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001111"
        )
    port map (
            in0 => \N__29278\,
            in1 => \N__27713\,
            in2 => \N__17678\,
            in3 => \N__17651\,
            lcout => \tok.n892\,
            ltout => \tok.n892_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_174_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011101"
        )
    port map (
            in0 => \N__26562\,
            in1 => \N__21989\,
            in2 => \N__17675\,
            in3 => \N__17672\,
            lcout => \tok.n13_adj_842\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_adj_165_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100110011"
        )
    port map (
            in0 => \N__29820\,
            in1 => \N__24456\,
            in2 => \N__24621\,
            in3 => \N__27986\,
            lcout => \tok.n8_adj_666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_1_lut_2_lut_4_lut_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__30390\,
            in1 => \N__29819\,
            in2 => \N__28013\,
            in3 => \N__30111\,
            lcout => \tok.n8_adj_777\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i54_3_lut_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27423\,
            in1 => \N__26563\,
            in2 => \_gnd_net_\,
            in3 => \N__17888\,
            lcout => OPEN,
            ltout => \tok.n4502_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_159_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100111111"
        )
    port map (
            in0 => \N__26919\,
            in1 => \N__26814\,
            in2 => \N__17609\,
            in3 => \N__29036\,
            lcout => \tok.n12_adj_830\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4678_4_lut_4_lut_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000111111"
        )
    port map (
            in0 => \N__30112\,
            in1 => \N__27987\,
            in2 => \N__29864\,
            in3 => \N__30391\,
            lcout => \tok.n4607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_11_i9_2_lut_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20870\,
            in2 => \_gnd_net_\,
            in3 => \N__29421\,
            lcout => \tok.n9_adj_689\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_99_i9_2_lut_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28324\,
            in2 => \_gnd_net_\,
            in3 => \N__27399\,
            lcout => OPEN,
            ltout => \tok.n181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_35_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__24844\,
            in1 => \N__17893\,
            in2 => \N__17963\,
            in3 => \N__26796\,
            lcout => OPEN,
            ltout => \tok.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__28283\,
            in1 => \N__21813\,
            in2 => \N__17960\,
            in3 => \N__24725\,
            lcout => OPEN,
            ltout => \tok.n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4670_4_lut_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__17957\,
            in1 => \N__21560\,
            in2 => \N__17948\,
            in3 => \N__17945\,
            lcout => \tok.n4684\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_99_i13_2_lut_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28323\,
            in2 => \_gnd_net_\,
            in3 => \N__24843\,
            lcout => OPEN,
            ltout => \tok.n177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_61_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__22994\,
            in1 => \N__17892\,
            in2 => \N__17834\,
            in3 => \N__26795\,
            lcout => OPEN,
            ltout => \tok.n12_adj_696_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_64_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__19826\,
            in1 => \N__27323\,
            in2 => \N__17831\,
            in3 => \N__24724\,
            lcout => \tok.n20_adj_700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_2_lut_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__17786\,
            in1 => \N__17785\,
            in2 => \N__19405\,
            in3 => \N__17753\,
            lcout => \tok.n33_adj_663\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \tok.n3888\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_3_lut_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__18407\,
            in1 => \N__18406\,
            in2 => \N__19430\,
            in3 => \N__18368\,
            lcout => \tok.n33_adj_841\,
            ltout => OPEN,
            carryin => \tok.n3888\,
            carryout => \tok.n3889\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_4_lut_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__18333\,
            in1 => \N__18332\,
            in2 => \N__19406\,
            in3 => \N__18299\,
            lcout => \tok.n33_adj_665\,
            ltout => OPEN,
            carryin => \tok.n3889\,
            carryout => \tok.n3890\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_5_lut_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__18263\,
            in1 => \N__18262\,
            in2 => \N__19431\,
            in3 => \N__18224\,
            lcout => \tok.n33_adj_755\,
            ltout => OPEN,
            carryin => \tok.n3890\,
            carryout => \tok.n3891\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_6_lut_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__18213\,
            in1 => \N__18212\,
            in2 => \N__19407\,
            in3 => \N__18140\,
            lcout => \tok.n33_adj_852\,
            ltout => OPEN,
            carryin => \tok.n3891\,
            carryout => \tok.n3892\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_7_lut_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__18113\,
            in1 => \N__18112\,
            in2 => \N__19432\,
            in3 => \N__18074\,
            lcout => \tok.n33_adj_817\,
            ltout => OPEN,
            carryin => \tok.n3892\,
            carryout => \tok.n3893\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_8_lut_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19214\,
            in1 => \N__19215\,
            in2 => \N__19408\,
            in3 => \N__18071\,
            lcout => \tok.n33\,
            ltout => OPEN,
            carryin => \tok.n3893\,
            carryout => \tok.n3894\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_9_lut_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__18044\,
            in1 => \N__18045\,
            in2 => \N__19433\,
            in3 => \N__18002\,
            lcout => \tok.n33_adj_643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i12_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25708\,
            in1 => \N__17990\,
            in2 => \_gnd_net_\,
            in3 => \N__25327\,
            lcout => \tok.tail_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26231\,
            ce => \N__25471\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i18_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25751\,
            in1 => \N__18536\,
            in2 => \_gnd_net_\,
            in3 => \N__25714\,
            lcout => \tok.C_stk.tail_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26231\,
            ce => \N__25471\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i15_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25709\,
            in1 => \N__22838\,
            in2 => \_gnd_net_\,
            in3 => \N__18562\,
            lcout => \tok.tail_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26231\,
            ce => \N__25471\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i0_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22874\,
            in1 => \N__25712\,
            in2 => \_gnd_net_\,
            in3 => \N__18604\,
            lcout => \tok.C_stk.tail_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26231\,
            ce => \N__25471\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i7_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25711\,
            in1 => \_gnd_net_\,
            in2 => \N__22855\,
            in3 => \N__18746\,
            lcout => \tok.C_stk.tail_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26231\,
            ce => \N__25471\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i4_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18524\,
            in1 => \N__25713\,
            in2 => \_gnd_net_\,
            in3 => \N__30538\,
            lcout => \tok.C_stk.tail_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26231\,
            ce => \N__25471\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i44_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25710\,
            in1 => \N__23231\,
            in2 => \_gnd_net_\,
            in3 => \N__18511\,
            lcout => \tok.tail_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26231\,
            ce => \N__25471\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i48_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18500\,
            in1 => \N__18481\,
            in2 => \_gnd_net_\,
            in3 => \N__25715\,
            lcout => \tok.tail_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26231\,
            ce => \N__25471\,
            sr => \_gnd_net_\
        );

    \tok.i4634_2_lut_3_lut_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18449\,
            in1 => \N__29035\,
            in2 => \_gnd_net_\,
            in3 => \N__29857\,
            lcout => OPEN,
            ltout => \tok.n4694_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__18572\,
            in1 => \N__28549\,
            in2 => \N__18440\,
            in3 => \N__30161\,
            lcout => OPEN,
            ltout => \tok.n13_adj_713_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_71_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__18672\,
            in1 => \N__25251\,
            in2 => \N__18611\,
            in3 => \N__25191\,
            lcout => n10_adj_875,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.n602_bdd_4_lut_4739_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__25106\,
            in1 => \N__26347\,
            in2 => \N__19469\,
            in3 => \N__18673\,
            lcout => OPEN,
            ltout => \tok.C_stk.n4894_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i0_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__26348\,
            in1 => \N__22888\,
            in2 => \N__18608\,
            in3 => \N__18602\,
            lcout => \tok.c_stk_r_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i4666_4_lut_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__26695\,
            in1 => \N__18671\,
            in2 => \N__18605\,
            in3 => \N__25996\,
            lcout => OPEN,
            ltout => \tok.ram.n4717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5_4_lut_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__18603\,
            in1 => \N__25884\,
            in2 => \N__18575\,
            in3 => \N__29856\,
            lcout => \tok.n1_adj_712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.n602_bdd_4_lut_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__18879\,
            in1 => \N__25101\,
            in2 => \N__18845\,
            in3 => \N__26359\,
            lcout => OPEN,
            ltout => \tok.C_stk.n4912_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i7_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__26360\,
            in1 => \N__18566\,
            in2 => \N__18551\,
            in3 => \N__18743\,
            lcout => \tok.c_stk_r_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_137_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18803\,
            in1 => \N__23518\,
            in2 => \_gnd_net_\,
            in3 => \N__18814\,
            lcout => \tok.tc_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i4637_4_lut_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__26694\,
            in1 => \N__25995\,
            in2 => \N__18745\,
            in3 => \N__18878\,
            lcout => OPEN,
            ltout => \tok.ram.n4696_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5_4_lut_adj_26_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__25873\,
            in1 => \N__18739\,
            in2 => \N__18710\,
            in3 => \N__29873\,
            lcout => OPEN,
            ltout => \tok.n1_adj_798_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_132_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__18707\,
            in1 => \N__28531\,
            in2 => \N__18701\,
            in3 => \N__30160\,
            lcout => \tok.n13_adj_799\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_148_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19468\,
            in1 => \N__19480\,
            in2 => \_gnd_net_\,
            in3 => \N__23517\,
            lcout => \tok.tc_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_2_lut_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19454\,
            in2 => \_gnd_net_\,
            in3 => \N__18653\,
            lcout => \tok.tc_plus_1_0\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \tok.n3895\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_3_lut_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18764\,
            in2 => \_gnd_net_\,
            in3 => \N__18626\,
            lcout => \tok.tc_plus_1_1\,
            ltout => OPEN,
            carryin => \tok.n3895\,
            carryout => \tok.n3896\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_4_lut_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25034\,
            in2 => \_gnd_net_\,
            in3 => \N__18623\,
            lcout => \tok.tc_plus_1_2\,
            ltout => OPEN,
            carryin => \tok.n3896\,
            carryout => \tok.n3897\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_5_lut_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23555\,
            in2 => \_gnd_net_\,
            in3 => \N__18620\,
            lcout => \tok.tc_plus_1_3\,
            ltout => OPEN,
            carryin => \tok.n3897\,
            carryout => \tok.n3898\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_6_lut_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25352\,
            in2 => \_gnd_net_\,
            in3 => \N__18617\,
            lcout => \tok.tc_plus_1_4\,
            ltout => OPEN,
            carryin => \tok.n3898\,
            carryout => \tok.n3899\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_7_lut_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23684\,
            in2 => \_gnd_net_\,
            in3 => \N__18614\,
            lcout => \tok.tc_plus_1_5\,
            ltout => OPEN,
            carryin => \tok.n3899\,
            carryout => \tok.n3900\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_8_lut_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18794\,
            in2 => \_gnd_net_\,
            in3 => \N__18896\,
            lcout => \tok.tc_plus_1_6\,
            ltout => OPEN,
            carryin => \tok.n3900\,
            carryout => \tok.n3901\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_9_lut_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18836\,
            in2 => \_gnd_net_\,
            in3 => \N__18893\,
            lcout => \tok.tc_plus_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i7_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23502\,
            in1 => \N__18860\,
            in2 => \_gnd_net_\,
            in3 => \N__18841\,
            lcout => \c_stk_w_7_N_18_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26252\,
            ce => 'H',
            sr => \N__19151\
        );

    \tok.tc_i6_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18801\,
            in1 => \N__23505\,
            in2 => \_gnd_net_\,
            in3 => \N__18815\,
            lcout => \c_stk_w_7_N_18_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26252\,
            ce => 'H',
            sr => \N__19151\
        );

    \tok.tc_i5_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23501\,
            in1 => \N__23711\,
            in2 => \_gnd_net_\,
            in3 => \N__23691\,
            lcout => \c_stk_w_7_N_18_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26252\,
            ce => 'H',
            sr => \N__19151\
        );

    \tok.tc_i4_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25151\,
            in1 => \N__25359\,
            in2 => \_gnd_net_\,
            in3 => \N__23506\,
            lcout => \c_stk_w_7_N_18_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26252\,
            ce => 'H',
            sr => \N__19151\
        );

    \tok.tc_i3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23500\,
            in1 => \_gnd_net_\,
            in2 => \N__23585\,
            in3 => \N__23562\,
            lcout => \c_stk_w_7_N_18_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26252\,
            ce => 'H',
            sr => \N__19151\
        );

    \tok.tc_i2_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23654\,
            in1 => \N__23504\,
            in2 => \_gnd_net_\,
            in3 => \N__25041\,
            lcout => \c_stk_w_7_N_18_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26252\,
            ce => 'H',
            sr => \N__19151\
        );

    \tok.tc_i1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23499\,
            in1 => \N__18773\,
            in2 => \_gnd_net_\,
            in3 => \N__18767\,
            lcout => \c_stk_w_7_N_18_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26252\,
            ce => 'H',
            sr => \N__19151\
        );

    \tok.tc_i0_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19484\,
            in1 => \N__23503\,
            in2 => \_gnd_net_\,
            in3 => \N__19461\,
            lcout => \c_stk_w_7_N_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26252\,
            ce => 'H',
            sr => \N__19151\
        );

    \tok.i1_2_lut_adj_37_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__22261\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19377\,
            lcout => \tok.n5_adj_655\,
            ltout => \tok.n5_adj_655_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_38_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010111011"
        )
    port map (
            in0 => \N__19005\,
            in1 => \N__18989\,
            in2 => \N__19349\,
            in3 => \N__22450\,
            lcout => \stall_\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_105_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101111"
        )
    port map (
            in0 => \N__19346\,
            in1 => \N__24066\,
            in2 => \N__19312\,
            in3 => \N__27050\,
            lcout => \tok.uart_stall\,
            ltout => \tok.uart_stall_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2655_2_lut_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19283\,
            in3 => \N__18990\,
            lcout => \tok.n2732\,
            ltout => \tok.n2732_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i6_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__19184\,
            in1 => \N__18940\,
            in2 => \N__19232\,
            in3 => \N__22748\,
            lcout => \tok.n43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26257\,
            ce => 'H',
            sr => \N__19143\
        );

    \tok.stall_200_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100001101"
        )
    port map (
            in0 => \N__22451\,
            in1 => \N__19157\,
            in2 => \N__18995\,
            in3 => \N__19007\,
            lcout => \tok.stall\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26257\,
            ce => 'H',
            sr => \N__19143\
        );

    \tok.i1_4_lut_adj_179_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__19006\,
            in1 => \N__22262\,
            in2 => \N__22489\,
            in3 => \N__18991\,
            lcout => \tok.n4431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_2_lut_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26900\,
            in2 => \N__29574\,
            in3 => \N__27661\,
            lcout => \tok.n5_adj_682\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \tok.n3925\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_3_lut_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27660\,
            in1 => \N__24173\,
            in2 => \N__20169\,
            in3 => \N__20072\,
            lcout => \tok.n4_adj_790\,
            ltout => OPEN,
            carryin => \tok.n3925\,
            carryout => \tok.n3926\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_4_lut_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27667\,
            in1 => \N__21981\,
            in2 => \N__20060\,
            in3 => \N__19961\,
            lcout => \tok.n5_adj_789\,
            ltout => OPEN,
            carryin => \tok.n3926\,
            carryout => \tok.n3927\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_5_lut_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27657\,
            in1 => \N__21824\,
            in2 => \N__21544\,
            in3 => \N__19958\,
            lcout => \tok.n23_adj_788\,
            ltout => OPEN,
            carryin => \tok.n3927\,
            carryout => \tok.n3928\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_6_lut_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27666\,
            in1 => \N__27411\,
            in2 => \N__24389\,
            in3 => \N__19955\,
            lcout => \tok.n13_adj_787\,
            ltout => OPEN,
            carryin => \tok.n3928\,
            carryout => \tok.n3929\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_7_lut_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27659\,
            in1 => \N__22389\,
            in2 => \N__19951\,
            in3 => \N__19844\,
            lcout => \tok.n5_adj_775\,
            ltout => OPEN,
            carryin => \tok.n3929\,
            carryout => \tok.n3930\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_8_lut_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27668\,
            in1 => \N__28232\,
            in2 => \N__21321\,
            in3 => \N__19829\,
            lcout => \tok.n5_adj_773\,
            ltout => OPEN,
            carryin => \tok.n3930\,
            carryout => \tok.n3931\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_9_lut_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27658\,
            in1 => \N__19775\,
            in2 => \N__19678\,
            in3 => \N__19574\,
            lcout => \tok.n5_adj_752\,
            ltout => OPEN,
            carryin => \tok.n3931\,
            carryout => \tok.n3932\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_10_lut_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27653\,
            in1 => \N__19562\,
            in2 => \N__24856\,
            in3 => \N__19487\,
            lcout => \tok.n5\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \tok.n3933\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_11_lut_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27664\,
            in1 => \N__22656\,
            in2 => \N__21182\,
            in3 => \N__21071\,
            lcout => \tok.n21\,
            ltout => OPEN,
            carryin => \tok.n3933\,
            carryout => \tok.n3934\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_12_lut_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27656\,
            in1 => \N__21055\,
            in2 => \N__20965\,
            in3 => \N__20873\,
            lcout => \tok.n5_adj_668\,
            ltout => OPEN,
            carryin => \tok.n3934\,
            carryout => \tok.n3935\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_13_lut_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27663\,
            in1 => \N__21434\,
            in2 => \N__20869\,
            in3 => \N__20765\,
            lcout => \tok.n5_adj_690\,
            ltout => OPEN,
            carryin => \tok.n3935\,
            carryout => \tok.n3936\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_14_lut_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27654\,
            in1 => \N__23005\,
            in2 => \N__20760\,
            in3 => \N__20684\,
            lcout => \tok.n5_adj_694\,
            ltout => OPEN,
            carryin => \tok.n3936\,
            carryout => \tok.n3937\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_15_lut_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27665\,
            in1 => \N__20676\,
            in2 => \N__20595\,
            in3 => \N__20513\,
            lcout => \tok.n5_adj_710\,
            ltout => OPEN,
            carryin => \tok.n3937\,
            carryout => \tok.n3938\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_16_lut_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27655\,
            in1 => \N__20510\,
            in2 => \N__24014\,
            in3 => \N__20405\,
            lcout => \tok.n5_adj_729\,
            ltout => OPEN,
            carryin => \tok.n3938\,
            carryout => \tok.n3939\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_17_lut_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__27662\,
            in1 => \N__20399\,
            in2 => \N__20321\,
            in3 => \N__20216\,
            lcout => \tok.n5_adj_750\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_167_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20198\,
            in2 => \_gnd_net_\,
            in3 => \N__20183\,
            lcout => OPEN,
            ltout => \tok.n5_adj_837_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_168_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010100"
        )
    port map (
            in0 => \N__29293\,
            in1 => \N__21347\,
            in2 => \N__21554\,
            in3 => \N__22004\,
            lcout => OPEN,
            ltout => \tok.n10_adj_838_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_170_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__21545\,
            in1 => \N__21461\,
            in2 => \N__21452\,
            in3 => \N__29392\,
            lcout => \tok.n12_adj_840\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_166_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__27781\,
            in1 => \N__21435\,
            in2 => \N__21194\,
            in3 => \N__27571\,
            lcout => \tok.n6_adj_835\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_99_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29292\,
            in2 => \_gnd_net_\,
            in3 => \N__27780\,
            lcout => \tok.n109\,
            ltout => \tok.n109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_120_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001100"
        )
    port map (
            in0 => \N__29393\,
            in1 => \N__21341\,
            in2 => \N__21326\,
            in3 => \N__21319\,
            lcout => \tok.n18_adj_782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_102_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27570\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29294\,
            lcout => \tok.n101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i3_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21193\,
            in1 => \N__21221\,
            in2 => \_gnd_net_\,
            in3 => \N__22123\,
            lcout => uart_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_2_lut_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__30322\,
            in1 => \N__30020\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n40\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \tok.n3902\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_3_lut_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__22176\,
            in1 => \N__30323\,
            in2 => \_gnd_net_\,
            in3 => \N__22019\,
            lcout => \tok.n13_adj_816\,
            ltout => OPEN,
            carryin => \tok.n3902\,
            carryout => \tok.n3903\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_4_lut_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__22177\,
            in1 => \N__29824\,
            in2 => \_gnd_net_\,
            in3 => \N__22007\,
            lcout => \tok.n2_adj_811\,
            ltout => OPEN,
            carryin => \tok.n3903\,
            carryout => \tok.n3904\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_5_lut_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__22175\,
            in1 => \N__27988\,
            in2 => \N__21689\,
            in3 => \N__21998\,
            lcout => \tok.n26_adj_808\,
            ltout => OPEN,
            carryin => \tok.n3904\,
            carryout => \tok.n3905\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_6_lut_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__26882\,
            in1 => \N__28973\,
            in2 => \_gnd_net_\,
            in3 => \N__21995\,
            lcout => \tok.n36\,
            ltout => OPEN,
            carryin => \tok.n3905\,
            carryout => \tok.n3906\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_7_lut_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__24180\,
            in1 => \N__28658\,
            in2 => \_gnd_net_\,
            in3 => \N__21992\,
            lcout => \tok.n211\,
            ltout => OPEN,
            carryin => \tok.n3906\,
            carryout => \tok.n3907\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_8_lut_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21986\,
            in1 => \N__28505\,
            in2 => \N__21691\,
            in3 => \N__21854\,
            lcout => \tok.n210\,
            ltout => OPEN,
            carryin => \tok.n3907\,
            carryout => \tok.n3908\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_9_lut_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21794\,
            in1 => \N__28808\,
            in2 => \N__21690\,
            in3 => \N__21704\,
            lcout => \tok.n209\,
            ltout => OPEN,
            carryin => \tok.n3908\,
            carryout => \tok.n3909\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_10_lut_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21665\,
            in2 => \_gnd_net_\,
            in3 => \N__21563\,
            lcout => \tok.n191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2546_2_lut_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24845\,
            in2 => \_gnd_net_\,
            in3 => \N__26599\,
            lcout => \tok.n2598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_5_i2_2_lut_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__22811\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24471\,
            lcout => \tok.n2_adj_810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4623_3_lut_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__22796\,
            in1 => \N__22787\,
            in2 => \_gnd_net_\,
            in3 => \N__22775\,
            lcout => \tok.n4663\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__22490\,
            in1 => \N__28252\,
            in2 => \N__22283\,
            in3 => \N__22754\,
            lcout => \tok.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i7_1_lut_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28251\,
            lcout => \tok.n296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_13_i2_3_lut_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__24472\,
            in1 => \N__22697\,
            in2 => \_gnd_net_\,
            in3 => \N__22657\,
            lcout => \tok.n2_adj_703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_218_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__22491\,
            in1 => \N__22393\,
            in2 => \N__22281\,
            in3 => \N__22196\,
            lcout => \tok.n27_adj_868\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i25_1_lut_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24469\,
            lcout => \tok.n82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i4_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23057\,
            in1 => \N__22148\,
            in2 => \_gnd_net_\,
            in3 => \N__22124\,
            lcout => uart_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_156_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__23069\,
            in1 => \N__23003\,
            in2 => \_gnd_net_\,
            in3 => \N__27575\,
            lcout => OPEN,
            ltout => \tok.n6_adj_827_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_157_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__23056\,
            in1 => \N__23048\,
            in2 => \N__23033\,
            in3 => \N__27795\,
            lcout => OPEN,
            ltout => \tok.n33_adj_828_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_160_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__23030\,
            in1 => \N__29285\,
            in2 => \N__23021\,
            in3 => \N__24470\,
            lcout => \tok.n11_adj_831\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2462_2_lut_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__23004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26600\,
            lcout => \tok.n2514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i8_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25727\,
            in1 => \N__23180\,
            in2 => \_gnd_net_\,
            in3 => \N__22892\,
            lcout => \tok.tail_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26238\,
            ce => \N__25465\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i16_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22867\,
            in1 => \N__23155\,
            in2 => \_gnd_net_\,
            in3 => \N__25728\,
            lcout => \tok.C_stk.tail_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26238\,
            ce => \N__25465\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i23_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25724\,
            in1 => \N__22820\,
            in2 => \_gnd_net_\,
            in3 => \N__22856\,
            lcout => \tok.C_stk.tail_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26238\,
            ce => \N__25465\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i31_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22831\,
            in1 => \N__23198\,
            in2 => \_gnd_net_\,
            in3 => \N__25730\,
            lcout => \tok.tail_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26238\,
            ce => \N__25465\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i39_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25725\,
            in1 => \N__23189\,
            in2 => \_gnd_net_\,
            in3 => \N__22819\,
            lcout => \tok.C_stk.tail_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26238\,
            ce => \N__25465\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i47_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23290\,
            in1 => \N__23197\,
            in2 => \_gnd_net_\,
            in3 => \N__25731\,
            lcout => \tok.tail_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26238\,
            ce => \N__25465\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i55_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25726\,
            in1 => \N__23270\,
            in2 => \_gnd_net_\,
            in3 => \N__23188\,
            lcout => \tok.tail_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26238\,
            ce => \N__25465\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i24_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23179\,
            in1 => \N__23171\,
            in2 => \_gnd_net_\,
            in3 => \N__25729\,
            lcout => \tok.tail_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26238\,
            ce => \N__25465\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i30_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24974\,
            in1 => \N__23129\,
            in2 => \_gnd_net_\,
            in3 => \N__25620\,
            lcout => \tok.tail_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26243\,
            ce => \N__25466\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i38_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23137\,
            in2 => \N__25706\,
            in3 => \N__23119\,
            lcout => \tok.C_stk.tail_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26243\,
            ce => \N__25466\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i22_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25619\,
            in2 => \N__23141\,
            in3 => \N__24940\,
            lcout => \tok.C_stk.tail_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26243\,
            ce => \N__25466\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i46_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__23128\,
            in1 => \N__23254\,
            in2 => \N__25707\,
            in3 => \_gnd_net_\,
            lcout => \tok.tail_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26243\,
            ce => \N__25466\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i54_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23120\,
            in1 => \N__23242\,
            in2 => \_gnd_net_\,
            in3 => \N__25622\,
            lcout => \tok.tail_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26243\,
            ce => \N__25466\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i6_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24941\,
            in1 => \_gnd_net_\,
            in2 => \N__25704\,
            in3 => \N__23111\,
            lcout => \tok.C_stk.tail_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26243\,
            ce => \N__25466\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i52_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23210\,
            in1 => \N__23348\,
            in2 => \_gnd_net_\,
            in3 => \N__25621\,
            lcout => \tok.tail_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26243\,
            ce => \N__25466\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i10_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__23330\,
            in1 => \N__26374\,
            in2 => \N__25705\,
            in3 => \_gnd_net_\,
            lcout => \tok.tail_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26243\,
            ce => \N__25466\,
            sr => \_gnd_net_\
        );

    \tok.i547_3_lut_4_lut_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010101010"
        )
    port map (
            in0 => \N__25459\,
            in1 => \N__24623\,
            in2 => \N__23312\,
            in3 => \N__28074\,
            lcout => \tok.n602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.i545_2_lut_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23311\,
            in2 => \_gnd_net_\,
            in3 => \N__25458\,
            lcout => \tok.C_stk.n600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i63_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__23266\,
            in1 => \N__25697\,
            in2 => \N__23291\,
            in3 => \N__25464\,
            lcout => \tok.tail_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i62_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__25461\,
            in1 => \N__23255\,
            in2 => \N__25733\,
            in3 => \N__23243\,
            lcout => \tok.tail_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i61_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__25015\,
            in1 => \N__25696\,
            in2 => \N__24995\,
            in3 => \N__25463\,
            lcout => \tok.tail_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i60_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__25460\,
            in1 => \N__23230\,
            in2 => \N__25732\,
            in3 => \N__23209\,
            lcout => \tok.tail_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i59_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__24895\,
            in1 => \N__25695\,
            in2 => \N__24875\,
            in3 => \N__25462\,
            lcout => \tok.tail_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.n602_bdd_4_lut_4744_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__25074\,
            in1 => \N__26304\,
            in2 => \N__23699\,
            in3 => \N__23373\,
            lcout => OPEN,
            ltout => \tok.C_stk.n4900_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i5_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__26305\,
            in1 => \N__24560\,
            in2 => \N__23438\,
            in3 => \N__24584\,
            lcout => \tok.c_stk_r_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_98_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__24583\,
            in1 => \N__30380\,
            in2 => \N__23435\,
            in3 => \N__30151\,
            lcout => OPEN,
            ltout => \tok.n83_adj_742_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4619_2_lut_3_lut_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28962\,
            in2 => \N__23402\,
            in3 => \N__29800\,
            lcout => OPEN,
            ltout => \tok.n4651_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_100_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__23393\,
            in1 => \N__28504\,
            in2 => \N__23399\,
            in3 => \N__30152\,
            lcout => \tok.n13_adj_758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.n602_bdd_4_lut_4729_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__26303\,
            in1 => \N__25073\,
            in2 => \N__23570\,
            in3 => \N__23615\,
            lcout => \tok.C_stk.n4882\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i4645_4_lut_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__26683\,
            in1 => \N__25994\,
            in2 => \N__24589\,
            in3 => \N__23372\,
            lcout => OPEN,
            ltout => \tok.ram.n4702_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5_4_lut_adj_24_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__24585\,
            in1 => \N__25899\,
            in2 => \N__23396\,
            in3 => \N__29799\,
            lcout => \tok.n1_adj_757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i4654_4_lut_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__26650\,
            in1 => \N__23619\,
            in2 => \N__30489\,
            in3 => \N__25978\,
            lcout => \tok.ram.n4708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_101_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__25265\,
            in1 => \N__25204\,
            in2 => \N__23387\,
            in3 => \N__23717\,
            lcout => n10_adj_873,
            ltout => \n10_adj_873_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_138_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23521\,
            in1 => \_gnd_net_\,
            in2 => \N__23702\,
            in3 => \N__23692\,
            lcout => \tok.tc_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_81_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__25916\,
            in1 => \N__25203\,
            in2 => \N__25275\,
            in3 => \N__26032\,
            lcout => n10_adj_874,
            ltout => \n10_adj_874_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_143_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23520\,
            in1 => \_gnd_net_\,
            in2 => \N__23642\,
            in3 => \N__25043\,
            lcout => \tok.tc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_88_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23620\,
            in1 => \N__25205\,
            in2 => \N__25276\,
            in3 => \N__25832\,
            lcout => n92_adj_870,
            ltout => \n92_adj_870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_141_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23519\,
            in1 => \_gnd_net_\,
            in2 => \N__23573\,
            in3 => \N__23563\,
            lcout => \tok.tc_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_139_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25144\,
            in1 => \N__25363\,
            in2 => \_gnd_net_\,
            in3 => \N__23522\,
            lcout => \tok.tc_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_113_i9_2_lut_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30286\,
            in2 => \_gnd_net_\,
            in3 => \N__29968\,
            lcout => \tok.n9_adj_645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_220_i11_2_lut_4_lut_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__30288\,
            in1 => \N__29683\,
            in2 => \N__30040\,
            in3 => \N__27884\,
            lcout => \tok.n11_adj_648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_142_i14_2_lut_3_lut_4_lut_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__28400\,
            in1 => \N__28590\,
            in2 => \N__28773\,
            in3 => \N__28904\,
            lcout => \tok.n14_adj_650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_119_i10_2_lut_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29681\,
            in2 => \_gnd_net_\,
            in3 => \N__27880\,
            lcout => \tok.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_120_i14_2_lut_3_lut_4_lut_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__28402\,
            in1 => \N__28594\,
            in2 => \N__28774\,
            in3 => \N__28905\,
            lcout => \tok.n14_adj_702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_121_i9_2_lut_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__30287\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29967\,
            lcout => \tok.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4403_3_lut_4_lut_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110111"
        )
    port map (
            in0 => \N__29682\,
            in1 => \N__29969\,
            in2 => \N__27927\,
            in3 => \_gnd_net_\,
            lcout => \tok.n4558\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__28903\,
            in1 => \N__28739\,
            in2 => \N__28625\,
            in3 => \N__28401\,
            lcout => \tok.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_119_i11_2_lut_4_lut_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__29674\,
            in1 => \N__30279\,
            in2 => \N__27923\,
            in3 => \N__29962\,
            lcout => \tok.n11_adj_647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_1_lut_2_lut_4_lut_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__29966\,
            in1 => \N__27879\,
            in2 => \N__30345\,
            in3 => \N__29680\,
            lcout => \tok.n9_adj_797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4315_2_lut_4_lut_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__29679\,
            in1 => \N__30282\,
            in2 => \N__27926\,
            in3 => \N__29965\,
            lcout => \tok.n4464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2534_2_lut_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29676\,
            in2 => \_gnd_net_\,
            in3 => \N__27868\,
            lcout => \tok.n2586\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_121_i11_2_lut_4_lut_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__29677\,
            in1 => \N__30280\,
            in2 => \N__27924\,
            in3 => \N__29963\,
            lcout => \tok.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_4_lut_adj_154_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__28906\,
            in1 => \N__28746\,
            in2 => \N__28634\,
            in3 => \N__28416\,
            lcout => \tok.n14_adj_825\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_114_i11_2_lut_4_lut_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__29678\,
            in1 => \N__30281\,
            in2 => \N__27925\,
            in3 => \N__29964\,
            lcout => \tok.n11_adj_649\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_123_i10_2_lut_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27869\,
            in2 => \_gnd_net_\,
            in3 => \N__29675\,
            lcout => \tok.n10_adj_646\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4417_4_lut_4_lut_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111010101"
        )
    port map (
            in0 => \N__30289\,
            in1 => \N__29684\,
            in2 => \N__27928\,
            in3 => \N__29973\,
            lcout => OPEN,
            ltout => \tok.n4575_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_32_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110111111"
        )
    port map (
            in0 => \N__23773\,
            in1 => \N__23801\,
            in2 => \N__23780\,
            in3 => \N__27266\,
            lcout => \tok.n4424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4373_4_lut_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111011"
        )
    port map (
            in0 => \N__23756\,
            in1 => \N__26441\,
            in2 => \N__27596\,
            in3 => \N__27500\,
            lcout => \tok.n83\,
            ltout => \tok.n83_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2669_2_lut_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__26730\,
            in1 => \_gnd_net_\,
            in2 => \N__23777\,
            in3 => \_gnd_net_\,
            lcout => \tok.n2746\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4413_4_lut_4_lut_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111110011"
        )
    port map (
            in0 => \N__30291\,
            in1 => \N__29685\,
            in2 => \N__27930\,
            in3 => \N__29974\,
            lcout => OPEN,
            ltout => \tok.n4571_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_34_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100111111"
        )
    port map (
            in0 => \N__23774\,
            in1 => \N__29121\,
            in2 => \N__23759\,
            in3 => \N__28056\,
            lcout => \tok.n4393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_3_lut_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110101"
        )
    port map (
            in0 => \N__30290\,
            in1 => \_gnd_net_\,
            in2 => \N__27929\,
            in3 => \N__29975\,
            lcout => OPEN,
            ltout => \tok.n4460_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2651_4_lut_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__27289\,
            in1 => \N__29122\,
            in2 => \N__24500\,
            in3 => \N__26455\,
            lcout => \tok.n2726\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_158_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__24659\,
            in1 => \N__29436\,
            in2 => \N__24393\,
            in3 => \N__28971\,
            lcout => OPEN,
            ltout => \tok.n10_adj_829_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_162_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__30571\,
            in1 => \N__24293\,
            in2 => \N__24281\,
            in3 => \N__27188\,
            lcout => \tok.n13_adj_833\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_169_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__28001\,
            in1 => \N__30184\,
            in2 => \N__27218\,
            in3 => \N__24261\,
            lcout => \tok.n8_adj_839\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_55_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__24068\,
            in1 => \N__24857\,
            in2 => \N__24226\,
            in3 => \N__27192\,
            lcout => \tok.n18_adj_681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.xor_103_i7_2_lut_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24186\,
            in2 => \_gnd_net_\,
            in3 => \N__28543\,
            lcout => OPEN,
            ltout => \tok.n244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_122_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__24069\,
            in1 => \N__23983\,
            in2 => \N__23912\,
            in3 => \N__24703\,
            lcout => \tok.n17_adj_785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_13_i3_2_lut_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24855\,
            in2 => \_gnd_net_\,
            in3 => \N__24704\,
            lcout => \tok.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_172_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28000\,
            in2 => \_gnd_net_\,
            in3 => \N__29782\,
            lcout => \tok.n40_adj_661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4329_2_lut_3_lut_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__30393\,
            in1 => \N__27530\,
            in2 => \_gnd_net_\,
            in3 => \N__30109\,
            lcout => \tok.n4478\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i13_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24533\,
            in1 => \N__24553\,
            in2 => \_gnd_net_\,
            in3 => \N__25639\,
            lcout => \tok.tail_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26249\,
            ce => \N__25467\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i5_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25638\,
            in1 => \N__24542\,
            in2 => \_gnd_net_\,
            in3 => \N__24590\,
            lcout => \tok.C_stk.tail_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26249\,
            ce => \N__25467\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i21_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24541\,
            in1 => \_gnd_net_\,
            in2 => \N__24524\,
            in3 => \N__25640\,
            lcout => \tok.C_stk.tail_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26249\,
            ce => \N__25467\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i29_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25636\,
            in1 => \N__24532\,
            in2 => \_gnd_net_\,
            in3 => \N__24509\,
            lcout => \tok.tail_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26249\,
            ce => \N__25467\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i37_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24520\,
            in1 => \N__25004\,
            in2 => \_gnd_net_\,
            in3 => \N__25641\,
            lcout => \tok.C_stk.tail_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26249\,
            ce => \N__25467\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i45_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25637\,
            in1 => \N__24985\,
            in2 => \_gnd_net_\,
            in3 => \N__24508\,
            lcout => \tok.tail_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26249\,
            ce => \N__25467\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i53_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25016\,
            in1 => \N__25003\,
            in2 => \_gnd_net_\,
            in3 => \N__25642\,
            lcout => \tok.tail_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26249\,
            ce => \N__25467\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i14_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25635\,
            in1 => \N__24973\,
            in2 => \_gnd_net_\,
            in3 => \N__24952\,
            lcout => \tok.tail_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26249\,
            ce => \N__25467\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i11_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25716\,
            in1 => \N__24923\,
            in2 => \_gnd_net_\,
            in3 => \N__25132\,
            lcout => \tok.tail_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26254\,
            ce => \N__25472\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i3_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24932\,
            in1 => \N__25721\,
            in2 => \_gnd_net_\,
            in3 => \N__30487\,
            lcout => \tok.C_stk.tail_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26254\,
            ce => \N__25472\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i19_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25717\,
            in1 => \N__24914\,
            in2 => \_gnd_net_\,
            in3 => \N__24931\,
            lcout => \tok.C_stk.tail_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26254\,
            ce => \N__25472\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i27_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24922\,
            in1 => \N__24905\,
            in2 => \_gnd_net_\,
            in3 => \N__25722\,
            lcout => \tok.tail_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26254\,
            ce => \N__25472\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i35_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25718\,
            in1 => \N__24884\,
            in2 => \_gnd_net_\,
            in3 => \N__24913\,
            lcout => \tok.C_stk.tail_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26254\,
            ce => \N__25472\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i43_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24868\,
            in1 => \N__24904\,
            in2 => \_gnd_net_\,
            in3 => \N__25723\,
            lcout => \tok.tail_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26254\,
            ce => \N__25472\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i51_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25719\,
            in1 => \N__24896\,
            in2 => \_gnd_net_\,
            in3 => \N__24883\,
            lcout => \tok.tail_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26254\,
            ce => \N__25472\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i2_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25747\,
            in1 => \N__25720\,
            in2 => \_gnd_net_\,
            in3 => \N__25826\,
            lcout => \tok.C_stk.tail_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26254\,
            ce => \N__25472\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.n602_bdd_4_lut_4734_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001011000"
        )
    port map (
            in0 => \N__26322\,
            in1 => \N__25297\,
            in2 => \N__25105\,
            in3 => \N__25364\,
            lcout => OPEN,
            ltout => \tok.C_stk.n4888_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i4_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__25334\,
            in1 => \N__30536\,
            in2 => \N__25316\,
            in3 => \N__26324\,
            lcout => \tok.c_stk_r_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i4650_4_lut_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__26682\,
            in1 => \N__25295\,
            in2 => \N__30539\,
            in3 => \N__26000\,
            lcout => OPEN,
            ltout => \tok.ram.n4705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5_4_lut_adj_23_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__29851\,
            in1 => \N__30535\,
            in2 => \N__25313\,
            in3 => \N__25910\,
            lcout => OPEN,
            ltout => \tok.n1_adj_745_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_92_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__27704\,
            in1 => \N__28556\,
            in2 => \N__25310\,
            in3 => \N__30153\,
            lcout => OPEN,
            ltout => \tok.n13_adj_746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_93_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__25296\,
            in1 => \N__25277\,
            in2 => \N__25208\,
            in3 => \N__25202\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i3_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__26323\,
            in1 => \N__25133\,
            in2 => \N__25121\,
            in3 => \N__30488\,
            lcout => \tok.c_stk_r_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26260\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.n602_bdd_4_lut_4724_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001011000"
        )
    port map (
            in0 => \N__26330\,
            in1 => \N__26031\,
            in2 => \N__25111\,
            in3 => \N__25042\,
            lcout => OPEN,
            ltout => \tok.C_stk.n4876_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i2_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__26378\,
            in1 => \N__25821\,
            in2 => \N__26363\,
            in3 => \N__26331\,
            lcout => \tok.c_stk_r_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i4658_4_lut_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__26673\,
            in1 => \N__26030\,
            in2 => \N__25825\,
            in3 => \N__25979\,
            lcout => OPEN,
            ltout => \tok.ram.n4711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5_4_lut_adj_21_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__25909\,
            in1 => \N__25820\,
            in2 => \N__25922\,
            in3 => \N__29863\,
            lcout => OPEN,
            ltout => \tok.n1_adj_724_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_78_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__25757\,
            in1 => \N__28532\,
            in2 => \N__25919\,
            in3 => \N__30136\,
            lcout => \tok.n13_adj_725\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5_4_lut_adj_22_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__25908\,
            in1 => \N__25844\,
            in2 => \N__30493\,
            in3 => \N__29862\,
            lcout => \tok.n1_adj_736\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i18_4_lut_adj_87_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__30105\,
            in1 => \N__25838\,
            in2 => \N__29606\,
            in3 => \N__28459\,
            lcout => \tok.n5_adj_737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_75_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__30384\,
            in1 => \N__25816\,
            in2 => \N__25796\,
            in3 => \N__30104\,
            lcout => OPEN,
            ltout => \tok.n83_adj_721_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4632_2_lut_3_lut_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__29859\,
            in1 => \_gnd_net_\,
            in2 => \N__25760\,
            in3 => \N__28941\,
            lcout => \tok.n4692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i2_4_lut_4_lut_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__30381\,
            in1 => \N__29858\,
            in2 => \N__28012\,
            in3 => \N__30102\,
            lcout => OPEN,
            ltout => \tok.ram.n14_adj_631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i2581_4_lut_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__26497\,
            in1 => \N__27556\,
            in2 => \N__26819\,
            in3 => \N__28057\,
            lcout => \tok.n2635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_130_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30383\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28940\,
            lcout => \tok.n4_adj_795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_150_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30103\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30382\,
            lcout => \tok.n41\,
            ltout => \tok.n41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_45_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__28058\,
            in1 => \N__29597\,
            in2 => \N__26627\,
            in3 => \N__28939\,
            lcout => \tok.n884\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_157_i15_2_lut_3_lut_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__28055\,
            in1 => \N__28103\,
            in2 => \_gnd_net_\,
            in3 => \N__26498\,
            lcout => \tok.n15_adj_662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4415_4_lut_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__28104\,
            in1 => \N__27528\,
            in2 => \N__26456\,
            in3 => \N__27267\,
            lcout => \tok.n4573\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011111111"
        )
    port map (
            in0 => \N__28102\,
            in1 => \N__28054\,
            in2 => \N__26434\,
            in3 => \N__26397\,
            lcout => OPEN,
            ltout => \tok.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110101"
        )
    port map (
            in0 => \N__27690\,
            in1 => \N__30352\,
            in2 => \N__26381\,
            in3 => \N__30044\,
            lcout => OPEN,
            ltout => \tok.n4422_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_33_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__27589\,
            in1 => \N__27538\,
            in2 => \N__27578\,
            in3 => \N__27555\,
            lcout => OPEN,
            ltout => \tok.n51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_36_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110001"
        )
    port map (
            in0 => \N__27539\,
            in1 => \N__27529\,
            in2 => \N__27509\,
            in3 => \N__27506\,
            lcout => \tok.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_adj_60_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__27494\,
            in1 => \N__27479\,
            in2 => \_gnd_net_\,
            in3 => \N__27168\,
            lcout => OPEN,
            ltout => \tok.n14_adj_695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_62_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__27045\,
            in1 => \N__27470\,
            in2 => \N__27455\,
            in3 => \N__27448\,
            lcout => \tok.n18_adj_698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2458_2_lut_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30412\,
            in2 => \_gnd_net_\,
            in3 => \N__30113\,
            lcout => \tok.n2177\,
            ltout => \tok.n2177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1_3_lut_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27290\,
            in2 => \N__27278\,
            in3 => \N__27268\,
            lcout => \tok.n132\,
            ltout => \tok.n132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27122\,
            in2 => \N__27110\,
            in3 => \N__27107\,
            lcout => \tok.n14_adj_651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101110"
        )
    port map (
            in0 => \N__27098\,
            in1 => \N__27083\,
            in2 => \N__27061\,
            in3 => \N__26933\,
            lcout => \tok.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_99_i11_2_lut_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28299\,
            in2 => \_gnd_net_\,
            in3 => \N__28260\,
            lcout => \tok.n179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_117_i10_2_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__27979\,
            in1 => \N__29802\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n10_adj_675\,
            ltout => \tok.n10_adj_675_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4335_3_lut_4_lut_4_lut_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__27762\,
            in1 => \N__28116\,
            in2 => \N__28079\,
            in3 => \N__28073\,
            lcout => \tok.n4484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_4_lut_adj_152_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__30392\,
            in1 => \N__29801\,
            in2 => \N__28011\,
            in3 => \N__30110\,
            lcout => \tok.n2178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_42_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__27737\,
            in1 => \N__27728\,
            in2 => \N__27722\,
            in3 => \N__27698\,
            lcout => \tok.n42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4585_2_lut_3_lut_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30500\,
            in1 => \N__28990\,
            in2 => \_gnd_net_\,
            in3 => \N__29860\,
            lcout => \tok.n4688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_233_i14_2_lut_3_lut_4_lut_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__28449\,
            in1 => \N__28626\,
            in2 => \N__28807\,
            in3 => \N__28934\,
            lcout => \tok.n14_adj_658\,
            ltout => \tok.n14_adj_658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_154_i16_3_lut_4_lut_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__27691\,
            in1 => \N__30385\,
            in2 => \N__27671\,
            in3 => \N__30106\,
            lcout => \tok.n399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_90_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101001000000"
        )
    port map (
            in0 => \N__30107\,
            in1 => \N__30572\,
            in2 => \N__30418\,
            in3 => \N__30537\,
            lcout => \tok.n83_adj_743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_84_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__30494\,
            in1 => \N__30389\,
            in2 => \N__30194\,
            in3 => \N__30108\,
            lcout => OPEN,
            ltout => \tok.n83_adj_733_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4584_2_lut_3_lut_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28935\,
            in2 => \N__29876\,
            in3 => \N__29861\,
            lcout => \tok.n4627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__28627\,
            in1 => \N__28775\,
            in2 => \_gnd_net_\,
            in3 => \N__28450\,
            lcout => \tok.n883\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_adj_53_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__29591\,
            in1 => \N__29573\,
            in2 => \_gnd_net_\,
            in3 => \N__29457\,
            lcout => \tok.n15_adj_680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4710_2_lut_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29149\,
            in2 => \_gnd_net_\,
            in3 => \N__29126\,
            lcout => \tok.write_flag\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i244_2_lut_3_lut_4_lut_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__28989\,
            in1 => \N__28830\,
            in2 => \N__28699\,
            in3 => \N__28542\,
            lcout => \tok.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
