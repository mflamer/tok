-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Dec 31 2020 17:42:06

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    tx : out std_logic;
    rx : in std_logic;
    reset : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__38690\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13042\ : std_logic;
signal \VCCG0\ : std_logic;
signal \tok.A_stk.tail_73\ : std_logic;
signal \tok.A_stk.tail_93\ : std_logic;
signal \tok.A_stk.tail_77\ : std_logic;
signal \tok.A_stk.tail_61\ : std_logic;
signal \tok.A_stk.tail_45\ : std_logic;
signal \tok.A_stk.tail_29\ : std_logic;
signal \tok.A_stk.tail_13\ : std_logic;
signal \tok.A_stk.tail_75\ : std_logic;
signal \tok.A_stk.tail_59\ : std_logic;
signal \tok.A_stk.tail_43\ : std_logic;
signal \tok.A_stk.tail_27\ : std_logic;
signal \tok.A_stk.tail_85\ : std_logic;
signal \tok.A_stk.tail_69\ : std_logic;
signal \tok.A_stk.tail_53\ : std_logic;
signal \tok.A_stk.tail_37\ : std_logic;
signal \tok.A_stk.tail_21\ : std_logic;
signal \tok.A_stk.tail_5\ : std_logic;
signal \tok.A_stk.tail_11\ : std_logic;
signal \tok.A_stk.tail_9\ : std_logic;
signal \tok.A_stk.tail_25\ : std_logic;
signal \tok.A_stk.tail_57\ : std_logic;
signal \tok.A_stk.tail_41\ : std_logic;
signal \tok.table_rd_10\ : std_logic;
signal \tok.n203_adj_866_cascade_\ : std_logic;
signal \tok.n212_adj_867_cascade_\ : std_logic;
signal \tok.n6426_cascade_\ : std_logic;
signal tail_80 : std_logic;
signal \tok.A_stk.tail_64\ : std_logic;
signal tail_48 : std_logic;
signal \tok.A_stk.tail_32\ : std_logic;
signal tail_16 : std_logic;
signal tail_96 : std_logic;
signal tail_112 : std_logic;
signal tail_118 : std_logic;
signal \tok.table_wr_data_8\ : std_logic;
signal \tok.A_stk.tail_89\ : std_logic;
signal tail_122 : std_logic;
signal tail_106 : std_logic;
signal \tok.A_stk.tail_90\ : std_logic;
signal \tok.A_stk.tail_74\ : std_logic;
signal \tok.A_stk.tail_58\ : std_logic;
signal \tok.A_stk.tail_42\ : std_logic;
signal tail_109 : std_logic;
signal tail_125 : std_logic;
signal \tok.n6274\ : std_logic;
signal \tok.n34_cascade_\ : std_logic;
signal \A_stk_delta_1_cascade_\ : std_logic;
signal tail_105 : std_logic;
signal tail_121 : std_logic;
signal tail_101 : std_logic;
signal tail_117 : std_logic;
signal \tok.n34\ : std_logic;
signal tail_100 : std_logic;
signal \rd_15__N_300_cascade_\ : std_logic;
signal tail_116 : std_logic;
signal \tok.A_stk.tail_91\ : std_logic;
signal tail_123 : std_logic;
signal tail_107 : std_logic;
signal \tok.A_stk.tail_84\ : std_logic;
signal \tok.A_stk.tail_68\ : std_logic;
signal \tok.A_stk.tail_52\ : std_logic;
signal \tok.A_stk.tail_36\ : std_logic;
signal \tok.A_stk.tail_20\ : std_logic;
signal \tok.A_stk.tail_0\ : std_logic;
signal \tok.A_stk.tail_4\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \tok.n4767\ : std_logic;
signal \tok.n4768\ : std_logic;
signal \tok.n4769\ : std_logic;
signal \tok.n4770\ : std_logic;
signal \tok.n4771\ : std_logic;
signal \tok.n4772\ : std_logic;
signal \tok.n4773\ : std_logic;
signal tail_120 : std_logic;
signal tail_104 : std_logic;
signal \tok.A_stk.tail_88\ : std_logic;
signal \tok.A_stk.tail_72\ : std_logic;
signal \tok.A_stk.tail_56\ : std_logic;
signal \tok.A_stk.tail_40\ : std_logic;
signal \tok.A_stk.tail_24\ : std_logic;
signal \tok.A_stk.tail_8\ : std_logic;
signal \tok.table_rd_13\ : std_logic;
signal \tok.n226_cascade_\ : std_logic;
signal \tok.n203_adj_643_cascade_\ : std_logic;
signal \tok.n226\ : std_logic;
signal \tok.n212_adj_646_cascade_\ : std_logic;
signal \tok.n6448_cascade_\ : std_logic;
signal \tok.n6388\ : std_logic;
signal \tok.n206_adj_649\ : std_logic;
signal \tok.table_rd_9\ : std_logic;
signal \tok.n203_adj_833_cascade_\ : std_logic;
signal \tok.n212_adj_835_cascade_\ : std_logic;
signal \tok.n206_adj_834\ : std_logic;
signal \tok.n6443_cascade_\ : std_logic;
signal \tok.n242_adj_839_cascade_\ : std_logic;
signal \tok.n230\ : std_logic;
signal \tok.n242_adj_874\ : std_logic;
signal \tok.n6431_cascade_\ : std_logic;
signal \tok.n206_adj_869\ : std_logic;
signal \tok.n206_adj_691\ : std_logic;
signal \tok.n212_adj_689_cascade_\ : std_logic;
signal \tok.n229_adj_863\ : std_logic;
signal \tok.uart.n6223_cascade_\ : std_logic;
signal \txtick_cascade_\ : std_logic;
signal \tok.uart.n12\ : std_logic;
signal \tok.uart.txclkcounter_0\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \tok.uart.txclkcounter_1\ : std_logic;
signal \tok.uart.n4830\ : std_logic;
signal \tok.uart.txclkcounter_2\ : std_logic;
signal \tok.uart.n4831\ : std_logic;
signal \tok.uart.txclkcounter_3\ : std_logic;
signal \tok.uart.n4832\ : std_logic;
signal \tok.uart.txclkcounter_4\ : std_logic;
signal \tok.uart.n4833\ : std_logic;
signal \tok.uart.txclkcounter_5\ : std_logic;
signal \tok.uart.n4834\ : std_logic;
signal \tok.uart.txclkcounter_6\ : std_logic;
signal \tok.uart.n4835\ : std_logic;
signal \tok.uart.txclkcounter_7\ : std_logic;
signal \tok.uart.n4836\ : std_logic;
signal \tok.uart.n4837\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \tok.uart.txclkcounter_8\ : std_logic;
signal tail_127 : std_logic;
signal tail_111 : std_logic;
signal \tok.A_stk.tail_95\ : std_logic;
signal \tok.A_stk.tail_79\ : std_logic;
signal \tok.A_stk.tail_63\ : std_logic;
signal \tok.A_stk.tail_47\ : std_logic;
signal \tok.A_stk.tail_31\ : std_logic;
signal \tok.A_stk.tail_15\ : std_logic;
signal \tok.A_stk.tail_26\ : std_logic;
signal tail_126 : std_logic;
signal tail_110 : std_logic;
signal \tok.A_stk.tail_94\ : std_logic;
signal \tok.A_stk.tail_78\ : std_logic;
signal \tok.A_stk.tail_62\ : std_logic;
signal \tok.A_stk.tail_46\ : std_logic;
signal \tok.A_stk.tail_30\ : std_logic;
signal \tok.A_stk.tail_14\ : std_logic;
signal \tok.A_stk.tail_34\ : std_logic;
signal \tok.A_stk.tail_50\ : std_logic;
signal \tok.A_stk.tail_66\ : std_logic;
signal \tok.A_stk.tail_82\ : std_logic;
signal table_wr_data_0 : std_logic;
signal tail_98 : std_logic;
signal tail_114 : std_logic;
signal \tok.n4_adj_642_cascade_\ : std_logic;
signal \tok.table_wr_data_13\ : std_logic;
signal \tok.table_wr_data_10\ : std_logic;
signal \tok.table_wr_data_15\ : std_logic;
signal \tok.n33_adj_631\ : std_logic;
signal \tok.n27_cascade_\ : std_logic;
signal \tok.n41\ : std_logic;
signal \tok.n33_adj_662\ : std_logic;
signal \tok.n27_adj_709_cascade_\ : std_logic;
signal \tok.n19\ : std_logic;
signal \tok.n33_adj_634\ : std_logic;
signal \tok.n27_adj_706_cascade_\ : std_logic;
signal \tok.n35\ : std_logic;
signal \tok.n6667_cascade_\ : std_logic;
signal \tok.n2532\ : std_logic;
signal \tok.n4_adj_642\ : std_logic;
signal \tok.found_slot_cascade_\ : std_logic;
signal \tok.write_slot\ : std_logic;
signal \tok.n21_cascade_\ : std_logic;
signal \tok.n30_adj_647\ : std_logic;
signal \tok.key_rd_10\ : std_logic;
signal \tok.key_rd_12\ : std_logic;
signal \tok.n26\ : std_logic;
signal \tok.n27_adj_639_cascade_\ : std_logic;
signal \tok.found_slot_N_144\ : std_logic;
signal \tok.n6322\ : std_logic;
signal \tok.n313_cascade_\ : std_logic;
signal \tok.key_rd_2\ : std_logic;
signal \tok.key_rd_7\ : std_logic;
signal \tok.n22\ : std_logic;
signal \tok.table_rd_12\ : std_logic;
signal \tok.n227\ : std_logic;
signal \tok.n203_cascade_\ : std_logic;
signal \tok.n212_cascade_\ : std_logic;
signal \tok.n206\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \tok.n4774\ : std_logic;
signal \tok.n4775\ : std_logic;
signal \tok.n4776\ : std_logic;
signal \tok.n4777\ : std_logic;
signal \tok.n4778\ : std_logic;
signal \tok.n4779\ : std_logic;
signal \tok.n4780\ : std_logic;
signal \tok.n4781\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \tok.n214_cascade_\ : std_logic;
signal \tok.n6358\ : std_logic;
signal \tok.n6402\ : std_logic;
signal \tok.table_rd_14\ : std_logic;
signal \tok.n225_cascade_\ : std_logic;
signal \tok.n203_adj_664_cascade_\ : std_logic;
signal \tok.n225\ : std_logic;
signal \tok.n224\ : std_logic;
signal \tok.table_rd_15\ : std_logic;
signal \tok.n224_cascade_\ : std_logic;
signal \tok.n203_adj_688\ : std_logic;
signal \tok.n6373_cascade_\ : std_logic;
signal \tok.n206_adj_666_cascade_\ : std_logic;
signal \tok.n212_adj_665\ : std_logic;
signal \tok.n281_cascade_\ : std_logic;
signal \tok.n236_adj_864_cascade_\ : std_logic;
signal \tok.n2648_cascade_\ : std_logic;
signal \tok.n226_adj_865\ : std_logic;
signal \tok.n6334\ : std_logic;
signal \tok.n4_adj_762\ : std_logic;
signal \tok.n6316\ : std_logic;
signal sender_1 : std_logic;
signal tx_c : std_logic;
signal \tok.A_stk.tail_65\ : std_logic;
signal tail_49 : std_logic;
signal tail_81 : std_logic;
signal \tok.A_stk.tail_33\ : std_logic;
signal tail_17 : std_logic;
signal \tok.A_stk.tail_1\ : std_logic;
signal tail_102 : std_logic;
signal \tok.A_stk.tail_86\ : std_logic;
signal \tok.A_stk.tail_70\ : std_logic;
signal \tok.A_stk.tail_54\ : std_logic;
signal \tok.A_stk.tail_38\ : std_logic;
signal \tok.A_stk.tail_22\ : std_logic;
signal \tok.A_stk.tail_28\ : std_logic;
signal \tok.A_stk.tail_44\ : std_logic;
signal \tok.A_stk.tail_92\ : std_logic;
signal \tok.A_stk.tail_60\ : std_logic;
signal \tok.A_stk.tail_76\ : std_logic;
signal \tok.A_stk.tail_6\ : std_logic;
signal \tok.A_stk.tail_12\ : std_logic;
signal \tok.A_stk.tail_10\ : std_logic;
signal \tok.A_stk.tail_83\ : std_logic;
signal \tok.A_stk.tail_67\ : std_logic;
signal \tok.A_stk.tail_51\ : std_logic;
signal \tok.A_stk.tail_35\ : std_logic;
signal \tok.A_stk.tail_19\ : std_logic;
signal \tok.A_stk.tail_3\ : std_logic;
signal \tok.n4_cascade_\ : std_logic;
signal \tok.n6273\ : std_logic;
signal \tok.table_wr_data_9\ : std_logic;
signal \tok.n4\ : std_logic;
signal \tok.n6252\ : std_logic;
signal \tok.n6253_cascade_\ : std_logic;
signal tail_99 : std_logic;
signal tail_115 : std_logic;
signal \tok.n33_adj_633\ : std_logic;
signal \tok.n27_adj_704_cascade_\ : std_logic;
signal \tok.n38\ : std_logic;
signal \tok.n33_adj_632\ : std_logic;
signal \tok.n33_adj_661\ : std_logic;
signal \tok.n27_adj_705_cascade_\ : std_logic;
signal \tok.n36\ : std_logic;
signal \tok.n27_adj_703\ : std_logic;
signal \tok.n40\ : std_logic;
signal \tok.n32\ : std_logic;
signal \tok.n33\ : std_logic;
signal \tok.n27_adj_707\ : std_logic;
signal \tok.n33_adj_663\ : std_logic;
signal \tok.n27_adj_708_cascade_\ : std_logic;
signal \tok.n29\ : std_logic;
signal \tok.search_clk\ : std_logic;
signal \tok.found_slot\ : std_logic;
signal \tok.n6670\ : std_logic;
signal \tok.key_rd_6\ : std_logic;
signal \tok.key_rd_0\ : std_logic;
signal \tok.n25\ : std_logic;
signal \tok.key_rd_4\ : std_logic;
signal \tok.key_rd_1\ : std_logic;
signal \tok.n18\ : std_logic;
signal \tok.n6575_cascade_\ : std_logic;
signal \tok.n177\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \tok.n4797\ : std_logic;
signal \tok.n4798\ : std_logic;
signal \tok.n4799\ : std_logic;
signal \tok.n6556\ : std_logic;
signal \tok.n4800\ : std_logic;
signal \tok.n4801\ : std_logic;
signal \tok.n4802\ : std_logic;
signal \tok.n4803\ : std_logic;
signal \tok.n4803_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \tok.n4804\ : std_logic;
signal \tok.n6437\ : std_logic;
signal \tok.n4805\ : std_logic;
signal \tok.n4806\ : std_logic;
signal \tok.n4807\ : std_logic;
signal \tok.n4808\ : std_logic;
signal \tok.n6377\ : std_logic;
signal \tok.n4809\ : std_logic;
signal \tok.n4810\ : std_logic;
signal \tok.n4810_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \tok.n4811\ : std_logic;
signal \tok.n6362\ : std_logic;
signal \tok.n83\ : std_logic;
signal \tok.n161_adj_836\ : std_logic;
signal \tok.n197_adj_837_cascade_\ : std_logic;
signal \tok.n248_adj_838\ : std_logic;
signal \tok.n161_adj_650\ : std_logic;
signal \tok.n6386_cascade_\ : std_logic;
signal \tok.n197_adj_652_cascade_\ : std_logic;
signal \tok.table_rd_11\ : std_logic;
signal \tok.n228_cascade_\ : std_logic;
signal \tok.n203_adj_879_cascade_\ : std_logic;
signal \tok.n228\ : std_logic;
signal \tok.n212_adj_880_cascade_\ : std_logic;
signal \tok.n6339\ : std_logic;
signal \tok.n161_adj_692_cascade_\ : std_logic;
signal \tok.n6356\ : std_logic;
signal \tok.n6417\ : std_logic;
signal \tok.n206_adj_881\ : std_logic;
signal \tok.n6412\ : std_logic;
signal tail_119 : std_logic;
signal tail_103 : std_logic;
signal \tok.A_stk.tail_87\ : std_logic;
signal \tok.A_stk.tail_71\ : std_logic;
signal \tok.A_stk.tail_55\ : std_logic;
signal \tok.A_stk.tail_39\ : std_logic;
signal \tok.A_stk.tail_23\ : std_logic;
signal \tok.A_stk.tail_7\ : std_logic;
signal tail_97 : std_logic;
signal tail_113 : std_logic;
signal tail_108 : std_logic;
signal tail_124 : std_logic;
signal \tok.table_wr_data_3\ : std_logic;
signal table_wr_data_1 : std_logic;
signal \tok.table_wr_data_6\ : std_logic;
signal \tok.table_wr_data_4\ : std_logic;
signal \tok.table_wr_data_2\ : std_logic;
signal \tok.ram.n6266_cascade_\ : std_logic;
signal \tok.n1495_cascade_\ : std_logic;
signal \tok.n13_adj_766\ : std_logic;
signal n10_adj_907 : std_logic;
signal \n10_adj_907_cascade_\ : std_logic;
signal \tok.tc_6\ : std_logic;
signal \tok.n83_adj_765_cascade_\ : std_logic;
signal \tok.n6435\ : std_logic;
signal \tok.n6283_cascade_\ : std_logic;
signal \tok.n80_cascade_\ : std_logic;
signal \tok.n89_cascade_\ : std_logic;
signal \tok.n83_adj_734_cascade_\ : std_logic;
signal \tok.n6279\ : std_logic;
signal \tok.table_rd_0\ : std_logic;
signal \tok.table_wr_data_14\ : std_logic;
signal \tok.table_wr_data_11\ : std_logic;
signal \tok.table_wr_data_12\ : std_logic;
signal \tok.n2696\ : std_logic;
signal \tok.n9_adj_651_cascade_\ : std_logic;
signal \tok.n13\ : std_logic;
signal \n15_cascade_\ : std_logic;
signal \tok.n6_adj_687_cascade_\ : std_logic;
signal \tok.n4_adj_641\ : std_logic;
signal \tok.n5\ : std_logic;
signal \tok.n796_cascade_\ : std_logic;
signal \tok.n12\ : std_logic;
signal \tok.n796\ : std_logic;
signal \tok.n2702\ : std_logic;
signal \tok.uart_stall\ : std_logic;
signal \tok.n6203\ : std_logic;
signal \tok.search_clk_N_137\ : std_logic;
signal \tok.n31_adj_637_cascade_\ : std_logic;
signal \tok.n6170\ : std_logic;
signal \tok.n30\ : std_logic;
signal \tok.n221_adj_753_cascade_\ : std_logic;
signal \tok.key_rd_3\ : std_logic;
signal \tok.key_rd_5\ : std_logic;
signal \tok.key_rd_8\ : std_logic;
signal \tok.n20_cascade_\ : std_logic;
signal \tok.n26_adj_645\ : std_logic;
signal \tok.key_rd_13\ : std_logic;
signal \tok.n14_adj_644\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \tok.n4782\ : std_logic;
signal \tok.n4783\ : std_logic;
signal \tok.n127\ : std_logic;
signal \tok.n4784\ : std_logic;
signal \tok.n6557\ : std_logic;
signal \tok.n4785\ : std_logic;
signal \tok.n320\ : std_logic;
signal \tok.n4786\ : std_logic;
signal \tok.n4787\ : std_logic;
signal \GNDG0\ : std_logic;
signal \tok.n4788\ : std_logic;
signal \tok.n4788_THRU_CRY_0_THRU_CO\ : std_logic;
signal \tok.n21_adj_660\ : std_logic;
signal \tok.n318\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \tok.n4789\ : std_logic;
signal \tok.n4790\ : std_logic;
signal \tok.n315\ : std_logic;
signal \tok.n4791\ : std_logic;
signal \tok.n4792\ : std_logic;
signal \tok.n313\ : std_logic;
signal \tok.n4793\ : std_logic;
signal \tok.n312\ : std_logic;
signal \tok.n295\ : std_logic;
signal \tok.n4794\ : std_logic;
signal \tok.n4795\ : std_logic;
signal \tok.n4796\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \tok.n293\ : std_logic;
signal \tok.n297\ : std_logic;
signal \tok.n310\ : std_logic;
signal \tok.n6452\ : std_logic;
signal \tok.n2579\ : std_logic;
signal \tok.n6392\ : std_logic;
signal \tok.n6421\ : std_logic;
signal \tok.n300\ : std_logic;
signal \tok.n6460\ : std_logic;
signal \tok.n161_adj_825\ : std_logic;
signal \tok.n197_adj_826\ : std_logic;
signal \tok.n18_adj_850\ : std_logic;
signal \tok.n17_adj_853\ : std_logic;
signal \tok.n31_cascade_\ : std_logic;
signal \tok.n299\ : std_logic;
signal \tok.n6446\ : std_logic;
signal \tok.n308\ : std_logic;
signal \tok.n294\ : std_logic;
signal \tok.n161_adj_667\ : std_logic;
signal \tok.n6371_cascade_\ : std_logic;
signal \tok.n248_adj_653\ : std_logic;
signal \tok.n200_adj_655_cascade_\ : std_logic;
signal \tok.n6_adj_658_cascade_\ : std_logic;
signal \tok.n6_adj_832_cascade_\ : std_logic;
signal \tok.n6383\ : std_logic;
signal \tok.n242_adj_654\ : std_logic;
signal \tok.S_13\ : std_logic;
signal \tok.S_8\ : std_logic;
signal \tok.n14_adj_844_cascade_\ : std_logic;
signal \tok.n20_adj_845\ : std_logic;
signal \tok.n26_adj_851\ : std_logic;
signal \tok.n6324_cascade_\ : std_logic;
signal \tok.n262_adj_858_cascade_\ : std_logic;
signal \tok.n268\ : std_logic;
signal \tok.n6315\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CONSTANT_ONE_NET_cascade_\ : std_logic;
signal \tok.n239\ : std_logic;
signal sender_2 : std_logic;
signal \tok.n6347\ : std_logic;
signal \tok.n197_adj_693\ : std_logic;
signal \tok.n248_adj_694_cascade_\ : std_logic;
signal \tok.n242_adj_695\ : std_logic;
signal \tok.n200_adj_696_cascade_\ : std_logic;
signal \tok.n6_adj_699_cascade_\ : std_logic;
signal \bfn_6_2_0_\ : std_logic;
signal \tok.n4812\ : std_logic;
signal \tok.n4813\ : std_logic;
signal \tok.n4814\ : std_logic;
signal \tok.n4815\ : std_logic;
signal \tok.n4816\ : std_logic;
signal \tok.n4817\ : std_logic;
signal \tok.n4818\ : std_logic;
signal \tok.n13_adj_760_cascade_\ : std_logic;
signal \n10_adj_905_cascade_\ : std_logic;
signal \tok.tc_5\ : std_logic;
signal \tok.ram.n6263_cascade_\ : std_logic;
signal \tok.n1530\ : std_logic;
signal \tok.n83_adj_759_cascade_\ : std_logic;
signal \tok.n6660\ : std_logic;
signal n10_adj_905 : std_logic;
signal \tok.n83_adj_764_cascade_\ : std_logic;
signal \tok.ram.n6277_cascade_\ : std_logic;
signal \n10_cascade_\ : std_logic;
signal \tok.tc_7\ : std_logic;
signal \tok.n1635\ : std_logic;
signal \tok.n6662\ : std_logic;
signal \tok.n13_adj_790\ : std_logic;
signal n10 : std_logic;
signal \tok.n5_adj_675\ : std_logic;
signal \tok.n6205_cascade_\ : std_logic;
signal \tok.n270\ : std_logic;
signal \tok.n270_cascade_\ : std_logic;
signal \tok.A_stk.tail_18\ : std_logic;
signal \A_stk_delta_1\ : std_logic;
signal \tok.A_stk.tail_2\ : std_logic;
signal \rd_15__N_300\ : std_logic;
signal \tok.n283_cascade_\ : std_logic;
signal \tok.n223_cascade_\ : std_logic;
signal \tok.n4_adj_752\ : std_logic;
signal \tok.n6586_cascade_\ : std_logic;
signal \tok.n226_adj_744\ : std_logic;
signal \tok.n254\ : std_logic;
signal \tok.n319\ : std_logic;
signal \tok.n6326\ : std_logic;
signal \tok.n387_cascade_\ : std_logic;
signal \tok.n254_adj_860_cascade_\ : std_logic;
signal \tok.n163\ : std_logic;
signal \tok.n256_adj_862\ : std_logic;
signal \tok.n5_adj_871\ : std_logic;
signal \tok.n6_adj_868_cascade_\ : std_logic;
signal \S_0\ : std_logic;
signal \tok.n28\ : std_logic;
signal \tok.key_rd_11\ : std_logic;
signal \tok.key_rd_14\ : std_logic;
signal \tok.n23_adj_638\ : std_logic;
signal \tok.key_rd_15\ : std_logic;
signal \tok.key_rd_9\ : std_logic;
signal \tok.n24\ : std_logic;
signal \tok.n26_adj_781\ : std_logic;
signal \tok.n28_adj_778_cascade_\ : std_logic;
signal \tok.n25_adj_788\ : std_logic;
signal \tok.S_15\ : std_logic;
signal \tok.n6634\ : std_logic;
signal \tok.n23_adj_848\ : std_logic;
signal \tok.n21_adj_849_cascade_\ : std_logic;
signal \tok.n24_adj_846\ : std_logic;
signal \tok.n30_adj_852\ : std_logic;
signal \tok.n323\ : std_logic;
signal \tok.n22_adj_847\ : std_logic;
signal \tok.n27_adj_782\ : std_logic;
signal \tok.n298\ : std_logic;
signal \tok.n161_adj_870\ : std_logic;
signal \tok.n6429_cascade_\ : std_logic;
signal \tok.n197_adj_872_cascade_\ : std_logic;
signal \tok.n248_adj_873\ : std_logic;
signal \tok.n296\ : std_logic;
signal \tok.n6400_cascade_\ : std_logic;
signal \tok.n161\ : std_logic;
signal \tok.n6406\ : std_logic;
signal \tok.n6415\ : std_logic;
signal \tok.n161_adj_882_cascade_\ : std_logic;
signal \tok.n208_adj_857\ : std_logic;
signal \tok.n6328\ : std_logic;
signal \tok.n250\ : std_logic;
signal \tok.n190_adj_774_cascade_\ : std_logic;
signal \tok.n6514\ : std_logic;
signal \tok.n833_cascade_\ : std_logic;
signal \tok.n6515\ : std_logic;
signal \tok.n6534_cascade_\ : std_logic;
signal \tok.n252_adj_783_cascade_\ : std_logic;
signal \tok.n255_adj_775\ : std_logic;
signal \tok.n190_adj_774\ : std_logic;
signal \tok.n258_adj_780\ : std_logic;
signal \tok.n177_adj_779\ : std_logic;
signal \tok.n6368\ : std_logic;
signal \tok.n197_adj_668\ : std_logic;
signal \tok.n248_adj_669_cascade_\ : std_logic;
signal \tok.n242_adj_670\ : std_logic;
signal \tok.n200_adj_671_cascade_\ : std_logic;
signal \tok.S_14\ : std_logic;
signal \tok.n6_adj_674_cascade_\ : std_logic;
signal \tok.table_rd_8\ : std_logic;
signal \tok.n7269\ : std_logic;
signal \tok.n203_adj_822_cascade_\ : std_logic;
signal \tok.n212_adj_824_cascade_\ : std_logic;
signal \tok.n6457_cascade_\ : std_logic;
signal \tok.n248_adj_827\ : std_logic;
signal \tok.n242_adj_828_cascade_\ : std_logic;
signal \tok.n200_adj_829\ : std_logic;
signal \tok.n231\ : std_logic;
signal \tok.n242_adj_885\ : std_logic;
signal \tok.n200_adj_886_cascade_\ : std_logic;
signal \tok.n6_adj_889_cascade_\ : std_logic;
signal \tok.n8_cascade_\ : std_logic;
signal \tok.S_11\ : std_logic;
signal \tok.n197_adj_883\ : std_logic;
signal \tok.n248_adj_884\ : std_logic;
signal \tok.n83_adj_756_cascade_\ : std_logic;
signal \tok.ram.n6260_cascade_\ : std_logic;
signal \tok.n6295\ : std_logic;
signal \tok.n1565_cascade_\ : std_logic;
signal \tok.n13_adj_757_cascade_\ : std_logic;
signal \n10_adj_906_cascade_\ : std_logic;
signal \tok.tc_4\ : std_logic;
signal n10_adj_906 : std_logic;
signal \tok.n324_cascade_\ : std_logic;
signal \tok.n225_adj_678\ : std_logic;
signal \tok.n225_adj_678_cascade_\ : std_logic;
signal \tok.n6351\ : std_logic;
signal \tok.n6632\ : std_logic;
signal \tok.n7456_cascade_\ : std_logic;
signal \tok.n176\ : std_logic;
signal \tok.n8_adj_686\ : std_logic;
signal \tok.n6622\ : std_logic;
signal \tok.n237_adj_724_cascade_\ : std_logic;
signal \tok.n4893\ : std_logic;
signal \tok.n286\ : std_logic;
signal \tok.n286_cascade_\ : std_logic;
signal \tok.n877\ : std_logic;
signal \tok.n394_cascade_\ : std_logic;
signal \tok.n6143\ : std_logic;
signal \tok.tc_3\ : std_logic;
signal \tok.tc_1\ : std_logic;
signal n92_adj_897 : std_logic;
signal \tok.tc_0\ : std_logic;
signal \stall_\ : std_logic;
signal \tok.tc_2\ : std_logic;
signal \tok.n6140\ : std_logic;
signal \tok.n6582\ : std_logic;
signal \tok.table_wr_data_5\ : std_logic;
signal \tok.n199_cascade_\ : std_logic;
signal \tok.n262\ : std_logic;
signal \tok.n4_adj_648_cascade_\ : std_logic;
signal \tok.n326\ : std_logic;
signal \tok.n234\ : std_logic;
signal \tok.table_rd_5\ : std_logic;
signal \tok.n4842_cascade_\ : std_logic;
signal \tok.n7451_cascade_\ : std_logic;
signal \tok.n6616\ : std_logic;
signal \tok.S_2\ : std_logic;
signal \tok.n164\ : std_logic;
signal \tok.n6597\ : std_logic;
signal \tok.n4_adj_711\ : std_logic;
signal \tok.n307\ : std_logic;
signal \tok.n6397\ : std_logic;
signal \tok.n242_cascade_\ : std_logic;
signal \tok.n197\ : std_logic;
signal \tok.n248\ : std_logic;
signal \tok.n6606_cascade_\ : std_logic;
signal \tok.n200\ : std_logic;
signal \tok.n6_cascade_\ : std_logic;
signal \tok.S_12\ : std_logic;
signal \tok.n200_adj_875\ : std_logic;
signal \tok.n6_adj_878_cascade_\ : std_logic;
signal \tok.S_10\ : std_logic;
signal \tok.n2600_cascade_\ : std_logic;
signal \tok.n6610_cascade_\ : std_logic;
signal \tok.n6344\ : std_logic;
signal \tok.n269_cascade_\ : std_logic;
signal \tok.n4_adj_786\ : std_logic;
signal \tok.n205_adj_789\ : std_logic;
signal \tok.n4_adj_635\ : std_logic;
signal \tok.n6341_cascade_\ : std_logic;
signal \tok.n170\ : std_logic;
signal \tok.n321\ : std_logic;
signal \tok.n4_adj_640\ : std_logic;
signal \tok.n4_adj_680\ : std_logic;
signal \tok.n239_adj_679\ : std_logic;
signal \tok.n238_adj_681_cascade_\ : std_logic;
signal \tok.n900\ : std_logic;
signal \tok.n317_adj_659\ : std_logic;
signal \tok.n2663\ : std_logic;
signal \tok.uart.sender_5\ : std_logic;
signal \tok.uart.sender_4\ : std_logic;
signal \tok.uart.sender_3\ : std_logic;
signal \tok.n2602\ : std_logic;
signal \tok.n6450\ : std_logic;
signal \tok.n215_adj_830_cascade_\ : std_logic;
signal \tok.n6605_cascade_\ : std_logic;
signal \tok.n6604\ : std_logic;
signal \tok.n6456\ : std_logic;
signal \tok.n179_adj_831\ : std_logic;
signal \tok.n214\ : std_logic;
signal \tok.n6462_cascade_\ : std_logic;
signal \tok.n786\ : std_logic;
signal \tok.n206_adj_823\ : std_logic;
signal \tok.n314\ : std_logic;
signal \tok.n6425\ : std_logic;
signal \tok.n6346\ : std_logic;
signal \tok.n215_adj_876\ : std_logic;
signal \tok.n179_adj_877\ : std_logic;
signal \tok.n6553_cascade_\ : std_logic;
signal \tok.n6552\ : std_logic;
signal \tok.n179_adj_698\ : std_logic;
signal \tok.n6537\ : std_logic;
signal \tok.n6541_cascade_\ : std_logic;
signal \tok.n6540\ : std_logic;
signal \tok.n6367\ : std_logic;
signal \tok.n179_adj_673\ : std_logic;
signal tc_plus_1_0 : std_logic;
signal \tok.C_stk.n6230_cascade_\ : std_logic;
signal tc_0 : std_logic;
signal c_stk_r_0 : std_logic;
signal \tok.C_stk.tail_0\ : std_logic;
signal \tok.tc_plus_1_4\ : std_logic;
signal \tok.C_stk.n6239_cascade_\ : std_logic;
signal tc_4 : std_logic;
signal \tok.c_stk_r_4\ : std_logic;
signal \tok.C_stk.tail_4\ : std_logic;
signal \tok.tail_12\ : std_logic;
signal \tok.C_stk.tail_20\ : std_logic;
signal \tok.tail_28\ : std_logic;
signal \tok.C_stk.tail_36\ : std_logic;
signal \tok.n83_adj_723_cascade_\ : std_logic;
signal n10_adj_908 : std_logic;
signal \tok.n4_adj_726_cascade_\ : std_logic;
signal \tok.ram.n6257_cascade_\ : std_logic;
signal \tok.n6664\ : std_logic;
signal \tok.n1600_cascade_\ : std_logic;
signal \tok.n13_adj_742\ : std_logic;
signal \tok.n6301_cascade_\ : std_logic;
signal \tok.n80_adj_751_cascade_\ : std_logic;
signal \tok.n83_adj_746_cascade_\ : std_logic;
signal \tok.n6297\ : std_logic;
signal \tok.n89_adj_754\ : std_logic;
signal n92_adj_898 : std_logic;
signal \tok.table_rd_3\ : std_logic;
signal \tok.n14_adj_683_cascade_\ : std_logic;
signal \tok.n9_adj_651\ : std_logic;
signal \tok.n15_adj_807_cascade_\ : std_logic;
signal \tok.n903\ : std_logic;
signal \tok.n14_adj_683\ : std_logic;
signal \tok.n6621\ : std_logic;
signal \tok.n241_adj_747\ : std_logic;
signal \tok.n6593\ : std_logic;
signal \tok.n236\ : std_logic;
signal \tok.n4925\ : std_logic;
signal \tok.n288\ : std_logic;
signal \tok.n2613\ : std_logic;
signal \tok.n6578_cascade_\ : std_logic;
signal \tok.n6581\ : std_logic;
signal \tok.n4_adj_739\ : std_logic;
signal \tok.n2611\ : std_logic;
signal \tok.n6580\ : std_logic;
signal \tok.n4_adj_684\ : std_logic;
signal \tok.n6620_cascade_\ : std_logic;
signal \tok.n311_adj_721\ : std_logic;
signal \tok.n167_cascade_\ : std_logic;
signal \tok.n6567\ : std_logic;
signal \tok.table_rd_2\ : std_logic;
signal \tok.n209_cascade_\ : std_logic;
signal \tok.n6625_cascade_\ : std_logic;
signal \tok.n6624\ : std_logic;
signal \tok.n168_adj_700_cascade_\ : std_logic;
signal \tok.n6569\ : std_logic;
signal \tok.n2548\ : std_logic;
signal \tok.n6396\ : std_logic;
signal \tok.n179_cascade_\ : std_logic;
signal \tok.n6546\ : std_logic;
signal \tok.table_rd_7\ : std_logic;
signal \tok.table_rd_4\ : std_logic;
signal \tok.n258_adj_814\ : std_logic;
signal \tok.n252_adj_815_cascade_\ : std_logic;
signal \tok.n232\ : std_logic;
signal \tok.n255_adj_808\ : std_logic;
signal \tok.n210_adj_816\ : std_logic;
signal \tok.n872_cascade_\ : std_logic;
signal \tok.n174_adj_817_cascade_\ : std_logic;
signal \tok.n4_adj_818\ : std_logic;
signal \tok.n205_adj_820\ : std_logic;
signal \tok.n200_adj_840\ : std_logic;
signal \tok.n6_adj_843_cascade_\ : std_logic;
signal \tok.S_9\ : std_logic;
signal \tok.n6440_cascade_\ : std_logic;
signal \tok.n6612_cascade_\ : std_logic;
signal \tok.n6365\ : std_logic;
signal \tok.n215_adj_672\ : std_logic;
signal \tok.n252\ : std_logic;
signal \tok.n4_adj_769_cascade_\ : std_logic;
signal \tok.n205_adj_770\ : std_logic;
signal \tok.n235\ : std_logic;
signal \tok.n190_cascade_\ : std_logic;
signal \tok.n190\ : std_logic;
signal \tok.n255_cascade_\ : std_logic;
signal \tok.n258\ : std_logic;
signal \tok.n6508_cascade_\ : std_logic;
signal \tok.n6532\ : std_logic;
signal \tok.n207_adj_771_cascade_\ : std_logic;
signal \tok.n6583\ : std_logic;
signal \tok.S_5\ : std_logic;
signal \tok.n213\ : std_logic;
signal \tok.n207_adj_776_cascade_\ : std_logic;
signal \tok.n6529_cascade_\ : std_logic;
signal \tok.n210_adj_784\ : std_logic;
signal \tok.n174_adj_785\ : std_logic;
signal \tok.n229_adj_861\ : std_logic;
signal \tok.n6320\ : std_logic;
signal \tok.n49\ : std_logic;
signal \tok.n6380_cascade_\ : std_logic;
signal \tok.n215_adj_656_cascade_\ : std_logic;
signal \tok.n2665\ : std_logic;
signal \tok.n4_adj_719\ : std_logic;
signal \tok.n4_adj_719_cascade_\ : std_logic;
signal \tok.n10_adj_809\ : std_logic;
signal \tok.n6411\ : std_logic;
signal \tok.n6404_cascade_\ : std_logic;
signal \tok.n179_adj_888\ : std_logic;
signal \tok.n6550_cascade_\ : std_logic;
signal \tok.n6549\ : std_logic;
signal \tok.n6419\ : std_logic;
signal \tok.n215_adj_697\ : std_logic;
signal \tok.n6337_cascade_\ : std_logic;
signal \tok.n6538\ : std_logic;
signal \tok.tc_plus_1_5\ : std_logic;
signal \tok.C_stk.n6236_cascade_\ : std_logic;
signal tc_5 : std_logic;
signal \tok.c_stk_r_5\ : std_logic;
signal \tok.C_stk.tail_5\ : std_logic;
signal \tok.tail_13\ : std_logic;
signal \tok.C_stk.tail_21\ : std_logic;
signal \tok.tail_29\ : std_logic;
signal \tok.C_stk.tail_37\ : std_logic;
signal \tok.tc_plus_1_2\ : std_logic;
signal \tok.C_stk.n6245_cascade_\ : std_logic;
signal tc_2 : std_logic;
signal \tok.c_stk_r_2\ : std_logic;
signal \tok.C_stk.tail_2\ : std_logic;
signal \tok.tail_10\ : std_logic;
signal \tok.C_stk.tail_18\ : std_logic;
signal \tok.tail_26\ : std_logic;
signal \tok.C_stk.tail_34\ : std_logic;
signal \tok.tc_plus_1_3\ : std_logic;
signal \tok.C_stk.n6242_cascade_\ : std_logic;
signal tc_3 : std_logic;
signal \tok.c_stk_r_3\ : std_logic;
signal \tok.C_stk.tail_3\ : std_logic;
signal \tok.C_stk.tail_11\ : std_logic;
signal \tok.C_stk.tail_19\ : std_logic;
signal \tok.C_stk.tail_27\ : std_logic;
signal \tok.C_stk.tail_35\ : std_logic;
signal \tok.n4_adj_726\ : std_logic;
signal \tok.tc__7__N_133\ : std_logic;
signal \tok.n2573\ : std_logic;
signal \tok.n6291_cascade_\ : std_logic;
signal \tok.n80_adj_735_cascade_\ : std_logic;
signal \tok.n83_adj_725_cascade_\ : std_logic;
signal \tok.n6287\ : std_logic;
signal \tok.n89_adj_736\ : std_logic;
signal n92 : std_logic;
signal \tok.n4926\ : std_logic;
signal \tok.n2692_cascade_\ : std_logic;
signal \tok.n217\ : std_logic;
signal \tok.n7154\ : std_logic;
signal \tok.n6_adj_701\ : std_logic;
signal \tok.n2700\ : std_logic;
signal \tok.n236_adj_737\ : std_logic;
signal \tok.n239_adj_738\ : std_logic;
signal \tok.n17\ : std_logic;
signal \tok.n5_adj_821\ : std_logic;
signal \tok.n2679\ : std_logic;
signal \tok.n17_cascade_\ : std_logic;
signal \tok.n864\ : std_logic;
signal \tok.n186\ : std_logic;
signal \tok.n6562_cascade_\ : std_logic;
signal \tok.n338\ : std_logic;
signal \tok.n162\ : std_logic;
signal \tok.n179_adj_730\ : std_logic;
signal \tok.n197_adj_729_cascade_\ : std_logic;
signal \tok.n7458\ : std_logic;
signal \tok.n2544\ : std_logic;
signal \tok.table_rd_1\ : std_logic;
signal \tok.n7475_cascade_\ : std_logic;
signal \tok.n237\ : std_logic;
signal \tok.n180\ : std_logic;
signal \tok.n6628\ : std_logic;
signal \tok.S_3\ : std_logic;
signal \tok.n241\ : std_logic;
signal \tok.n6637\ : std_logic;
signal \tok.n284_cascade_\ : std_logic;
signal \tok.n244_cascade_\ : std_logic;
signal \tok.n4_adj_720_cascade_\ : std_logic;
signal \tok.n145\ : std_logic;
signal \tok.n251\ : std_logic;
signal \tok.n2557\ : std_logic;
signal \tok.n4_adj_714_cascade_\ : std_logic;
signal \tok.n218\ : std_logic;
signal \tok.n39\ : std_logic;
signal \tok.n6269_cascade_\ : std_logic;
signal \tok.n6466\ : std_logic;
signal \tok.n6467\ : std_logic;
signal \tok.n6486\ : std_logic;
signal \tok.n833\ : std_logic;
signal \tok.n6490\ : std_logic;
signal \tok.n6491\ : std_logic;
signal \S_1\ : std_logic;
signal \tok.n208\ : std_logic;
signal \tok.n6589\ : std_logic;
signal \tok.n239_adj_727\ : std_logic;
signal \tok.n6_adj_728_cascade_\ : std_logic;
signal \tok.n200_adj_732_cascade_\ : std_logic;
signal \tok.n203_adj_731\ : std_logic;
signal \tok.n6_adj_733\ : std_logic;
signal \tok.n206_adj_794\ : std_logic;
signal \tok.n207_adj_811_cascade_\ : std_logic;
signal \tok.n6481\ : std_logic;
signal \tok.n6484\ : std_logic;
signal \tok.n213_adj_810\ : std_logic;
signal \tok.S_4\ : std_logic;
signal \tok.n207_cascade_\ : std_logic;
signal \tok.n210\ : std_logic;
signal \tok.n6572_cascade_\ : std_logic;
signal \tok.n174_adj_768\ : std_logic;
signal \tok.n31\ : std_logic;
signal \tok.n26_adj_763\ : std_logic;
signal \tok.n26_adj_763_cascade_\ : std_logic;
signal \tok.n4_adj_636\ : std_logic;
signal \tok.n213_adj_795\ : std_logic;
signal \tok.n207_adj_796_cascade_\ : std_logic;
signal \tok.n872\ : std_logic;
signal \tok.n6505_cascade_\ : std_logic;
signal \tok.n42\ : std_logic;
signal \tok.n6360\ : std_logic;
signal \tok.table_rd_6\ : std_logic;
signal \tok.n210_adj_802\ : std_logic;
signal \tok.n316\ : std_logic;
signal \tok.n6409_cascade_\ : std_logic;
signal \tok.n46\ : std_logic;
signal \tok.n215_adj_887\ : std_logic;
signal \tok.n6442\ : std_logic;
signal \tok.n6433_cascade_\ : std_logic;
signal \tok.n215_adj_841\ : std_logic;
signal \tok.n179_adj_842\ : std_logic;
signal \tok.n6602_cascade_\ : std_logic;
signal \tok.n6601\ : std_logic;
signal \tok.n6375\ : std_logic;
signal \tok.n847\ : std_logic;
signal \tok.n6544\ : std_logic;
signal \tok.n179_adj_657_cascade_\ : std_logic;
signal \tok.n6543\ : std_logic;
signal \tok.n464\ : std_logic;
signal \tok.n8\ : std_logic;
signal \tok.n6382\ : std_logic;
signal tail_40 : std_logic;
signal tail_8 : std_logic;
signal \tok.C_stk.tail_32\ : std_logic;
signal \tok.C_stk.tail_16\ : std_logic;
signal tail_24 : std_logic;
signal \tok.C_stk.tail_43\ : std_logic;
signal \tok.tail_45\ : std_logic;
signal \tok.tail_44\ : std_logic;
signal \tok.tail_42\ : std_logic;
signal tail_51 : std_logic;
signal tail_59 : std_logic;
signal tail_48_adj_900 : std_logic;
signal tail_56 : std_logic;
signal \C_stk_delta_1_cascade_\ : std_logic;
signal tail_57 : std_logic;
signal \tok.tail_52\ : std_logic;
signal \tok.tail_60\ : std_logic;
signal \tok.tail_62\ : std_logic;
signal \tok.n37\ : std_logic;
signal \tok.n2559\ : std_logic;
signal \tok.tail_53\ : std_logic;
signal \rd_7__N_373_cascade_\ : std_logic;
signal \tok.tail_61\ : std_logic;
signal tc_plus_1_1 : std_logic;
signal \tok.C_stk.n6248_cascade_\ : std_logic;
signal tc_1 : std_logic;
signal c_stk_r_1 : std_logic;
signal \tok.C_stk.tail_1\ : std_logic;
signal tail_9 : std_logic;
signal \tok.C_stk.tail_17\ : std_logic;
signal tail_25 : std_logic;
signal tail_49_adj_899 : std_logic;
signal \tok.C_stk.tail_33\ : std_logic;
signal tail_41 : std_logic;
signal \tok.n156\ : std_logic;
signal \tok.n211_adj_741_cascade_\ : std_logic;
signal \tok.n277_cascade_\ : std_logic;
signal \tok.n265\ : std_logic;
signal \tok.n6_adj_748\ : std_logic;
signal \tok.n6331\ : std_logic;
signal \tok.n238_adj_855_cascade_\ : std_logic;
signal \tok.n4_adj_859\ : std_logic;
signal \tok.n6_adj_676\ : std_logic;
signal \tok.n298_adj_856\ : std_logic;
signal \tok.n53_cascade_\ : std_logic;
signal \tok.n992\ : std_logic;
signal \tok.n2_cascade_\ : std_logic;
signal \tok.n23\ : std_logic;
signal \tok.n174_cascade_\ : std_logic;
signal \tok.stall\ : std_logic;
signal \tok.n6189\ : std_logic;
signal \tok.n6_adj_722\ : std_logic;
signal \tok.n127_adj_772\ : std_logic;
signal \tok.n10_adj_773_cascade_\ : std_logic;
signal \tok.n6146_cascade_\ : std_logic;
signal \tok.n86\ : std_logic;
signal \tok.n5_adj_715\ : std_logic;
signal \tok.n369_cascade_\ : std_logic;
signal \tok.n278\ : std_logic;
signal \tok.n233_adj_716_cascade_\ : std_logic;
signal \tok.n229\ : std_logic;
signal \tok.n6156\ : std_logic;
signal \tok.n7\ : std_logic;
signal \tok.n4_adj_648\ : std_logic;
signal \tok.n2635\ : std_logic;
signal \tok.n6653_cascade_\ : std_logic;
signal \tok.n6646_cascade_\ : std_logic;
signal \tok.n6167\ : std_logic;
signal \tok.n6645\ : std_logic;
signal \tok.n247\ : std_logic;
signal \tok.n6639\ : std_logic;
signal \tok.n280\ : std_logic;
signal \tok.n6638_cascade_\ : std_logic;
signal \tok.n6636\ : std_logic;
signal \tok.n260_adj_717\ : std_logic;
signal \tok.S_6\ : std_logic;
signal \tok.n815\ : std_logic;
signal \tok.n6510\ : std_logic;
signal \tok.n177_adj_799_cascade_\ : std_logic;
signal \tok.n252_adj_801_cascade_\ : std_logic;
signal \tok.n867\ : std_logic;
signal \tok.n233\ : std_logic;
signal \tok.n5_adj_745\ : std_logic;
signal \tok.n255_adj_793_cascade_\ : std_logic;
signal \tok.n258_adj_800\ : std_logic;
signal \tok.n6183\ : std_logic;
signal \tok.n6162_cascade_\ : std_logic;
signal \tok.n865_cascade_\ : std_logic;
signal \tok.n222_cascade_\ : std_logic;
signal \tok.n245\ : std_logic;
signal \tok.n6501\ : std_logic;
signal \tok.n186_adj_798_cascade_\ : std_logic;
signal \tok.n6496\ : std_logic;
signal \tok.n194\ : std_logic;
signal \tok.n338_adj_805_cascade_\ : std_logic;
signal \tok.n6608\ : std_logic;
signal \tok.n219\ : std_logic;
signal \tok.n190_adj_792\ : std_logic;
signal \tok.n4_adj_804\ : std_logic;
signal \tok.n174_adj_803\ : std_logic;
signal \tok.n205_adj_806\ : std_logic;
signal \tok.n177_adj_813\ : std_logic;
signal \tok.n2598_cascade_\ : std_logic;
signal \tok.n45\ : std_logic;
signal \tok.n6390\ : std_logic;
signal \tok.n821\ : std_logic;
signal \tok.n215_cascade_\ : std_logic;
signal \tok.n6547\ : std_logic;
signal \tok.n4_adj_712\ : std_logic;
signal \tok.n238\ : std_logic;
signal \tok.n6650_cascade_\ : std_logic;
signal \tok.n48\ : std_logic;
signal \tok.n211_cascade_\ : std_logic;
signal \tok.n6644\ : std_logic;
signal \tok.n260_cascade_\ : std_logic;
signal \tok.n6641\ : std_logic;
signal \tok.n266_cascade_\ : std_logic;
signal \tok.n5_adj_713\ : std_logic;
signal \tok.n256\ : std_logic;
signal \tok.n4_adj_718_cascade_\ : std_logic;
signal \tok.n221\ : std_logic;
signal \tok.A_low_1\ : std_logic;
signal \tok.n2637\ : std_logic;
signal \tok.A_low_4\ : std_logic;
signal \tok.uart.sender_6\ : std_logic;
signal \tok.uart.sender_7\ : std_logic;
signal \tok.uart.sender_8\ : std_logic;
signal \tok.uart.n950\ : std_logic;
signal \tok.n274\ : std_logic;
signal \tok.n185\ : std_logic;
signal \tok.n7410\ : std_logic;
signal reset_c : std_logic;
signal \tok.tail_50\ : std_logic;
signal \tok.tail_58\ : std_logic;
signal \tok.tc_plus_1_6\ : std_logic;
signal \tok.C_stk.n6233_cascade_\ : std_logic;
signal tc_6 : std_logic;
signal \tok.c_stk_r_6\ : std_logic;
signal \tok.C_stk.tail_6\ : std_logic;
signal \tok.tail_14\ : std_logic;
signal \tok.C_stk.tail_22\ : std_logic;
signal \tok.tail_30\ : std_logic;
signal \tok.tail_54\ : std_logic;
signal \tok.C_stk.tail_38\ : std_logic;
signal \tok.tail_46\ : std_logic;
signal \tok.C_stk.n449\ : std_logic;
signal \tok.n273\ : std_logic;
signal tc_7 : std_logic;
signal \tok.C_stk.n6227_cascade_\ : std_logic;
signal \tok.n15\ : std_logic;
signal \tok.c_stk_r_7\ : std_logic;
signal \tok.C_stk.tail_7\ : std_logic;
signal \tok.tail_15\ : std_logic;
signal \tok.C_stk.tail_23\ : std_logic;
signal \tok.tail_31\ : std_logic;
signal \tok.C_stk.tail_39\ : std_logic;
signal \tok.tail_47\ : std_logic;
signal \rd_7__N_373\ : std_logic;
signal \tok.tail_55\ : std_logic;
signal \C_stk_delta_1\ : std_logic;
signal \tok.tail_63\ : std_logic;
signal n15 : std_logic;
signal \tok.tc_plus_1_7\ : std_logic;
signal \tok.S_7\ : std_logic;
signal \tok.table_wr_data_7\ : std_logic;
signal uart_rx_data_4 : std_logic;
signal uart_rx_data_2 : std_logic;
signal uart_rx_data_1 : std_logic;
signal capture_2 : std_logic;
signal \tok.A_stk_delta_1__N_4\ : std_logic;
signal \tok.A_stk_delta_1__N_4_cascade_\ : std_logic;
signal \tok.n1\ : std_logic;
signal \tok.n4_adj_702_cascade_\ : std_logic;
signal \tok.n52\ : std_logic;
signal \tok.n51_cascade_\ : std_logic;
signal \tok.n50\ : std_logic;
signal \tok.n8_adj_854\ : std_logic;
signal \tok.n174\ : std_logic;
signal \tok.n4_adj_702\ : std_logic;
signal \tok.reset_N_2\ : std_logic;
signal \tok.n256_adj_749\ : std_logic;
signal \tok.n367\ : std_logic;
signal \tok.n215_adj_750\ : std_logic;
signal \tok.depth_2\ : std_logic;
signal \tok.depth_1\ : std_logic;
signal \tok.n741\ : std_logic;
signal \tok.n806\ : std_logic;
signal \tok.depth_0\ : std_logic;
signal \tok.n6213\ : std_logic;
signal \tok.n806_cascade_\ : std_logic;
signal \tok.depth_3\ : std_logic;
signal \tok.n748\ : std_logic;
signal \tok.n47\ : std_logic;
signal \tok.n6615\ : std_logic;
signal \tok.n158_cascade_\ : std_logic;
signal \tok.n6627\ : std_logic;
signal \tok.uart_stall_N_46\ : std_logic;
signal \tok.n9\ : std_logic;
signal \tok.n10\ : std_logic;
signal \tok.n10_cascade_\ : std_logic;
signal \tok.write_flag\ : std_logic;
signal \tok.n14\ : std_logic;
signal \tok.uart.n10_cascade_\ : std_logic;
signal \n23_cascade_\ : std_logic;
signal \tok.n168_adj_710_cascade_\ : std_logic;
signal \tok.A_low_6\ : std_logic;
signal \tok.n6502\ : std_logic;
signal uart_rx_data_6 : std_logic;
signal \tok.n43\ : std_logic;
signal \tok.n311\ : std_logic;
signal \tok.n190_adj_797\ : std_logic;
signal \tok.n44\ : std_logic;
signal \tok.T_2\ : std_logic;
signal \tok.T_0\ : std_logic;
signal \tok.n168_adj_690\ : std_logic;
signal \tok.n6525\ : std_logic;
signal \tok.n6526_cascade_\ : std_logic;
signal \tok.n186_adj_777_cascade_\ : std_logic;
signal \tok.n338_adj_787\ : std_logic;
signal \tok.A_low_0\ : std_logic;
signal \tok.A_low_5\ : std_logic;
signal \tok.n866_cascade_\ : std_logic;
signal \tok.n6520\ : std_logic;
signal \tok.T_5\ : std_logic;
signal \tok.n317\ : std_logic;
signal \tok.n317_cascade_\ : std_logic;
signal \tok.A_low_3\ : std_logic;
signal \tok.n168\ : std_logic;
signal \tok.n5_adj_682\ : std_logic;
signal \tok.T_4\ : std_logic;
signal \tok.n6478_cascade_\ : std_logic;
signal \tok.T_6\ : std_logic;
signal \tok.n186_adj_812_cascade_\ : std_logic;
signal \tok.T_3\ : std_logic;
signal \tok.n338_adj_819\ : std_logic;
signal \tok.T_7\ : std_logic;
signal \tok.A_low_2\ : std_logic;
signal \tok.n289\ : std_logic;
signal \tok.T_1\ : std_logic;
signal \tok.n222\ : std_logic;
signal \tok.n838\ : std_logic;
signal \tok.n863_cascade_\ : std_logic;
signal \tok.n6472\ : std_logic;
signal \tok.n9_adj_677\ : std_logic;
signal \tok.n205\ : std_logic;
signal \tok.n6477\ : std_logic;
signal capture_8 : std_logic;
signal uart_rx_data_7 : std_logic;
signal txtick : std_logic;
signal n23 : std_logic;
signal \A_low_7\ : std_logic;
signal sender_9 : std_logic;
signal capture_3 : std_logic;
signal capture_5 : std_logic;
signal \tok.n891\ : std_logic;
signal \tok.uart_rx_valid\ : std_logic;
signal \tok.uart.n922\ : std_logic;
signal capture_7 : std_logic;
signal capture_0 : std_logic;
signal capture_4 : std_logic;
signal \rx_data_7__N_510_cascade_\ : std_logic;
signal uart_rx_data_3 : std_logic;
signal capture_9 : std_logic;
signal capture_6 : std_logic;
signal uart_rx_data_5 : std_logic;
signal capture_1 : std_logic;
signal \rx_data_7__N_510\ : std_logic;
signal uart_rx_data_0 : std_logic;
signal \tok.uart_tx_busy\ : std_logic;
signal \tok.uart.sentbits_3\ : std_logic;
signal \tok.uart.sentbits_2\ : std_logic;
signal \tok.uart.sentbits_1\ : std_logic;
signal \tok.uart.sentbits_0\ : std_logic;
signal \tok.uart.n994\ : std_logic;
signal \tok.uart.n1013\ : std_logic;
signal rx_c : std_logic;
signal \tok.uart.n4977\ : std_logic;
signal \tok.uart.n4977_cascade_\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \tok.uart.n4819\ : std_logic;
signal \tok.uart.n4820\ : std_logic;
signal \tok.uart.bytephase_3\ : std_logic;
signal \tok.uart.n4821\ : std_logic;
signal \tok.uart.bytephase_4\ : std_logic;
signal \tok.uart.n4822\ : std_logic;
signal \tok.uart.n4823\ : std_logic;
signal \tok.uart.bytephase_5\ : std_logic;
signal n4928 : std_logic;
signal \tok.uart.n6_cascade_\ : std_logic;
signal \n746_cascade_\ : std_logic;
signal \bytephase_5__N_509\ : std_logic;
signal n974 : std_logic;
signal \tok.uart.n6211\ : std_logic;
signal \tok.uart.n2356\ : std_logic;
signal \tok.uart.n809\ : std_logic;
signal \tok.uart.n2356_cascade_\ : std_logic;
signal n746 : std_logic;
signal \tok.uart.bytephase_2\ : std_logic;
signal \tok.uart.bytephase_0\ : std_logic;
signal \tok.uart.bytephase_1\ : std_logic;
signal \tok.uart.n2357\ : std_logic;
signal \tok.uart.rxclkcounter_0\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \tok.uart.rxclkcounter_1\ : std_logic;
signal \tok.uart.n4824\ : std_logic;
signal \tok.uart.rxclkcounter_2\ : std_logic;
signal \tok.uart.n4825\ : std_logic;
signal \tok.uart.rxclkcounter_3\ : std_logic;
signal \tok.uart.n4826\ : std_logic;
signal \tok.uart.rxclkcounter_4\ : std_logic;
signal \tok.uart.n4827\ : std_logic;
signal \tok.uart.rxclkcounter_5\ : std_logic;
signal \tok.uart.n4828\ : std_logic;
signal \tok.uart.n4829\ : std_logic;
signal \tok.uart.rxclkcounter_6\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk : std_logic;
signal \tok.uart.rxclkcounter_6__N_476\ : std_logic;

signal rx_wire : std_logic;
signal reset_wire : std_logic;
signal tx_wire : std_logic;
signal \tok.vals.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.vals.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.vals.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.vals.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \tok.vals.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.keys.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.keys.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.keys.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.keys.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \tok.keys.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.ram.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.ram.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.ram.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.ram.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \tok.ram.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    rx_wire <= rx;
    reset_wire <= reset;
    tx <= tx_wire;
    \tok.table_rd_15\ <= \tok.vals.mem1_physical_RDATA_wire\(15);
    \tok.table_rd_14\ <= \tok.vals.mem1_physical_RDATA_wire\(14);
    \tok.table_rd_13\ <= \tok.vals.mem1_physical_RDATA_wire\(13);
    \tok.table_rd_12\ <= \tok.vals.mem1_physical_RDATA_wire\(12);
    \tok.table_rd_11\ <= \tok.vals.mem1_physical_RDATA_wire\(11);
    \tok.table_rd_10\ <= \tok.vals.mem1_physical_RDATA_wire\(10);
    \tok.table_rd_9\ <= \tok.vals.mem1_physical_RDATA_wire\(9);
    \tok.table_rd_8\ <= \tok.vals.mem1_physical_RDATA_wire\(8);
    \tok.table_rd_7\ <= \tok.vals.mem1_physical_RDATA_wire\(7);
    \tok.table_rd_6\ <= \tok.vals.mem1_physical_RDATA_wire\(6);
    \tok.table_rd_5\ <= \tok.vals.mem1_physical_RDATA_wire\(5);
    \tok.table_rd_4\ <= \tok.vals.mem1_physical_RDATA_wire\(4);
    \tok.table_rd_3\ <= \tok.vals.mem1_physical_RDATA_wire\(3);
    \tok.table_rd_2\ <= \tok.vals.mem1_physical_RDATA_wire\(2);
    \tok.table_rd_1\ <= \tok.vals.mem1_physical_RDATA_wire\(1);
    \tok.table_rd_0\ <= \tok.vals.mem1_physical_RDATA_wire\(0);
    \tok.vals.mem1_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__14469\&\N__15849\&\N__15402\&\N__14700\&\N__15539\&\N__15633\&\N__15465\&\N__14532\;
    \tok.vals.mem1_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__14466\&\N__15852\&\N__15399\&\N__14697\&\N__15536\&\N__15636\&\N__15468\&\N__14529\;
    \tok.vals.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \tok.vals.mem1_physical_WDATA_wire\ <= \N__14563\&\N__16507\&\N__14590\&\N__16477\&\N__16492\&\N__14578\&\N__15319\&\N__13384\&\N__28243\&\N__16309\&\N__19966\&\N__16294\&\N__16339\&\N__16282\&\N__16324\&\N__14389\;
    \tok.key_rd_15\ <= \tok.keys.mem0_physical_RDATA_wire\(15);
    \tok.key_rd_14\ <= \tok.keys.mem0_physical_RDATA_wire\(14);
    \tok.key_rd_13\ <= \tok.keys.mem0_physical_RDATA_wire\(13);
    \tok.key_rd_12\ <= \tok.keys.mem0_physical_RDATA_wire\(12);
    \tok.key_rd_11\ <= \tok.keys.mem0_physical_RDATA_wire\(11);
    \tok.key_rd_10\ <= \tok.keys.mem0_physical_RDATA_wire\(10);
    \tok.key_rd_9\ <= \tok.keys.mem0_physical_RDATA_wire\(9);
    \tok.key_rd_8\ <= \tok.keys.mem0_physical_RDATA_wire\(8);
    \tok.key_rd_7\ <= \tok.keys.mem0_physical_RDATA_wire\(7);
    \tok.key_rd_6\ <= \tok.keys.mem0_physical_RDATA_wire\(6);
    \tok.key_rd_5\ <= \tok.keys.mem0_physical_RDATA_wire\(5);
    \tok.key_rd_4\ <= \tok.keys.mem0_physical_RDATA_wire\(4);
    \tok.key_rd_3\ <= \tok.keys.mem0_physical_RDATA_wire\(3);
    \tok.key_rd_2\ <= \tok.keys.mem0_physical_RDATA_wire\(2);
    \tok.key_rd_1\ <= \tok.keys.mem0_physical_RDATA_wire\(1);
    \tok.key_rd_0\ <= \tok.keys.mem0_physical_RDATA_wire\(0);
    \tok.keys.mem0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__14479\&\N__15861\&\N__15412\&\N__14710\&\N__15550\&\N__15645\&\N__15477\&\N__14542\;
    \tok.keys.mem0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__14478\&\N__15862\&\N__15411\&\N__14709\&\N__15549\&\N__15646\&\N__15478\&\N__14541\;
    \tok.keys.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \tok.keys.mem0_physical_WDATA_wire\ <= \N__24196\&\N__32379\&\N__32233\&\N__27043\&\N__24001\&\N__29629\&\N__26793\&\N__22255\&\N__37442\&\N__30038\&\N__30320\&\N__27388\&\N__36532\&\N__33642\&\N__27514\&\N__30511\;
    \tok.T_7\ <= \tok.ram.mem2_physical_RDATA_wire\(14);
    \tok.T_6\ <= \tok.ram.mem2_physical_RDATA_wire\(12);
    \tok.T_5\ <= \tok.ram.mem2_physical_RDATA_wire\(10);
    \tok.T_4\ <= \tok.ram.mem2_physical_RDATA_wire\(8);
    \tok.T_3\ <= \tok.ram.mem2_physical_RDATA_wire\(6);
    \tok.T_2\ <= \tok.ram.mem2_physical_RDATA_wire\(4);
    \tok.T_1\ <= \tok.ram.mem2_physical_RDATA_wire\(2);
    \tok.T_0\ <= \tok.ram.mem2_physical_RDATA_wire\(0);
    \tok.ram.mem2_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__17680\&\N__16438\&\N__17623\&\N__19555\&\N__19831\&\N__19669\&\N__19813\&\N__19771\;
    \tok.ram.mem2_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__37466\&\N__30065\&\N__30342\&\N__27394\&\N__36556\&\N__33645\&\N__27561\&\N__30527\;
    \tok.ram.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \tok.ram.mem2_physical_WDATA_wire\ <= '0'&\N__37468\&'0'&\N__30085\&'0'&\N__30318\&'0'&\N__27391\&'0'&\N__36553\&'0'&\N__33643\&'0'&\N__27551\&'0'&\N__30507\;

    \tok.vals.mem1_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \tok.vals.mem1_physical_RDATA_wire\,
            RADDR => \tok.vals.mem1_physical_RADDR_wire\,
            WADDR => \tok.vals.mem1_physical_WADDR_wire\,
            MASK => \tok.vals.mem1_physical_MASK_wire\,
            WDATA => \tok.vals.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__38468\,
            RE => \N__17518\,
            WCLKE => 'H',
            WCLK => \N__38467\,
            WE => \N__14631\
        );

    \tok.keys.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \tok.keys.mem0_physical_RDATA_wire\,
            RADDR => \tok.keys.mem0_physical_RADDR_wire\,
            WADDR => \tok.keys.mem0_physical_WADDR_wire\,
            MASK => \tok.keys.mem0_physical_MASK_wire\,
            WDATA => \tok.keys.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__38455\,
            RE => \N__17528\,
            WCLKE => 'H',
            WCLK => \N__38456\,
            WE => \N__14632\
        );

    \tok.ram.mem2_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010001000001000000010000000100000101010001010101000101",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \tok.ram.mem2_physical_RDATA_wire\,
            RADDR => \tok.ram.mem2_physical_RADDR_wire\,
            WADDR => \tok.ram.mem2_physical_WADDR_wire\,
            MASK => \tok.ram.mem2_physical_MASK_wire\,
            WDATA => \tok.ram.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__38478\,
            RE => \N__17497\,
            WCLKE => 'H',
            WCLK => \N__38479\,
            WE => \N__30169\
        );

    \rx_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38690\,
            DIN => \N__38689\,
            DOUT => \N__38688\,
            PACKAGEPIN => rx_wire
        );

    \rx_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38690\,
            PADOUT => \N__38689\,
            PADIN => \N__38688\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => rx_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \reset_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38681\,
            DIN => \N__38680\,
            DOUT => \N__38679\,
            PACKAGEPIN => reset_wire
        );

    \reset_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38681\,
            PADOUT => \N__38680\,
            PADIN => \N__38679\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => reset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \tx_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38672\,
            DIN => \N__38671\,
            DOUT => \N__38670\,
            PACKAGEPIN => tx_wire
        );

    \tx_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38672\,
            PADOUT => \N__38671\,
            PADIN => \N__38670\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14953\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__9608\ : InMux
    port map (
            O => \N__38653\,
            I => \N__38646\
        );

    \I__9607\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38643\
        );

    \I__9606\ : InMux
    port map (
            O => \N__38651\,
            I => \N__38636\
        );

    \I__9605\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38636\
        );

    \I__9604\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38636\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__38646\,
            I => \tok.uart.bytephase_1\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__38643\,
            I => \tok.uart.bytephase_1\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__38636\,
            I => \tok.uart.bytephase_1\
        );

    \I__9600\ : InMux
    port map (
            O => \N__38629\,
            I => \N__38626\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__38626\,
            I => \N__38623\
        );

    \I__9598\ : Odrv4
    port map (
            O => \N__38623\,
            I => \tok.uart.n2357\
        );

    \I__9597\ : InMux
    port map (
            O => \N__38620\,
            I => \N__38616\
        );

    \I__9596\ : InMux
    port map (
            O => \N__38619\,
            I => \N__38613\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__38616\,
            I => \tok.uart.rxclkcounter_0\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__38613\,
            I => \tok.uart.rxclkcounter_0\
        );

    \I__9593\ : InMux
    port map (
            O => \N__38608\,
            I => \bfn_13_11_0_\
        );

    \I__9592\ : InMux
    port map (
            O => \N__38605\,
            I => \N__38601\
        );

    \I__9591\ : InMux
    port map (
            O => \N__38604\,
            I => \N__38598\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__38601\,
            I => \N__38595\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__38598\,
            I => \tok.uart.rxclkcounter_1\
        );

    \I__9588\ : Odrv4
    port map (
            O => \N__38595\,
            I => \tok.uart.rxclkcounter_1\
        );

    \I__9587\ : InMux
    port map (
            O => \N__38590\,
            I => \tok.uart.n4824\
        );

    \I__9586\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38583\
        );

    \I__9585\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38580\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__38583\,
            I => \tok.uart.rxclkcounter_2\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__38580\,
            I => \tok.uart.rxclkcounter_2\
        );

    \I__9582\ : InMux
    port map (
            O => \N__38575\,
            I => \tok.uart.n4825\
        );

    \I__9581\ : InMux
    port map (
            O => \N__38572\,
            I => \N__38568\
        );

    \I__9580\ : InMux
    port map (
            O => \N__38571\,
            I => \N__38565\
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__38568\,
            I => \tok.uart.rxclkcounter_3\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__38565\,
            I => \tok.uart.rxclkcounter_3\
        );

    \I__9577\ : InMux
    port map (
            O => \N__38560\,
            I => \tok.uart.n4826\
        );

    \I__9576\ : CascadeMux
    port map (
            O => \N__38557\,
            I => \N__38553\
        );

    \I__9575\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38550\
        );

    \I__9574\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38547\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__38550\,
            I => \tok.uart.rxclkcounter_4\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__38547\,
            I => \tok.uart.rxclkcounter_4\
        );

    \I__9571\ : InMux
    port map (
            O => \N__38542\,
            I => \tok.uart.n4827\
        );

    \I__9570\ : InMux
    port map (
            O => \N__38539\,
            I => \N__38535\
        );

    \I__9569\ : InMux
    port map (
            O => \N__38538\,
            I => \N__38532\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__38535\,
            I => \tok.uart.rxclkcounter_5\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__38532\,
            I => \tok.uart.rxclkcounter_5\
        );

    \I__9566\ : InMux
    port map (
            O => \N__38527\,
            I => \tok.uart.n4828\
        );

    \I__9565\ : InMux
    port map (
            O => \N__38524\,
            I => \tok.uart.n4829\
        );

    \I__9564\ : InMux
    port map (
            O => \N__38521\,
            I => \N__38517\
        );

    \I__9563\ : InMux
    port map (
            O => \N__38520\,
            I => \N__38514\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__38517\,
            I => \tok.uart.rxclkcounter_6\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__38514\,
            I => \tok.uart.rxclkcounter_6\
        );

    \I__9560\ : ClkMux
    port map (
            O => \N__38509\,
            I => \N__38257\
        );

    \I__9559\ : ClkMux
    port map (
            O => \N__38508\,
            I => \N__38257\
        );

    \I__9558\ : ClkMux
    port map (
            O => \N__38507\,
            I => \N__38257\
        );

    \I__9557\ : ClkMux
    port map (
            O => \N__38506\,
            I => \N__38257\
        );

    \I__9556\ : ClkMux
    port map (
            O => \N__38505\,
            I => \N__38257\
        );

    \I__9555\ : ClkMux
    port map (
            O => \N__38504\,
            I => \N__38257\
        );

    \I__9554\ : ClkMux
    port map (
            O => \N__38503\,
            I => \N__38257\
        );

    \I__9553\ : ClkMux
    port map (
            O => \N__38502\,
            I => \N__38257\
        );

    \I__9552\ : ClkMux
    port map (
            O => \N__38501\,
            I => \N__38257\
        );

    \I__9551\ : ClkMux
    port map (
            O => \N__38500\,
            I => \N__38257\
        );

    \I__9550\ : ClkMux
    port map (
            O => \N__38499\,
            I => \N__38257\
        );

    \I__9549\ : ClkMux
    port map (
            O => \N__38498\,
            I => \N__38257\
        );

    \I__9548\ : ClkMux
    port map (
            O => \N__38497\,
            I => \N__38257\
        );

    \I__9547\ : ClkMux
    port map (
            O => \N__38496\,
            I => \N__38257\
        );

    \I__9546\ : ClkMux
    port map (
            O => \N__38495\,
            I => \N__38257\
        );

    \I__9545\ : ClkMux
    port map (
            O => \N__38494\,
            I => \N__38257\
        );

    \I__9544\ : ClkMux
    port map (
            O => \N__38493\,
            I => \N__38257\
        );

    \I__9543\ : ClkMux
    port map (
            O => \N__38492\,
            I => \N__38257\
        );

    \I__9542\ : ClkMux
    port map (
            O => \N__38491\,
            I => \N__38257\
        );

    \I__9541\ : ClkMux
    port map (
            O => \N__38490\,
            I => \N__38257\
        );

    \I__9540\ : ClkMux
    port map (
            O => \N__38489\,
            I => \N__38257\
        );

    \I__9539\ : ClkMux
    port map (
            O => \N__38488\,
            I => \N__38257\
        );

    \I__9538\ : ClkMux
    port map (
            O => \N__38487\,
            I => \N__38257\
        );

    \I__9537\ : ClkMux
    port map (
            O => \N__38486\,
            I => \N__38257\
        );

    \I__9536\ : ClkMux
    port map (
            O => \N__38485\,
            I => \N__38257\
        );

    \I__9535\ : ClkMux
    port map (
            O => \N__38484\,
            I => \N__38257\
        );

    \I__9534\ : ClkMux
    port map (
            O => \N__38483\,
            I => \N__38257\
        );

    \I__9533\ : ClkMux
    port map (
            O => \N__38482\,
            I => \N__38257\
        );

    \I__9532\ : ClkMux
    port map (
            O => \N__38481\,
            I => \N__38257\
        );

    \I__9531\ : ClkMux
    port map (
            O => \N__38480\,
            I => \N__38257\
        );

    \I__9530\ : ClkMux
    port map (
            O => \N__38479\,
            I => \N__38257\
        );

    \I__9529\ : ClkMux
    port map (
            O => \N__38478\,
            I => \N__38257\
        );

    \I__9528\ : ClkMux
    port map (
            O => \N__38477\,
            I => \N__38257\
        );

    \I__9527\ : ClkMux
    port map (
            O => \N__38476\,
            I => \N__38257\
        );

    \I__9526\ : ClkMux
    port map (
            O => \N__38475\,
            I => \N__38257\
        );

    \I__9525\ : ClkMux
    port map (
            O => \N__38474\,
            I => \N__38257\
        );

    \I__9524\ : ClkMux
    port map (
            O => \N__38473\,
            I => \N__38257\
        );

    \I__9523\ : ClkMux
    port map (
            O => \N__38472\,
            I => \N__38257\
        );

    \I__9522\ : ClkMux
    port map (
            O => \N__38471\,
            I => \N__38257\
        );

    \I__9521\ : ClkMux
    port map (
            O => \N__38470\,
            I => \N__38257\
        );

    \I__9520\ : ClkMux
    port map (
            O => \N__38469\,
            I => \N__38257\
        );

    \I__9519\ : ClkMux
    port map (
            O => \N__38468\,
            I => \N__38257\
        );

    \I__9518\ : ClkMux
    port map (
            O => \N__38467\,
            I => \N__38257\
        );

    \I__9517\ : ClkMux
    port map (
            O => \N__38466\,
            I => \N__38257\
        );

    \I__9516\ : ClkMux
    port map (
            O => \N__38465\,
            I => \N__38257\
        );

    \I__9515\ : ClkMux
    port map (
            O => \N__38464\,
            I => \N__38257\
        );

    \I__9514\ : ClkMux
    port map (
            O => \N__38463\,
            I => \N__38257\
        );

    \I__9513\ : ClkMux
    port map (
            O => \N__38462\,
            I => \N__38257\
        );

    \I__9512\ : ClkMux
    port map (
            O => \N__38461\,
            I => \N__38257\
        );

    \I__9511\ : ClkMux
    port map (
            O => \N__38460\,
            I => \N__38257\
        );

    \I__9510\ : ClkMux
    port map (
            O => \N__38459\,
            I => \N__38257\
        );

    \I__9509\ : ClkMux
    port map (
            O => \N__38458\,
            I => \N__38257\
        );

    \I__9508\ : ClkMux
    port map (
            O => \N__38457\,
            I => \N__38257\
        );

    \I__9507\ : ClkMux
    port map (
            O => \N__38456\,
            I => \N__38257\
        );

    \I__9506\ : ClkMux
    port map (
            O => \N__38455\,
            I => \N__38257\
        );

    \I__9505\ : ClkMux
    port map (
            O => \N__38454\,
            I => \N__38257\
        );

    \I__9504\ : ClkMux
    port map (
            O => \N__38453\,
            I => \N__38257\
        );

    \I__9503\ : ClkMux
    port map (
            O => \N__38452\,
            I => \N__38257\
        );

    \I__9502\ : ClkMux
    port map (
            O => \N__38451\,
            I => \N__38257\
        );

    \I__9501\ : ClkMux
    port map (
            O => \N__38450\,
            I => \N__38257\
        );

    \I__9500\ : ClkMux
    port map (
            O => \N__38449\,
            I => \N__38257\
        );

    \I__9499\ : ClkMux
    port map (
            O => \N__38448\,
            I => \N__38257\
        );

    \I__9498\ : ClkMux
    port map (
            O => \N__38447\,
            I => \N__38257\
        );

    \I__9497\ : ClkMux
    port map (
            O => \N__38446\,
            I => \N__38257\
        );

    \I__9496\ : ClkMux
    port map (
            O => \N__38445\,
            I => \N__38257\
        );

    \I__9495\ : ClkMux
    port map (
            O => \N__38444\,
            I => \N__38257\
        );

    \I__9494\ : ClkMux
    port map (
            O => \N__38443\,
            I => \N__38257\
        );

    \I__9493\ : ClkMux
    port map (
            O => \N__38442\,
            I => \N__38257\
        );

    \I__9492\ : ClkMux
    port map (
            O => \N__38441\,
            I => \N__38257\
        );

    \I__9491\ : ClkMux
    port map (
            O => \N__38440\,
            I => \N__38257\
        );

    \I__9490\ : ClkMux
    port map (
            O => \N__38439\,
            I => \N__38257\
        );

    \I__9489\ : ClkMux
    port map (
            O => \N__38438\,
            I => \N__38257\
        );

    \I__9488\ : ClkMux
    port map (
            O => \N__38437\,
            I => \N__38257\
        );

    \I__9487\ : ClkMux
    port map (
            O => \N__38436\,
            I => \N__38257\
        );

    \I__9486\ : ClkMux
    port map (
            O => \N__38435\,
            I => \N__38257\
        );

    \I__9485\ : ClkMux
    port map (
            O => \N__38434\,
            I => \N__38257\
        );

    \I__9484\ : ClkMux
    port map (
            O => \N__38433\,
            I => \N__38257\
        );

    \I__9483\ : ClkMux
    port map (
            O => \N__38432\,
            I => \N__38257\
        );

    \I__9482\ : ClkMux
    port map (
            O => \N__38431\,
            I => \N__38257\
        );

    \I__9481\ : ClkMux
    port map (
            O => \N__38430\,
            I => \N__38257\
        );

    \I__9480\ : ClkMux
    port map (
            O => \N__38429\,
            I => \N__38257\
        );

    \I__9479\ : ClkMux
    port map (
            O => \N__38428\,
            I => \N__38257\
        );

    \I__9478\ : ClkMux
    port map (
            O => \N__38427\,
            I => \N__38257\
        );

    \I__9477\ : ClkMux
    port map (
            O => \N__38426\,
            I => \N__38257\
        );

    \I__9476\ : GlobalMux
    port map (
            O => \N__38257\,
            I => \N__38254\
        );

    \I__9475\ : DummyBuf
    port map (
            O => \N__38254\,
            I => clk
        );

    \I__9474\ : SRMux
    port map (
            O => \N__38251\,
            I => \N__38248\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38245\
        );

    \I__9472\ : Span4Mux_s0_h
    port map (
            O => \N__38245\,
            I => \N__38242\
        );

    \I__9471\ : Span4Mux_h
    port map (
            O => \N__38242\,
            I => \N__38239\
        );

    \I__9470\ : Odrv4
    port map (
            O => \N__38239\,
            I => \tok.uart.rxclkcounter_6__N_476\
        );

    \I__9469\ : InMux
    port map (
            O => \N__38236\,
            I => \tok.uart.n4823\
        );

    \I__9468\ : InMux
    port map (
            O => \N__38233\,
            I => \N__38228\
        );

    \I__9467\ : InMux
    port map (
            O => \N__38232\,
            I => \N__38223\
        );

    \I__9466\ : InMux
    port map (
            O => \N__38231\,
            I => \N__38223\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__38228\,
            I => \tok.uart.bytephase_5\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__38223\,
            I => \tok.uart.bytephase_5\
        );

    \I__9463\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38209\
        );

    \I__9462\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38209\
        );

    \I__9461\ : InMux
    port map (
            O => \N__38216\,
            I => \N__38198\
        );

    \I__9460\ : InMux
    port map (
            O => \N__38215\,
            I => \N__38198\
        );

    \I__9459\ : InMux
    port map (
            O => \N__38214\,
            I => \N__38198\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__38209\,
            I => \N__38195\
        );

    \I__9457\ : InMux
    port map (
            O => \N__38208\,
            I => \N__38192\
        );

    \I__9456\ : InMux
    port map (
            O => \N__38207\,
            I => \N__38185\
        );

    \I__9455\ : InMux
    port map (
            O => \N__38206\,
            I => \N__38185\
        );

    \I__9454\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38185\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__38198\,
            I => \N__38181\
        );

    \I__9452\ : Span4Mux_v
    port map (
            O => \N__38195\,
            I => \N__38174\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__38192\,
            I => \N__38174\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__38185\,
            I => \N__38174\
        );

    \I__9449\ : InMux
    port map (
            O => \N__38184\,
            I => \N__38171\
        );

    \I__9448\ : Odrv12
    port map (
            O => \N__38181\,
            I => n4928
        );

    \I__9447\ : Odrv4
    port map (
            O => \N__38174\,
            I => n4928
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__38171\,
            I => n4928
        );

    \I__9445\ : CascadeMux
    port map (
            O => \N__38164\,
            I => \tok.uart.n6_cascade_\
        );

    \I__9444\ : CascadeMux
    port map (
            O => \N__38161\,
            I => \n746_cascade_\
        );

    \I__9443\ : SRMux
    port map (
            O => \N__38158\,
            I => \N__38154\
        );

    \I__9442\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38151\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__38154\,
            I => \N__38148\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__38151\,
            I => \N__38145\
        );

    \I__9439\ : Odrv12
    port map (
            O => \N__38148\,
            I => \bytephase_5__N_509\
        );

    \I__9438\ : Odrv4
    port map (
            O => \N__38145\,
            I => \bytephase_5__N_509\
        );

    \I__9437\ : CEMux
    port map (
            O => \N__38140\,
            I => \N__38137\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__38137\,
            I => n974
        );

    \I__9435\ : InMux
    port map (
            O => \N__38134\,
            I => \N__38131\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__38131\,
            I => \tok.uart.n6211\
        );

    \I__9433\ : InMux
    port map (
            O => \N__38128\,
            I => \N__38125\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__38125\,
            I => \N__38122\
        );

    \I__9431\ : Odrv4
    port map (
            O => \N__38122\,
            I => \tok.uart.n2356\
        );

    \I__9430\ : InMux
    port map (
            O => \N__38119\,
            I => \N__38116\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__38116\,
            I => \N__38112\
        );

    \I__9428\ : InMux
    port map (
            O => \N__38115\,
            I => \N__38109\
        );

    \I__9427\ : Odrv12
    port map (
            O => \N__38112\,
            I => \tok.uart.n809\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__38109\,
            I => \tok.uart.n809\
        );

    \I__9425\ : CascadeMux
    port map (
            O => \N__38104\,
            I => \tok.uart.n2356_cascade_\
        );

    \I__9424\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38095\
        );

    \I__9423\ : InMux
    port map (
            O => \N__38100\,
            I => \N__38095\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__38095\,
            I => n746
        );

    \I__9421\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38087\
        );

    \I__9420\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38082\
        );

    \I__9419\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38082\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__38087\,
            I => \tok.uart.bytephase_2\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__38082\,
            I => \tok.uart.bytephase_2\
        );

    \I__9416\ : CascadeMux
    port map (
            O => \N__38077\,
            I => \N__38073\
        );

    \I__9415\ : InMux
    port map (
            O => \N__38076\,
            I => \N__38068\
        );

    \I__9414\ : InMux
    port map (
            O => \N__38073\,
            I => \N__38061\
        );

    \I__9413\ : InMux
    port map (
            O => \N__38072\,
            I => \N__38061\
        );

    \I__9412\ : InMux
    port map (
            O => \N__38071\,
            I => \N__38061\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__38068\,
            I => \tok.uart.bytephase_0\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__38061\,
            I => \tok.uart.bytephase_0\
        );

    \I__9409\ : CascadeMux
    port map (
            O => \N__38056\,
            I => \N__38052\
        );

    \I__9408\ : CascadeMux
    port map (
            O => \N__38055\,
            I => \N__38048\
        );

    \I__9407\ : InMux
    port map (
            O => \N__38052\,
            I => \N__38035\
        );

    \I__9406\ : InMux
    port map (
            O => \N__38051\,
            I => \N__38035\
        );

    \I__9405\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38035\
        );

    \I__9404\ : InMux
    port map (
            O => \N__38047\,
            I => \N__38035\
        );

    \I__9403\ : InMux
    port map (
            O => \N__38046\,
            I => \N__38035\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__38035\,
            I => \tok.uart.sentbits_0\
        );

    \I__9401\ : CEMux
    port map (
            O => \N__38032\,
            I => \N__38029\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__38029\,
            I => \N__38026\
        );

    \I__9399\ : Span4Mux_s0_h
    port map (
            O => \N__38026\,
            I => \N__38023\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__38023\,
            I => \tok.uart.n994\
        );

    \I__9397\ : SRMux
    port map (
            O => \N__38020\,
            I => \N__38017\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__38017\,
            I => \N__38014\
        );

    \I__9395\ : Odrv4
    port map (
            O => \N__38014\,
            I => \tok.uart.n1013\
        );

    \I__9394\ : CascadeMux
    port map (
            O => \N__38011\,
            I => \N__38007\
        );

    \I__9393\ : InMux
    port map (
            O => \N__38010\,
            I => \N__38004\
        );

    \I__9392\ : InMux
    port map (
            O => \N__38007\,
            I => \N__38001\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__38004\,
            I => \N__37996\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__38001\,
            I => \N__37996\
        );

    \I__9389\ : Span4Mux_v
    port map (
            O => \N__37996\,
            I => \N__37993\
        );

    \I__9388\ : Span4Mux_v
    port map (
            O => \N__37993\,
            I => \N__37990\
        );

    \I__9387\ : IoSpan4Mux
    port map (
            O => \N__37990\,
            I => \N__37987\
        );

    \I__9386\ : Odrv4
    port map (
            O => \N__37987\,
            I => rx_c
        );

    \I__9385\ : InMux
    port map (
            O => \N__37984\,
            I => \N__37981\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__37981\,
            I => \tok.uart.n4977\
        );

    \I__9383\ : CascadeMux
    port map (
            O => \N__37978\,
            I => \tok.uart.n4977_cascade_\
        );

    \I__9382\ : InMux
    port map (
            O => \N__37975\,
            I => \bfn_13_9_0_\
        );

    \I__9381\ : InMux
    port map (
            O => \N__37972\,
            I => \tok.uart.n4819\
        );

    \I__9380\ : InMux
    port map (
            O => \N__37969\,
            I => \tok.uart.n4820\
        );

    \I__9379\ : CascadeMux
    port map (
            O => \N__37966\,
            I => \N__37963\
        );

    \I__9378\ : InMux
    port map (
            O => \N__37963\,
            I => \N__37956\
        );

    \I__9377\ : InMux
    port map (
            O => \N__37962\,
            I => \N__37956\
        );

    \I__9376\ : InMux
    port map (
            O => \N__37961\,
            I => \N__37953\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__37956\,
            I => \N__37950\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__37953\,
            I => \tok.uart.bytephase_3\
        );

    \I__9373\ : Odrv4
    port map (
            O => \N__37950\,
            I => \tok.uart.bytephase_3\
        );

    \I__9372\ : InMux
    port map (
            O => \N__37945\,
            I => \tok.uart.n4821\
        );

    \I__9371\ : InMux
    port map (
            O => \N__37942\,
            I => \N__37937\
        );

    \I__9370\ : InMux
    port map (
            O => \N__37941\,
            I => \N__37932\
        );

    \I__9369\ : InMux
    port map (
            O => \N__37940\,
            I => \N__37932\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__37937\,
            I => \tok.uart.bytephase_4\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__37932\,
            I => \tok.uart.bytephase_4\
        );

    \I__9366\ : InMux
    port map (
            O => \N__37927\,
            I => \tok.uart.n4822\
        );

    \I__9365\ : InMux
    port map (
            O => \N__37924\,
            I => \N__37918\
        );

    \I__9364\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37918\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__37918\,
            I => capture_0
        );

    \I__9362\ : InMux
    port map (
            O => \N__37915\,
            I => \N__37912\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__37912\,
            I => \N__37907\
        );

    \I__9360\ : InMux
    port map (
            O => \N__37911\,
            I => \N__37904\
        );

    \I__9359\ : InMux
    port map (
            O => \N__37910\,
            I => \N__37901\
        );

    \I__9358\ : Odrv4
    port map (
            O => \N__37907\,
            I => capture_4
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__37904\,
            I => capture_4
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__37901\,
            I => capture_4
        );

    \I__9355\ : CascadeMux
    port map (
            O => \N__37894\,
            I => \rx_data_7__N_510_cascade_\
        );

    \I__9354\ : CascadeMux
    port map (
            O => \N__37891\,
            I => \N__37888\
        );

    \I__9353\ : InMux
    port map (
            O => \N__37888\,
            I => \N__37885\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__37885\,
            I => \N__37881\
        );

    \I__9351\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37878\
        );

    \I__9350\ : Span4Mux_h
    port map (
            O => \N__37881\,
            I => \N__37875\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__37878\,
            I => uart_rx_data_3
        );

    \I__9348\ : Odrv4
    port map (
            O => \N__37875\,
            I => uart_rx_data_3
        );

    \I__9347\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37865\
        );

    \I__9346\ : InMux
    port map (
            O => \N__37869\,
            I => \N__37860\
        );

    \I__9345\ : InMux
    port map (
            O => \N__37868\,
            I => \N__37860\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__37865\,
            I => capture_9
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__37860\,
            I => capture_9
        );

    \I__9342\ : InMux
    port map (
            O => \N__37855\,
            I => \N__37851\
        );

    \I__9341\ : CascadeMux
    port map (
            O => \N__37854\,
            I => \N__37848\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__37851\,
            I => \N__37844\
        );

    \I__9339\ : InMux
    port map (
            O => \N__37848\,
            I => \N__37839\
        );

    \I__9338\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37839\
        );

    \I__9337\ : Odrv4
    port map (
            O => \N__37844\,
            I => capture_6
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__37839\,
            I => capture_6
        );

    \I__9335\ : CascadeMux
    port map (
            O => \N__37834\,
            I => \N__37831\
        );

    \I__9334\ : InMux
    port map (
            O => \N__37831\,
            I => \N__37827\
        );

    \I__9333\ : InMux
    port map (
            O => \N__37830\,
            I => \N__37824\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__37827\,
            I => \N__37821\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__37824\,
            I => uart_rx_data_5
        );

    \I__9330\ : Odrv4
    port map (
            O => \N__37821\,
            I => uart_rx_data_5
        );

    \I__9329\ : InMux
    port map (
            O => \N__37816\,
            I => \N__37812\
        );

    \I__9328\ : InMux
    port map (
            O => \N__37815\,
            I => \N__37809\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__37812\,
            I => \N__37803\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__37809\,
            I => \N__37803\
        );

    \I__9325\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37800\
        );

    \I__9324\ : Odrv4
    port map (
            O => \N__37803\,
            I => capture_1
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__37800\,
            I => capture_1
        );

    \I__9322\ : InMux
    port map (
            O => \N__37795\,
            I => \N__37792\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__37792\,
            I => \N__37784\
        );

    \I__9320\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37781\
        );

    \I__9319\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37772\
        );

    \I__9318\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37772\
        );

    \I__9317\ : InMux
    port map (
            O => \N__37788\,
            I => \N__37772\
        );

    \I__9316\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37769\
        );

    \I__9315\ : Span4Mux_v
    port map (
            O => \N__37784\,
            I => \N__37764\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__37781\,
            I => \N__37764\
        );

    \I__9313\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37759\
        );

    \I__9312\ : InMux
    port map (
            O => \N__37779\,
            I => \N__37759\
        );

    \I__9311\ : LocalMux
    port map (
            O => \N__37772\,
            I => \N__37754\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__37769\,
            I => \N__37754\
        );

    \I__9309\ : Odrv4
    port map (
            O => \N__37764\,
            I => \rx_data_7__N_510\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__37759\,
            I => \rx_data_7__N_510\
        );

    \I__9307\ : Odrv4
    port map (
            O => \N__37754\,
            I => \rx_data_7__N_510\
        );

    \I__9306\ : CascadeMux
    port map (
            O => \N__37747\,
            I => \N__37744\
        );

    \I__9305\ : InMux
    port map (
            O => \N__37744\,
            I => \N__37741\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__37741\,
            I => \N__37738\
        );

    \I__9303\ : Span4Mux_h
    port map (
            O => \N__37738\,
            I => \N__37734\
        );

    \I__9302\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37731\
        );

    \I__9301\ : Span4Mux_h
    port map (
            O => \N__37734\,
            I => \N__37728\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__37731\,
            I => uart_rx_data_0
        );

    \I__9299\ : Odrv4
    port map (
            O => \N__37728\,
            I => uart_rx_data_0
        );

    \I__9298\ : InMux
    port map (
            O => \N__37723\,
            I => \N__37711\
        );

    \I__9297\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37711\
        );

    \I__9296\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37711\
        );

    \I__9295\ : InMux
    port map (
            O => \N__37720\,
            I => \N__37711\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__37711\,
            I => \tok.uart_tx_busy\
        );

    \I__9293\ : InMux
    port map (
            O => \N__37708\,
            I => \N__37702\
        );

    \I__9292\ : InMux
    port map (
            O => \N__37707\,
            I => \N__37702\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__37702\,
            I => \tok.uart.sentbits_3\
        );

    \I__9290\ : CascadeMux
    port map (
            O => \N__37699\,
            I => \N__37694\
        );

    \I__9289\ : InMux
    port map (
            O => \N__37698\,
            I => \N__37687\
        );

    \I__9288\ : InMux
    port map (
            O => \N__37697\,
            I => \N__37687\
        );

    \I__9287\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37687\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__37687\,
            I => \tok.uart.sentbits_2\
        );

    \I__9285\ : InMux
    port map (
            O => \N__37684\,
            I => \N__37672\
        );

    \I__9284\ : InMux
    port map (
            O => \N__37683\,
            I => \N__37672\
        );

    \I__9283\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37672\
        );

    \I__9282\ : InMux
    port map (
            O => \N__37681\,
            I => \N__37672\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__37672\,
            I => \tok.uart.sentbits_1\
        );

    \I__9280\ : InMux
    port map (
            O => \N__37669\,
            I => \N__37665\
        );

    \I__9279\ : InMux
    port map (
            O => \N__37668\,
            I => \N__37662\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__37665\,
            I => \N__37658\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__37662\,
            I => \N__37655\
        );

    \I__9276\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37652\
        );

    \I__9275\ : Odrv12
    port map (
            O => \N__37658\,
            I => capture_8
        );

    \I__9274\ : Odrv4
    port map (
            O => \N__37655\,
            I => capture_8
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__37652\,
            I => capture_8
        );

    \I__9272\ : CascadeMux
    port map (
            O => \N__37645\,
            I => \N__37642\
        );

    \I__9271\ : InMux
    port map (
            O => \N__37642\,
            I => \N__37638\
        );

    \I__9270\ : InMux
    port map (
            O => \N__37641\,
            I => \N__37635\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__37638\,
            I => \N__37632\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__37635\,
            I => uart_rx_data_7
        );

    \I__9267\ : Odrv4
    port map (
            O => \N__37632\,
            I => uart_rx_data_7
        );

    \I__9266\ : InMux
    port map (
            O => \N__37627\,
            I => \N__37624\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__37624\,
            I => \N__37620\
        );

    \I__9264\ : CascadeMux
    port map (
            O => \N__37623\,
            I => \N__37617\
        );

    \I__9263\ : Span4Mux_s2_v
    port map (
            O => \N__37620\,
            I => \N__37613\
        );

    \I__9262\ : InMux
    port map (
            O => \N__37617\,
            I => \N__37608\
        );

    \I__9261\ : InMux
    port map (
            O => \N__37616\,
            I => \N__37608\
        );

    \I__9260\ : Span4Mux_v
    port map (
            O => \N__37613\,
            I => \N__37602\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__37608\,
            I => \N__37602\
        );

    \I__9258\ : SRMux
    port map (
            O => \N__37607\,
            I => \N__37598\
        );

    \I__9257\ : Span4Mux_h
    port map (
            O => \N__37602\,
            I => \N__37595\
        );

    \I__9256\ : SRMux
    port map (
            O => \N__37601\,
            I => \N__37592\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__37598\,
            I => \N__37588\
        );

    \I__9254\ : Span4Mux_h
    port map (
            O => \N__37595\,
            I => \N__37585\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__37592\,
            I => \N__37582\
        );

    \I__9252\ : InMux
    port map (
            O => \N__37591\,
            I => \N__37579\
        );

    \I__9251\ : Span4Mux_s2_v
    port map (
            O => \N__37588\,
            I => \N__37574\
        );

    \I__9250\ : Span4Mux_h
    port map (
            O => \N__37585\,
            I => \N__37574\
        );

    \I__9249\ : Odrv4
    port map (
            O => \N__37582\,
            I => txtick
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__37579\,
            I => txtick
        );

    \I__9247\ : Odrv4
    port map (
            O => \N__37574\,
            I => txtick
        );

    \I__9246\ : CascadeMux
    port map (
            O => \N__37567\,
            I => \N__37562\
        );

    \I__9245\ : SRMux
    port map (
            O => \N__37566\,
            I => \N__37558\
        );

    \I__9244\ : InMux
    port map (
            O => \N__37565\,
            I => \N__37549\
        );

    \I__9243\ : InMux
    port map (
            O => \N__37562\,
            I => \N__37549\
        );

    \I__9242\ : InMux
    port map (
            O => \N__37561\,
            I => \N__37549\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__37558\,
            I => \N__37546\
        );

    \I__9240\ : InMux
    port map (
            O => \N__37557\,
            I => \N__37541\
        );

    \I__9239\ : InMux
    port map (
            O => \N__37556\,
            I => \N__37541\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__37549\,
            I => \N__37537\
        );

    \I__9237\ : Span4Mux_s2_v
    port map (
            O => \N__37546\,
            I => \N__37529\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__37541\,
            I => \N__37529\
        );

    \I__9235\ : InMux
    port map (
            O => \N__37540\,
            I => \N__37526\
        );

    \I__9234\ : Span4Mux_v
    port map (
            O => \N__37537\,
            I => \N__37523\
        );

    \I__9233\ : InMux
    port map (
            O => \N__37536\,
            I => \N__37516\
        );

    \I__9232\ : InMux
    port map (
            O => \N__37535\,
            I => \N__37516\
        );

    \I__9231\ : InMux
    port map (
            O => \N__37534\,
            I => \N__37516\
        );

    \I__9230\ : Span4Mux_v
    port map (
            O => \N__37529\,
            I => \N__37512\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__37526\,
            I => \N__37509\
        );

    \I__9228\ : Span4Mux_h
    port map (
            O => \N__37523\,
            I => \N__37504\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__37516\,
            I => \N__37504\
        );

    \I__9226\ : InMux
    port map (
            O => \N__37515\,
            I => \N__37501\
        );

    \I__9225\ : Span4Mux_h
    port map (
            O => \N__37512\,
            I => \N__37497\
        );

    \I__9224\ : Span12Mux_h
    port map (
            O => \N__37509\,
            I => \N__37490\
        );

    \I__9223\ : Sp12to4
    port map (
            O => \N__37504\,
            I => \N__37490\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__37501\,
            I => \N__37490\
        );

    \I__9221\ : InMux
    port map (
            O => \N__37500\,
            I => \N__37487\
        );

    \I__9220\ : Span4Mux_h
    port map (
            O => \N__37497\,
            I => \N__37484\
        );

    \I__9219\ : Odrv12
    port map (
            O => \N__37490\,
            I => n23
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__37487\,
            I => n23
        );

    \I__9217\ : Odrv4
    port map (
            O => \N__37484\,
            I => n23
        );

    \I__9216\ : InMux
    port map (
            O => \N__37477\,
            I => \N__37471\
        );

    \I__9215\ : InMux
    port map (
            O => \N__37476\,
            I => \N__37460\
        );

    \I__9214\ : InMux
    port map (
            O => \N__37475\,
            I => \N__37460\
        );

    \I__9213\ : InMux
    port map (
            O => \N__37474\,
            I => \N__37457\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__37471\,
            I => \N__37452\
        );

    \I__9211\ : InMux
    port map (
            O => \N__37470\,
            I => \N__37449\
        );

    \I__9210\ : CascadeMux
    port map (
            O => \N__37469\,
            I => \N__37446\
        );

    \I__9209\ : InMux
    port map (
            O => \N__37468\,
            I => \N__37439\
        );

    \I__9208\ : InMux
    port map (
            O => \N__37467\,
            I => \N__37436\
        );

    \I__9207\ : CascadeMux
    port map (
            O => \N__37466\,
            I => \N__37433\
        );

    \I__9206\ : InMux
    port map (
            O => \N__37465\,
            I => \N__37430\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__37460\,
            I => \N__37427\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__37457\,
            I => \N__37424\
        );

    \I__9203\ : InMux
    port map (
            O => \N__37456\,
            I => \N__37419\
        );

    \I__9202\ : InMux
    port map (
            O => \N__37455\,
            I => \N__37419\
        );

    \I__9201\ : Span4Mux_s0_v
    port map (
            O => \N__37452\,
            I => \N__37416\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__37449\,
            I => \N__37413\
        );

    \I__9199\ : InMux
    port map (
            O => \N__37446\,
            I => \N__37406\
        );

    \I__9198\ : InMux
    port map (
            O => \N__37445\,
            I => \N__37406\
        );

    \I__9197\ : InMux
    port map (
            O => \N__37444\,
            I => \N__37406\
        );

    \I__9196\ : InMux
    port map (
            O => \N__37443\,
            I => \N__37403\
        );

    \I__9195\ : InMux
    port map (
            O => \N__37442\,
            I => \N__37397\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__37439\,
            I => \N__37394\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__37436\,
            I => \N__37391\
        );

    \I__9192\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37388\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__37430\,
            I => \N__37383\
        );

    \I__9190\ : Span4Mux_s1_h
    port map (
            O => \N__37427\,
            I => \N__37380\
        );

    \I__9189\ : Span4Mux_s3_v
    port map (
            O => \N__37424\,
            I => \N__37375\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__37419\,
            I => \N__37375\
        );

    \I__9187\ : Span4Mux_v
    port map (
            O => \N__37416\,
            I => \N__37372\
        );

    \I__9186\ : Span4Mux_s1_v
    port map (
            O => \N__37413\,
            I => \N__37365\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__37406\,
            I => \N__37365\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__37403\,
            I => \N__37365\
        );

    \I__9183\ : InMux
    port map (
            O => \N__37402\,
            I => \N__37360\
        );

    \I__9182\ : InMux
    port map (
            O => \N__37401\,
            I => \N__37360\
        );

    \I__9181\ : CascadeMux
    port map (
            O => \N__37400\,
            I => \N__37356\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__37397\,
            I => \N__37349\
        );

    \I__9179\ : Span4Mux_v
    port map (
            O => \N__37394\,
            I => \N__37349\
        );

    \I__9178\ : Span4Mux_v
    port map (
            O => \N__37391\,
            I => \N__37349\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__37388\,
            I => \N__37346\
        );

    \I__9176\ : InMux
    port map (
            O => \N__37387\,
            I => \N__37341\
        );

    \I__9175\ : InMux
    port map (
            O => \N__37386\,
            I => \N__37341\
        );

    \I__9174\ : Span4Mux_s3_v
    port map (
            O => \N__37383\,
            I => \N__37334\
        );

    \I__9173\ : Span4Mux_h
    port map (
            O => \N__37380\,
            I => \N__37334\
        );

    \I__9172\ : Span4Mux_h
    port map (
            O => \N__37375\,
            I => \N__37334\
        );

    \I__9171\ : Span4Mux_v
    port map (
            O => \N__37372\,
            I => \N__37329\
        );

    \I__9170\ : Span4Mux_v
    port map (
            O => \N__37365\,
            I => \N__37329\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__37360\,
            I => \N__37326\
        );

    \I__9168\ : InMux
    port map (
            O => \N__37359\,
            I => \N__37321\
        );

    \I__9167\ : InMux
    port map (
            O => \N__37356\,
            I => \N__37321\
        );

    \I__9166\ : Span4Mux_h
    port map (
            O => \N__37349\,
            I => \N__37316\
        );

    \I__9165\ : Span4Mux_h
    port map (
            O => \N__37346\,
            I => \N__37316\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__37341\,
            I => \A_low_7\
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__37334\,
            I => \A_low_7\
        );

    \I__9162\ : Odrv4
    port map (
            O => \N__37329\,
            I => \A_low_7\
        );

    \I__9161\ : Odrv12
    port map (
            O => \N__37326\,
            I => \A_low_7\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__37321\,
            I => \A_low_7\
        );

    \I__9159\ : Odrv4
    port map (
            O => \N__37316\,
            I => \A_low_7\
        );

    \I__9158\ : CascadeMux
    port map (
            O => \N__37303\,
            I => \N__37300\
        );

    \I__9157\ : InMux
    port map (
            O => \N__37300\,
            I => \N__37296\
        );

    \I__9156\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37293\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__37296\,
            I => sender_9
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__37293\,
            I => sender_9
        );

    \I__9153\ : CascadeMux
    port map (
            O => \N__37288\,
            I => \N__37285\
        );

    \I__9152\ : InMux
    port map (
            O => \N__37285\,
            I => \N__37278\
        );

    \I__9151\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37278\
        );

    \I__9150\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37275\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__37278\,
            I => capture_3
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__37275\,
            I => capture_3
        );

    \I__9147\ : InMux
    port map (
            O => \N__37270\,
            I => \N__37267\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__37267\,
            I => \N__37262\
        );

    \I__9145\ : InMux
    port map (
            O => \N__37266\,
            I => \N__37257\
        );

    \I__9144\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37257\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__37262\,
            I => capture_5
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__37257\,
            I => capture_5
        );

    \I__9141\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37249\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__37249\,
            I => \N__37246\
        );

    \I__9139\ : Span4Mux_s0_h
    port map (
            O => \N__37246\,
            I => \N__37243\
        );

    \I__9138\ : Span4Mux_h
    port map (
            O => \N__37243\,
            I => \N__37238\
        );

    \I__9137\ : InMux
    port map (
            O => \N__37242\,
            I => \N__37235\
        );

    \I__9136\ : CascadeMux
    port map (
            O => \N__37241\,
            I => \N__37231\
        );

    \I__9135\ : Span4Mux_h
    port map (
            O => \N__37238\,
            I => \N__37227\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__37235\,
            I => \N__37224\
        );

    \I__9133\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37221\
        );

    \I__9132\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37216\
        );

    \I__9131\ : InMux
    port map (
            O => \N__37230\,
            I => \N__37216\
        );

    \I__9130\ : Odrv4
    port map (
            O => \N__37227\,
            I => \tok.n891\
        );

    \I__9129\ : Odrv12
    port map (
            O => \N__37224\,
            I => \tok.n891\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__37221\,
            I => \tok.n891\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__37216\,
            I => \tok.n891\
        );

    \I__9126\ : CascadeMux
    port map (
            O => \N__37207\,
            I => \N__37204\
        );

    \I__9125\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37195\
        );

    \I__9124\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37195\
        );

    \I__9123\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37195\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__37195\,
            I => \N__37192\
        );

    \I__9121\ : Span4Mux_h
    port map (
            O => \N__37192\,
            I => \N__37187\
        );

    \I__9120\ : InMux
    port map (
            O => \N__37191\,
            I => \N__37184\
        );

    \I__9119\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37181\
        );

    \I__9118\ : Span4Mux_h
    port map (
            O => \N__37187\,
            I => \N__37178\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__37184\,
            I => \tok.uart_rx_valid\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__37181\,
            I => \tok.uart_rx_valid\
        );

    \I__9115\ : Odrv4
    port map (
            O => \N__37178\,
            I => \tok.uart_rx_valid\
        );

    \I__9114\ : CEMux
    port map (
            O => \N__37171\,
            I => \N__37168\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__37168\,
            I => \N__37165\
        );

    \I__9112\ : Sp12to4
    port map (
            O => \N__37165\,
            I => \N__37162\
        );

    \I__9111\ : Odrv12
    port map (
            O => \N__37162\,
            I => \tok.uart.n922\
        );

    \I__9110\ : InMux
    port map (
            O => \N__37159\,
            I => \N__37156\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__37156\,
            I => \N__37153\
        );

    \I__9108\ : Span4Mux_v
    port map (
            O => \N__37153\,
            I => \N__37148\
        );

    \I__9107\ : InMux
    port map (
            O => \N__37152\,
            I => \N__37143\
        );

    \I__9106\ : InMux
    port map (
            O => \N__37151\,
            I => \N__37143\
        );

    \I__9105\ : Odrv4
    port map (
            O => \N__37148\,
            I => capture_7
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__37143\,
            I => capture_7
        );

    \I__9103\ : CascadeMux
    port map (
            O => \N__37138\,
            I => \N__37131\
        );

    \I__9102\ : InMux
    port map (
            O => \N__37137\,
            I => \N__37117\
        );

    \I__9101\ : InMux
    port map (
            O => \N__37136\,
            I => \N__37117\
        );

    \I__9100\ : CascadeMux
    port map (
            O => \N__37135\,
            I => \N__37114\
        );

    \I__9099\ : InMux
    port map (
            O => \N__37134\,
            I => \N__37107\
        );

    \I__9098\ : InMux
    port map (
            O => \N__37131\,
            I => \N__37100\
        );

    \I__9097\ : InMux
    port map (
            O => \N__37130\,
            I => \N__37100\
        );

    \I__9096\ : InMux
    port map (
            O => \N__37129\,
            I => \N__37100\
        );

    \I__9095\ : CascadeMux
    port map (
            O => \N__37128\,
            I => \N__37088\
        );

    \I__9094\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37079\
        );

    \I__9093\ : CascadeMux
    port map (
            O => \N__37126\,
            I => \N__37070\
        );

    \I__9092\ : InMux
    port map (
            O => \N__37125\,
            I => \N__37058\
        );

    \I__9091\ : InMux
    port map (
            O => \N__37124\,
            I => \N__37058\
        );

    \I__9090\ : InMux
    port map (
            O => \N__37123\,
            I => \N__37053\
        );

    \I__9089\ : InMux
    port map (
            O => \N__37122\,
            I => \N__37053\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__37117\,
            I => \N__37050\
        );

    \I__9087\ : InMux
    port map (
            O => \N__37114\,
            I => \N__37047\
        );

    \I__9086\ : InMux
    port map (
            O => \N__37113\,
            I => \N__37039\
        );

    \I__9085\ : InMux
    port map (
            O => \N__37112\,
            I => \N__37034\
        );

    \I__9084\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37034\
        );

    \I__9083\ : InMux
    port map (
            O => \N__37110\,
            I => \N__37031\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__37107\,
            I => \N__37026\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__37100\,
            I => \N__37026\
        );

    \I__9080\ : CascadeMux
    port map (
            O => \N__37099\,
            I => \N__37023\
        );

    \I__9079\ : InMux
    port map (
            O => \N__37098\,
            I => \N__37018\
        );

    \I__9078\ : InMux
    port map (
            O => \N__37097\,
            I => \N__37018\
        );

    \I__9077\ : InMux
    port map (
            O => \N__37096\,
            I => \N__37011\
        );

    \I__9076\ : InMux
    port map (
            O => \N__37095\,
            I => \N__37011\
        );

    \I__9075\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37011\
        );

    \I__9074\ : InMux
    port map (
            O => \N__37093\,
            I => \N__37004\
        );

    \I__9073\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37004\
        );

    \I__9072\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37004\
        );

    \I__9071\ : InMux
    port map (
            O => \N__37088\,
            I => \N__36994\
        );

    \I__9070\ : InMux
    port map (
            O => \N__37087\,
            I => \N__36994\
        );

    \I__9069\ : InMux
    port map (
            O => \N__37086\,
            I => \N__36994\
        );

    \I__9068\ : InMux
    port map (
            O => \N__37085\,
            I => \N__36989\
        );

    \I__9067\ : InMux
    port map (
            O => \N__37084\,
            I => \N__36989\
        );

    \I__9066\ : InMux
    port map (
            O => \N__37083\,
            I => \N__36973\
        );

    \I__9065\ : InMux
    port map (
            O => \N__37082\,
            I => \N__36973\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__37079\,
            I => \N__36970\
        );

    \I__9063\ : InMux
    port map (
            O => \N__37078\,
            I => \N__36959\
        );

    \I__9062\ : InMux
    port map (
            O => \N__37077\,
            I => \N__36959\
        );

    \I__9061\ : InMux
    port map (
            O => \N__37076\,
            I => \N__36959\
        );

    \I__9060\ : InMux
    port map (
            O => \N__37075\,
            I => \N__36959\
        );

    \I__9059\ : InMux
    port map (
            O => \N__37074\,
            I => \N__36959\
        );

    \I__9058\ : InMux
    port map (
            O => \N__37073\,
            I => \N__36942\
        );

    \I__9057\ : InMux
    port map (
            O => \N__37070\,
            I => \N__36937\
        );

    \I__9056\ : InMux
    port map (
            O => \N__37069\,
            I => \N__36937\
        );

    \I__9055\ : InMux
    port map (
            O => \N__37068\,
            I => \N__36932\
        );

    \I__9054\ : InMux
    port map (
            O => \N__37067\,
            I => \N__36929\
        );

    \I__9053\ : InMux
    port map (
            O => \N__37066\,
            I => \N__36926\
        );

    \I__9052\ : InMux
    port map (
            O => \N__37065\,
            I => \N__36923\
        );

    \I__9051\ : InMux
    port map (
            O => \N__37064\,
            I => \N__36918\
        );

    \I__9050\ : InMux
    port map (
            O => \N__37063\,
            I => \N__36918\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__37058\,
            I => \N__36909\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__37053\,
            I => \N__36909\
        );

    \I__9047\ : Span4Mux_h
    port map (
            O => \N__37050\,
            I => \N__36909\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__37047\,
            I => \N__36909\
        );

    \I__9045\ : InMux
    port map (
            O => \N__37046\,
            I => \N__36904\
        );

    \I__9044\ : InMux
    port map (
            O => \N__37045\,
            I => \N__36904\
        );

    \I__9043\ : InMux
    port map (
            O => \N__37044\,
            I => \N__36901\
        );

    \I__9042\ : InMux
    port map (
            O => \N__37043\,
            I => \N__36898\
        );

    \I__9041\ : InMux
    port map (
            O => \N__37042\,
            I => \N__36894\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__37039\,
            I => \N__36889\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__37034\,
            I => \N__36889\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__37031\,
            I => \N__36884\
        );

    \I__9037\ : Span4Mux_v
    port map (
            O => \N__37026\,
            I => \N__36884\
        );

    \I__9036\ : InMux
    port map (
            O => \N__37023\,
            I => \N__36881\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__37018\,
            I => \N__36874\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__37011\,
            I => \N__36874\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__37004\,
            I => \N__36874\
        );

    \I__9032\ : InMux
    port map (
            O => \N__37003\,
            I => \N__36867\
        );

    \I__9031\ : InMux
    port map (
            O => \N__37002\,
            I => \N__36867\
        );

    \I__9030\ : InMux
    port map (
            O => \N__37001\,
            I => \N__36867\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__36994\,
            I => \N__36862\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__36989\,
            I => \N__36862\
        );

    \I__9027\ : InMux
    port map (
            O => \N__36988\,
            I => \N__36853\
        );

    \I__9026\ : InMux
    port map (
            O => \N__36987\,
            I => \N__36853\
        );

    \I__9025\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36853\
        );

    \I__9024\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36853\
        );

    \I__9023\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36845\
        );

    \I__9022\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36845\
        );

    \I__9021\ : InMux
    port map (
            O => \N__36982\,
            I => \N__36845\
        );

    \I__9020\ : InMux
    port map (
            O => \N__36981\,
            I => \N__36842\
        );

    \I__9019\ : CascadeMux
    port map (
            O => \N__36980\,
            I => \N__36838\
        );

    \I__9018\ : InMux
    port map (
            O => \N__36979\,
            I => \N__36833\
        );

    \I__9017\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36833\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__36973\,
            I => \N__36826\
        );

    \I__9015\ : Span4Mux_h
    port map (
            O => \N__36970\,
            I => \N__36826\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__36959\,
            I => \N__36826\
        );

    \I__9013\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36819\
        );

    \I__9012\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36819\
        );

    \I__9011\ : InMux
    port map (
            O => \N__36956\,
            I => \N__36819\
        );

    \I__9010\ : InMux
    port map (
            O => \N__36955\,
            I => \N__36810\
        );

    \I__9009\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36810\
        );

    \I__9008\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36810\
        );

    \I__9007\ : InMux
    port map (
            O => \N__36952\,
            I => \N__36810\
        );

    \I__9006\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36805\
        );

    \I__9005\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36805\
        );

    \I__9004\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36798\
        );

    \I__9003\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36798\
        );

    \I__9002\ : InMux
    port map (
            O => \N__36947\,
            I => \N__36798\
        );

    \I__9001\ : InMux
    port map (
            O => \N__36946\,
            I => \N__36790\
        );

    \I__9000\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36790\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__36942\,
            I => \N__36785\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__36937\,
            I => \N__36785\
        );

    \I__8997\ : CascadeMux
    port map (
            O => \N__36936\,
            I => \N__36781\
        );

    \I__8996\ : CascadeMux
    port map (
            O => \N__36935\,
            I => \N__36777\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__36932\,
            I => \N__36774\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__36929\,
            I => \N__36771\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__36926\,
            I => \N__36768\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__36923\,
            I => \N__36759\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__36918\,
            I => \N__36759\
        );

    \I__8990\ : Span4Mux_v
    port map (
            O => \N__36909\,
            I => \N__36759\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__36904\,
            I => \N__36759\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__36901\,
            I => \N__36754\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__36898\,
            I => \N__36754\
        );

    \I__8986\ : InMux
    port map (
            O => \N__36897\,
            I => \N__36750\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__36894\,
            I => \N__36733\
        );

    \I__8984\ : Span4Mux_v
    port map (
            O => \N__36889\,
            I => \N__36733\
        );

    \I__8983\ : Span4Mux_h
    port map (
            O => \N__36884\,
            I => \N__36733\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__36881\,
            I => \N__36733\
        );

    \I__8981\ : Span4Mux_h
    port map (
            O => \N__36874\,
            I => \N__36733\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__36867\,
            I => \N__36733\
        );

    \I__8979\ : Span4Mux_v
    port map (
            O => \N__36862\,
            I => \N__36728\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__36853\,
            I => \N__36728\
        );

    \I__8977\ : InMux
    port map (
            O => \N__36852\,
            I => \N__36724\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__36845\,
            I => \N__36719\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__36842\,
            I => \N__36719\
        );

    \I__8974\ : InMux
    port map (
            O => \N__36841\,
            I => \N__36716\
        );

    \I__8973\ : InMux
    port map (
            O => \N__36838\,
            I => \N__36713\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__36833\,
            I => \N__36704\
        );

    \I__8971\ : Sp12to4
    port map (
            O => \N__36826\,
            I => \N__36704\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__36819\,
            I => \N__36704\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__36810\,
            I => \N__36704\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__36805\,
            I => \N__36699\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__36798\,
            I => \N__36699\
        );

    \I__8966\ : InMux
    port map (
            O => \N__36797\,
            I => \N__36694\
        );

    \I__8965\ : InMux
    port map (
            O => \N__36796\,
            I => \N__36689\
        );

    \I__8964\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36689\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__36790\,
            I => \N__36686\
        );

    \I__8962\ : Span4Mux_v
    port map (
            O => \N__36785\,
            I => \N__36683\
        );

    \I__8961\ : InMux
    port map (
            O => \N__36784\,
            I => \N__36678\
        );

    \I__8960\ : InMux
    port map (
            O => \N__36781\,
            I => \N__36678\
        );

    \I__8959\ : InMux
    port map (
            O => \N__36780\,
            I => \N__36673\
        );

    \I__8958\ : InMux
    port map (
            O => \N__36777\,
            I => \N__36673\
        );

    \I__8957\ : Span4Mux_v
    port map (
            O => \N__36774\,
            I => \N__36662\
        );

    \I__8956\ : Span4Mux_s3_v
    port map (
            O => \N__36771\,
            I => \N__36662\
        );

    \I__8955\ : Span4Mux_s3_v
    port map (
            O => \N__36768\,
            I => \N__36662\
        );

    \I__8954\ : Span4Mux_s3_v
    port map (
            O => \N__36759\,
            I => \N__36662\
        );

    \I__8953\ : Span4Mux_v
    port map (
            O => \N__36754\,
            I => \N__36662\
        );

    \I__8952\ : InMux
    port map (
            O => \N__36753\,
            I => \N__36659\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__36750\,
            I => \N__36656\
        );

    \I__8950\ : InMux
    port map (
            O => \N__36749\,
            I => \N__36647\
        );

    \I__8949\ : InMux
    port map (
            O => \N__36748\,
            I => \N__36647\
        );

    \I__8948\ : InMux
    port map (
            O => \N__36747\,
            I => \N__36647\
        );

    \I__8947\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36647\
        );

    \I__8946\ : Span4Mux_h
    port map (
            O => \N__36733\,
            I => \N__36644\
        );

    \I__8945\ : Span4Mux_h
    port map (
            O => \N__36728\,
            I => \N__36641\
        );

    \I__8944\ : CascadeMux
    port map (
            O => \N__36727\,
            I => \N__36638\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__36724\,
            I => \N__36635\
        );

    \I__8942\ : Span4Mux_s3_h
    port map (
            O => \N__36719\,
            I => \N__36632\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__36716\,
            I => \N__36627\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__36713\,
            I => \N__36627\
        );

    \I__8939\ : Span12Mux_s3_v
    port map (
            O => \N__36704\,
            I => \N__36622\
        );

    \I__8938\ : Span12Mux_s10_v
    port map (
            O => \N__36699\,
            I => \N__36622\
        );

    \I__8937\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36617\
        );

    \I__8936\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36617\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__36694\,
            I => \N__36596\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36596\
        );

    \I__8933\ : Span12Mux_s3_v
    port map (
            O => \N__36686\,
            I => \N__36596\
        );

    \I__8932\ : Sp12to4
    port map (
            O => \N__36683\,
            I => \N__36596\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__36678\,
            I => \N__36596\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__36673\,
            I => \N__36596\
        );

    \I__8929\ : Sp12to4
    port map (
            O => \N__36662\,
            I => \N__36596\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__36659\,
            I => \N__36596\
        );

    \I__8927\ : Span12Mux_s2_h
    port map (
            O => \N__36656\,
            I => \N__36596\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__36647\,
            I => \N__36596\
        );

    \I__8925\ : Span4Mux_v
    port map (
            O => \N__36644\,
            I => \N__36591\
        );

    \I__8924\ : Span4Mux_h
    port map (
            O => \N__36641\,
            I => \N__36591\
        );

    \I__8923\ : InMux
    port map (
            O => \N__36638\,
            I => \N__36588\
        );

    \I__8922\ : Odrv4
    port map (
            O => \N__36635\,
            I => \tok.T_5\
        );

    \I__8921\ : Odrv4
    port map (
            O => \N__36632\,
            I => \tok.T_5\
        );

    \I__8920\ : Odrv4
    port map (
            O => \N__36627\,
            I => \tok.T_5\
        );

    \I__8919\ : Odrv12
    port map (
            O => \N__36622\,
            I => \tok.T_5\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__36617\,
            I => \tok.T_5\
        );

    \I__8917\ : Odrv12
    port map (
            O => \N__36596\,
            I => \tok.T_5\
        );

    \I__8916\ : Odrv4
    port map (
            O => \N__36591\,
            I => \tok.T_5\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__36588\,
            I => \tok.T_5\
        );

    \I__8914\ : InMux
    port map (
            O => \N__36571\,
            I => \N__36568\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__36568\,
            I => \N__36565\
        );

    \I__8912\ : Span4Mux_h
    port map (
            O => \N__36565\,
            I => \N__36562\
        );

    \I__8911\ : Odrv4
    port map (
            O => \N__36562\,
            I => \tok.n317\
        );

    \I__8910\ : CascadeMux
    port map (
            O => \N__36559\,
            I => \tok.n317_cascade_\
        );

    \I__8909\ : CascadeMux
    port map (
            O => \N__36556\,
            I => \N__36550\
        );

    \I__8908\ : InMux
    port map (
            O => \N__36555\,
            I => \N__36545\
        );

    \I__8907\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36542\
        );

    \I__8906\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36536\
        );

    \I__8905\ : InMux
    port map (
            O => \N__36550\,
            I => \N__36536\
        );

    \I__8904\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36529\
        );

    \I__8903\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36525\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__36545\,
            I => \N__36520\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__36542\,
            I => \N__36520\
        );

    \I__8900\ : CascadeMux
    port map (
            O => \N__36541\,
            I => \N__36517\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__36536\,
            I => \N__36514\
        );

    \I__8898\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36510\
        );

    \I__8897\ : CascadeMux
    port map (
            O => \N__36534\,
            I => \N__36506\
        );

    \I__8896\ : InMux
    port map (
            O => \N__36533\,
            I => \N__36503\
        );

    \I__8895\ : InMux
    port map (
            O => \N__36532\,
            I => \N__36500\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__36529\,
            I => \N__36497\
        );

    \I__8893\ : InMux
    port map (
            O => \N__36528\,
            I => \N__36494\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__36525\,
            I => \N__36489\
        );

    \I__8891\ : Span4Mux_h
    port map (
            O => \N__36520\,
            I => \N__36489\
        );

    \I__8890\ : InMux
    port map (
            O => \N__36517\,
            I => \N__36486\
        );

    \I__8889\ : Span4Mux_h
    port map (
            O => \N__36514\,
            I => \N__36483\
        );

    \I__8888\ : InMux
    port map (
            O => \N__36513\,
            I => \N__36480\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__36510\,
            I => \N__36476\
        );

    \I__8886\ : InMux
    port map (
            O => \N__36509\,
            I => \N__36473\
        );

    \I__8885\ : InMux
    port map (
            O => \N__36506\,
            I => \N__36470\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__36503\,
            I => \N__36467\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__36500\,
            I => \N__36464\
        );

    \I__8882\ : Span4Mux_v
    port map (
            O => \N__36497\,
            I => \N__36461\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__36494\,
            I => \N__36458\
        );

    \I__8880\ : Span4Mux_s2_v
    port map (
            O => \N__36489\,
            I => \N__36446\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__36486\,
            I => \N__36446\
        );

    \I__8878\ : Span4Mux_s2_v
    port map (
            O => \N__36483\,
            I => \N__36446\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__36480\,
            I => \N__36443\
        );

    \I__8876\ : InMux
    port map (
            O => \N__36479\,
            I => \N__36440\
        );

    \I__8875\ : Span4Mux_v
    port map (
            O => \N__36476\,
            I => \N__36435\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__36473\,
            I => \N__36435\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__36470\,
            I => \N__36430\
        );

    \I__8872\ : Span4Mux_h
    port map (
            O => \N__36467\,
            I => \N__36430\
        );

    \I__8871\ : Span4Mux_v
    port map (
            O => \N__36464\,
            I => \N__36425\
        );

    \I__8870\ : Span4Mux_h
    port map (
            O => \N__36461\,
            I => \N__36425\
        );

    \I__8869\ : Span4Mux_h
    port map (
            O => \N__36458\,
            I => \N__36422\
        );

    \I__8868\ : InMux
    port map (
            O => \N__36457\,
            I => \N__36413\
        );

    \I__8867\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36413\
        );

    \I__8866\ : InMux
    port map (
            O => \N__36455\,
            I => \N__36413\
        );

    \I__8865\ : InMux
    port map (
            O => \N__36454\,
            I => \N__36413\
        );

    \I__8864\ : InMux
    port map (
            O => \N__36453\,
            I => \N__36410\
        );

    \I__8863\ : Span4Mux_v
    port map (
            O => \N__36446\,
            I => \N__36407\
        );

    \I__8862\ : Odrv4
    port map (
            O => \N__36443\,
            I => \tok.A_low_3\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__36440\,
            I => \tok.A_low_3\
        );

    \I__8860\ : Odrv4
    port map (
            O => \N__36435\,
            I => \tok.A_low_3\
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__36430\,
            I => \tok.A_low_3\
        );

    \I__8858\ : Odrv4
    port map (
            O => \N__36425\,
            I => \tok.A_low_3\
        );

    \I__8857\ : Odrv4
    port map (
            O => \N__36422\,
            I => \tok.A_low_3\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__36413\,
            I => \tok.A_low_3\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__36410\,
            I => \tok.A_low_3\
        );

    \I__8854\ : Odrv4
    port map (
            O => \N__36407\,
            I => \tok.A_low_3\
        );

    \I__8853\ : InMux
    port map (
            O => \N__36388\,
            I => \N__36385\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__36385\,
            I => \N__36382\
        );

    \I__8851\ : Span4Mux_v
    port map (
            O => \N__36382\,
            I => \N__36379\
        );

    \I__8850\ : Odrv4
    port map (
            O => \N__36379\,
            I => \tok.n168\
        );

    \I__8849\ : CascadeMux
    port map (
            O => \N__36376\,
            I => \N__36371\
        );

    \I__8848\ : InMux
    port map (
            O => \N__36375\,
            I => \N__36368\
        );

    \I__8847\ : InMux
    port map (
            O => \N__36374\,
            I => \N__36365\
        );

    \I__8846\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36361\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__36368\,
            I => \N__36358\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__36365\,
            I => \N__36355\
        );

    \I__8843\ : InMux
    port map (
            O => \N__36364\,
            I => \N__36352\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__36361\,
            I => \N__36349\
        );

    \I__8841\ : Span4Mux_h
    port map (
            O => \N__36358\,
            I => \N__36342\
        );

    \I__8840\ : Span4Mux_v
    port map (
            O => \N__36355\,
            I => \N__36342\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__36352\,
            I => \N__36342\
        );

    \I__8838\ : Span4Mux_h
    port map (
            O => \N__36349\,
            I => \N__36338\
        );

    \I__8837\ : Span4Mux_h
    port map (
            O => \N__36342\,
            I => \N__36335\
        );

    \I__8836\ : InMux
    port map (
            O => \N__36341\,
            I => \N__36332\
        );

    \I__8835\ : Odrv4
    port map (
            O => \N__36338\,
            I => \tok.n5_adj_682\
        );

    \I__8834\ : Odrv4
    port map (
            O => \N__36335\,
            I => \tok.n5_adj_682\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__36332\,
            I => \tok.n5_adj_682\
        );

    \I__8832\ : CascadeMux
    port map (
            O => \N__36325\,
            I => \N__36312\
        );

    \I__8831\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36307\
        );

    \I__8830\ : CascadeMux
    port map (
            O => \N__36323\,
            I => \N__36288\
        );

    \I__8829\ : CascadeMux
    port map (
            O => \N__36322\,
            I => \N__36276\
        );

    \I__8828\ : CascadeMux
    port map (
            O => \N__36321\,
            I => \N__36273\
        );

    \I__8827\ : CascadeMux
    port map (
            O => \N__36320\,
            I => \N__36270\
        );

    \I__8826\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36262\
        );

    \I__8825\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36262\
        );

    \I__8824\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36262\
        );

    \I__8823\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36246\
        );

    \I__8822\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36239\
        );

    \I__8821\ : InMux
    port map (
            O => \N__36312\,
            I => \N__36239\
        );

    \I__8820\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36239\
        );

    \I__8819\ : CascadeMux
    port map (
            O => \N__36310\,
            I => \N__36236\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__36307\,
            I => \N__36224\
        );

    \I__8817\ : InMux
    port map (
            O => \N__36306\,
            I => \N__36221\
        );

    \I__8816\ : CascadeMux
    port map (
            O => \N__36305\,
            I => \N__36216\
        );

    \I__8815\ : CascadeMux
    port map (
            O => \N__36304\,
            I => \N__36210\
        );

    \I__8814\ : CascadeMux
    port map (
            O => \N__36303\,
            I => \N__36207\
        );

    \I__8813\ : InMux
    port map (
            O => \N__36302\,
            I => \N__36199\
        );

    \I__8812\ : InMux
    port map (
            O => \N__36301\,
            I => \N__36199\
        );

    \I__8811\ : InMux
    port map (
            O => \N__36300\,
            I => \N__36199\
        );

    \I__8810\ : InMux
    port map (
            O => \N__36299\,
            I => \N__36196\
        );

    \I__8809\ : InMux
    port map (
            O => \N__36298\,
            I => \N__36191\
        );

    \I__8808\ : InMux
    port map (
            O => \N__36297\,
            I => \N__36191\
        );

    \I__8807\ : InMux
    port map (
            O => \N__36296\,
            I => \N__36186\
        );

    \I__8806\ : InMux
    port map (
            O => \N__36295\,
            I => \N__36186\
        );

    \I__8805\ : CascadeMux
    port map (
            O => \N__36294\,
            I => \N__36180\
        );

    \I__8804\ : InMux
    port map (
            O => \N__36293\,
            I => \N__36174\
        );

    \I__8803\ : InMux
    port map (
            O => \N__36292\,
            I => \N__36169\
        );

    \I__8802\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36169\
        );

    \I__8801\ : InMux
    port map (
            O => \N__36288\,
            I => \N__36166\
        );

    \I__8800\ : InMux
    port map (
            O => \N__36287\,
            I => \N__36157\
        );

    \I__8799\ : InMux
    port map (
            O => \N__36286\,
            I => \N__36157\
        );

    \I__8798\ : InMux
    port map (
            O => \N__36285\,
            I => \N__36157\
        );

    \I__8797\ : InMux
    port map (
            O => \N__36284\,
            I => \N__36157\
        );

    \I__8796\ : CascadeMux
    port map (
            O => \N__36283\,
            I => \N__36139\
        );

    \I__8795\ : InMux
    port map (
            O => \N__36282\,
            I => \N__36135\
        );

    \I__8794\ : InMux
    port map (
            O => \N__36281\,
            I => \N__36132\
        );

    \I__8793\ : InMux
    port map (
            O => \N__36280\,
            I => \N__36121\
        );

    \I__8792\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36121\
        );

    \I__8791\ : InMux
    port map (
            O => \N__36276\,
            I => \N__36121\
        );

    \I__8790\ : InMux
    port map (
            O => \N__36273\,
            I => \N__36121\
        );

    \I__8789\ : InMux
    port map (
            O => \N__36270\,
            I => \N__36121\
        );

    \I__8788\ : InMux
    port map (
            O => \N__36269\,
            I => \N__36118\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__36262\,
            I => \N__36115\
        );

    \I__8786\ : InMux
    port map (
            O => \N__36261\,
            I => \N__36108\
        );

    \I__8785\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36108\
        );

    \I__8784\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36108\
        );

    \I__8783\ : InMux
    port map (
            O => \N__36258\,
            I => \N__36103\
        );

    \I__8782\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36103\
        );

    \I__8781\ : CascadeMux
    port map (
            O => \N__36256\,
            I => \N__36099\
        );

    \I__8780\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36092\
        );

    \I__8779\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36092\
        );

    \I__8778\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36089\
        );

    \I__8777\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36086\
        );

    \I__8776\ : InMux
    port map (
            O => \N__36251\,
            I => \N__36079\
        );

    \I__8775\ : InMux
    port map (
            O => \N__36250\,
            I => \N__36079\
        );

    \I__8774\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36079\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__36246\,
            I => \N__36074\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__36239\,
            I => \N__36074\
        );

    \I__8771\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36065\
        );

    \I__8770\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36065\
        );

    \I__8769\ : InMux
    port map (
            O => \N__36234\,
            I => \N__36065\
        );

    \I__8768\ : InMux
    port map (
            O => \N__36233\,
            I => \N__36065\
        );

    \I__8767\ : InMux
    port map (
            O => \N__36232\,
            I => \N__36062\
        );

    \I__8766\ : CascadeMux
    port map (
            O => \N__36231\,
            I => \N__36059\
        );

    \I__8765\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36056\
        );

    \I__8764\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36053\
        );

    \I__8763\ : CascadeMux
    port map (
            O => \N__36228\,
            I => \N__36045\
        );

    \I__8762\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36041\
        );

    \I__8761\ : Span4Mux_h
    port map (
            O => \N__36224\,
            I => \N__36036\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__36221\,
            I => \N__36036\
        );

    \I__8759\ : InMux
    port map (
            O => \N__36220\,
            I => \N__36033\
        );

    \I__8758\ : InMux
    port map (
            O => \N__36219\,
            I => \N__36024\
        );

    \I__8757\ : InMux
    port map (
            O => \N__36216\,
            I => \N__36024\
        );

    \I__8756\ : InMux
    port map (
            O => \N__36215\,
            I => \N__36019\
        );

    \I__8755\ : InMux
    port map (
            O => \N__36214\,
            I => \N__36019\
        );

    \I__8754\ : CascadeMux
    port map (
            O => \N__36213\,
            I => \N__36011\
        );

    \I__8753\ : InMux
    port map (
            O => \N__36210\,
            I => \N__36002\
        );

    \I__8752\ : InMux
    port map (
            O => \N__36207\,
            I => \N__36002\
        );

    \I__8751\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36002\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__36199\,
            I => \N__35999\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__36196\,
            I => \N__35992\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__36191\,
            I => \N__35992\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__36186\,
            I => \N__35992\
        );

    \I__8746\ : InMux
    port map (
            O => \N__36185\,
            I => \N__35989\
        );

    \I__8745\ : InMux
    port map (
            O => \N__36184\,
            I => \N__35986\
        );

    \I__8744\ : InMux
    port map (
            O => \N__36183\,
            I => \N__35983\
        );

    \I__8743\ : InMux
    port map (
            O => \N__36180\,
            I => \N__35976\
        );

    \I__8742\ : InMux
    port map (
            O => \N__36179\,
            I => \N__35976\
        );

    \I__8741\ : InMux
    port map (
            O => \N__36178\,
            I => \N__35976\
        );

    \I__8740\ : InMux
    port map (
            O => \N__36177\,
            I => \N__35973\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__36174\,
            I => \N__35969\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__36169\,
            I => \N__35962\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__36166\,
            I => \N__35962\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__36157\,
            I => \N__35962\
        );

    \I__8735\ : InMux
    port map (
            O => \N__36156\,
            I => \N__35953\
        );

    \I__8734\ : InMux
    port map (
            O => \N__36155\,
            I => \N__35953\
        );

    \I__8733\ : InMux
    port map (
            O => \N__36154\,
            I => \N__35953\
        );

    \I__8732\ : InMux
    port map (
            O => \N__36153\,
            I => \N__35953\
        );

    \I__8731\ : InMux
    port map (
            O => \N__36152\,
            I => \N__35944\
        );

    \I__8730\ : InMux
    port map (
            O => \N__36151\,
            I => \N__35944\
        );

    \I__8729\ : InMux
    port map (
            O => \N__36150\,
            I => \N__35944\
        );

    \I__8728\ : InMux
    port map (
            O => \N__36149\,
            I => \N__35939\
        );

    \I__8727\ : InMux
    port map (
            O => \N__36148\,
            I => \N__35939\
        );

    \I__8726\ : InMux
    port map (
            O => \N__36147\,
            I => \N__35936\
        );

    \I__8725\ : InMux
    port map (
            O => \N__36146\,
            I => \N__35927\
        );

    \I__8724\ : InMux
    port map (
            O => \N__36145\,
            I => \N__35927\
        );

    \I__8723\ : InMux
    port map (
            O => \N__36144\,
            I => \N__35927\
        );

    \I__8722\ : InMux
    port map (
            O => \N__36143\,
            I => \N__35927\
        );

    \I__8721\ : InMux
    port map (
            O => \N__36142\,
            I => \N__35922\
        );

    \I__8720\ : InMux
    port map (
            O => \N__36139\,
            I => \N__35922\
        );

    \I__8719\ : CascadeMux
    port map (
            O => \N__36138\,
            I => \N__35919\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__36135\,
            I => \N__35915\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__36132\,
            I => \N__35910\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__36121\,
            I => \N__35910\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__36118\,
            I => \N__35901\
        );

    \I__8714\ : Span4Mux_v
    port map (
            O => \N__36115\,
            I => \N__35901\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__36108\,
            I => \N__35901\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__36103\,
            I => \N__35901\
        );

    \I__8711\ : InMux
    port map (
            O => \N__36102\,
            I => \N__35896\
        );

    \I__8710\ : InMux
    port map (
            O => \N__36099\,
            I => \N__35896\
        );

    \I__8709\ : InMux
    port map (
            O => \N__36098\,
            I => \N__35891\
        );

    \I__8708\ : InMux
    port map (
            O => \N__36097\,
            I => \N__35891\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__36092\,
            I => \N__35882\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__36089\,
            I => \N__35882\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__36086\,
            I => \N__35882\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__36079\,
            I => \N__35882\
        );

    \I__8703\ : Span4Mux_s2_v
    port map (
            O => \N__36074\,
            I => \N__35875\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__36065\,
            I => \N__35875\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__36062\,
            I => \N__35875\
        );

    \I__8700\ : InMux
    port map (
            O => \N__36059\,
            I => \N__35871\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__36056\,
            I => \N__35868\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__36053\,
            I => \N__35865\
        );

    \I__8697\ : InMux
    port map (
            O => \N__36052\,
            I => \N__35858\
        );

    \I__8696\ : InMux
    port map (
            O => \N__36051\,
            I => \N__35858\
        );

    \I__8695\ : InMux
    port map (
            O => \N__36050\,
            I => \N__35858\
        );

    \I__8694\ : InMux
    port map (
            O => \N__36049\,
            I => \N__35855\
        );

    \I__8693\ : InMux
    port map (
            O => \N__36048\,
            I => \N__35852\
        );

    \I__8692\ : InMux
    port map (
            O => \N__36045\,
            I => \N__35849\
        );

    \I__8691\ : InMux
    port map (
            O => \N__36044\,
            I => \N__35846\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__36041\,
            I => \N__35839\
        );

    \I__8689\ : Span4Mux_h
    port map (
            O => \N__36036\,
            I => \N__35839\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__36033\,
            I => \N__35839\
        );

    \I__8687\ : InMux
    port map (
            O => \N__36032\,
            I => \N__35836\
        );

    \I__8686\ : CascadeMux
    port map (
            O => \N__36031\,
            I => \N__35832\
        );

    \I__8685\ : InMux
    port map (
            O => \N__36030\,
            I => \N__35825\
        );

    \I__8684\ : InMux
    port map (
            O => \N__36029\,
            I => \N__35822\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__36024\,
            I => \N__35817\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__36019\,
            I => \N__35817\
        );

    \I__8681\ : InMux
    port map (
            O => \N__36018\,
            I => \N__35804\
        );

    \I__8680\ : InMux
    port map (
            O => \N__36017\,
            I => \N__35804\
        );

    \I__8679\ : InMux
    port map (
            O => \N__36016\,
            I => \N__35804\
        );

    \I__8678\ : InMux
    port map (
            O => \N__36015\,
            I => \N__35804\
        );

    \I__8677\ : InMux
    port map (
            O => \N__36014\,
            I => \N__35804\
        );

    \I__8676\ : InMux
    port map (
            O => \N__36011\,
            I => \N__35804\
        );

    \I__8675\ : InMux
    port map (
            O => \N__36010\,
            I => \N__35799\
        );

    \I__8674\ : InMux
    port map (
            O => \N__36009\,
            I => \N__35799\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__36002\,
            I => \N__35792\
        );

    \I__8672\ : Span4Mux_s3_h
    port map (
            O => \N__35999\,
            I => \N__35792\
        );

    \I__8671\ : Span4Mux_v
    port map (
            O => \N__35992\,
            I => \N__35792\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__35989\,
            I => \N__35783\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__35986\,
            I => \N__35783\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__35983\,
            I => \N__35783\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__35976\,
            I => \N__35783\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__35973\,
            I => \N__35780\
        );

    \I__8665\ : InMux
    port map (
            O => \N__35972\,
            I => \N__35775\
        );

    \I__8664\ : Span4Mux_v
    port map (
            O => \N__35969\,
            I => \N__35768\
        );

    \I__8663\ : Span4Mux_v
    port map (
            O => \N__35962\,
            I => \N__35768\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__35953\,
            I => \N__35768\
        );

    \I__8661\ : InMux
    port map (
            O => \N__35952\,
            I => \N__35758\
        );

    \I__8660\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35758\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__35944\,
            I => \N__35749\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__35939\,
            I => \N__35749\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__35936\,
            I => \N__35749\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__35927\,
            I => \N__35749\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__35922\,
            I => \N__35746\
        );

    \I__8654\ : InMux
    port map (
            O => \N__35919\,
            I => \N__35741\
        );

    \I__8653\ : InMux
    port map (
            O => \N__35918\,
            I => \N__35741\
        );

    \I__8652\ : Span4Mux_s3_v
    port map (
            O => \N__35915\,
            I => \N__35734\
        );

    \I__8651\ : Span4Mux_s3_v
    port map (
            O => \N__35910\,
            I => \N__35734\
        );

    \I__8650\ : Span4Mux_v
    port map (
            O => \N__35901\,
            I => \N__35734\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__35896\,
            I => \N__35725\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__35891\,
            I => \N__35725\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__35882\,
            I => \N__35725\
        );

    \I__8646\ : Span4Mux_v
    port map (
            O => \N__35875\,
            I => \N__35725\
        );

    \I__8645\ : CascadeMux
    port map (
            O => \N__35874\,
            I => \N__35718\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__35871\,
            I => \N__35712\
        );

    \I__8643\ : Span4Mux_v
    port map (
            O => \N__35868\,
            I => \N__35707\
        );

    \I__8642\ : Span4Mux_s3_v
    port map (
            O => \N__35865\,
            I => \N__35707\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__35858\,
            I => \N__35704\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__35855\,
            I => \N__35701\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__35852\,
            I => \N__35692\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__35849\,
            I => \N__35692\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__35846\,
            I => \N__35692\
        );

    \I__8636\ : Span4Mux_v
    port map (
            O => \N__35839\,
            I => \N__35692\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__35836\,
            I => \N__35689\
        );

    \I__8634\ : InMux
    port map (
            O => \N__35835\,
            I => \N__35676\
        );

    \I__8633\ : InMux
    port map (
            O => \N__35832\,
            I => \N__35676\
        );

    \I__8632\ : InMux
    port map (
            O => \N__35831\,
            I => \N__35676\
        );

    \I__8631\ : InMux
    port map (
            O => \N__35830\,
            I => \N__35676\
        );

    \I__8630\ : InMux
    port map (
            O => \N__35829\,
            I => \N__35676\
        );

    \I__8629\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35676\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__35825\,
            I => \N__35671\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__35822\,
            I => \N__35671\
        );

    \I__8626\ : Span4Mux_h
    port map (
            O => \N__35817\,
            I => \N__35668\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__35804\,
            I => \N__35659\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__35799\,
            I => \N__35659\
        );

    \I__8623\ : Span4Mux_h
    port map (
            O => \N__35792\,
            I => \N__35659\
        );

    \I__8622\ : Span4Mux_v
    port map (
            O => \N__35783\,
            I => \N__35659\
        );

    \I__8621\ : Span4Mux_s3_v
    port map (
            O => \N__35780\,
            I => \N__35656\
        );

    \I__8620\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35653\
        );

    \I__8619\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35650\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__35775\,
            I => \N__35647\
        );

    \I__8617\ : Span4Mux_s3_v
    port map (
            O => \N__35768\,
            I => \N__35644\
        );

    \I__8616\ : InMux
    port map (
            O => \N__35767\,
            I => \N__35641\
        );

    \I__8615\ : InMux
    port map (
            O => \N__35766\,
            I => \N__35632\
        );

    \I__8614\ : InMux
    port map (
            O => \N__35765\,
            I => \N__35632\
        );

    \I__8613\ : InMux
    port map (
            O => \N__35764\,
            I => \N__35632\
        );

    \I__8612\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35632\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35629\
        );

    \I__8610\ : Span4Mux_s3_v
    port map (
            O => \N__35749\,
            I => \N__35618\
        );

    \I__8609\ : Span4Mux_s3_v
    port map (
            O => \N__35746\,
            I => \N__35618\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__35741\,
            I => \N__35618\
        );

    \I__8607\ : Span4Mux_h
    port map (
            O => \N__35734\,
            I => \N__35618\
        );

    \I__8606\ : Span4Mux_v
    port map (
            O => \N__35725\,
            I => \N__35618\
        );

    \I__8605\ : InMux
    port map (
            O => \N__35724\,
            I => \N__35613\
        );

    \I__8604\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35613\
        );

    \I__8603\ : InMux
    port map (
            O => \N__35722\,
            I => \N__35607\
        );

    \I__8602\ : InMux
    port map (
            O => \N__35721\,
            I => \N__35598\
        );

    \I__8601\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35598\
        );

    \I__8600\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35598\
        );

    \I__8599\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35598\
        );

    \I__8598\ : InMux
    port map (
            O => \N__35715\,
            I => \N__35595\
        );

    \I__8597\ : Span12Mux_s10_v
    port map (
            O => \N__35712\,
            I => \N__35592\
        );

    \I__8596\ : Span4Mux_h
    port map (
            O => \N__35707\,
            I => \N__35573\
        );

    \I__8595\ : Span4Mux_s3_v
    port map (
            O => \N__35704\,
            I => \N__35573\
        );

    \I__8594\ : Span4Mux_v
    port map (
            O => \N__35701\,
            I => \N__35573\
        );

    \I__8593\ : Span4Mux_v
    port map (
            O => \N__35692\,
            I => \N__35573\
        );

    \I__8592\ : Span4Mux_s3_v
    port map (
            O => \N__35689\,
            I => \N__35573\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__35676\,
            I => \N__35573\
        );

    \I__8590\ : Span4Mux_s3_v
    port map (
            O => \N__35671\,
            I => \N__35573\
        );

    \I__8589\ : Span4Mux_v
    port map (
            O => \N__35668\,
            I => \N__35573\
        );

    \I__8588\ : Span4Mux_v
    port map (
            O => \N__35659\,
            I => \N__35573\
        );

    \I__8587\ : Sp12to4
    port map (
            O => \N__35656\,
            I => \N__35552\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__35653\,
            I => \N__35552\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__35650\,
            I => \N__35552\
        );

    \I__8584\ : Span12Mux_s10_v
    port map (
            O => \N__35647\,
            I => \N__35552\
        );

    \I__8583\ : Sp12to4
    port map (
            O => \N__35644\,
            I => \N__35552\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__35641\,
            I => \N__35552\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__35632\,
            I => \N__35552\
        );

    \I__8580\ : Span12Mux_s1_h
    port map (
            O => \N__35629\,
            I => \N__35552\
        );

    \I__8579\ : Sp12to4
    port map (
            O => \N__35618\,
            I => \N__35552\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__35613\,
            I => \N__35552\
        );

    \I__8577\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35549\
        );

    \I__8576\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35544\
        );

    \I__8575\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35544\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__35607\,
            I => \tok.T_4\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__35598\,
            I => \tok.T_4\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__35595\,
            I => \tok.T_4\
        );

    \I__8571\ : Odrv12
    port map (
            O => \N__35592\,
            I => \tok.T_4\
        );

    \I__8570\ : Odrv4
    port map (
            O => \N__35573\,
            I => \tok.T_4\
        );

    \I__8569\ : Odrv12
    port map (
            O => \N__35552\,
            I => \tok.T_4\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__35549\,
            I => \tok.T_4\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__35544\,
            I => \tok.T_4\
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__35527\,
            I => \tok.n6478_cascade_\
        );

    \I__8565\ : CascadeMux
    port map (
            O => \N__35524\,
            I => \N__35511\
        );

    \I__8564\ : CascadeMux
    port map (
            O => \N__35523\,
            I => \N__35497\
        );

    \I__8563\ : InMux
    port map (
            O => \N__35522\,
            I => \N__35475\
        );

    \I__8562\ : InMux
    port map (
            O => \N__35521\,
            I => \N__35469\
        );

    \I__8561\ : InMux
    port map (
            O => \N__35520\,
            I => \N__35469\
        );

    \I__8560\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35460\
        );

    \I__8559\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35460\
        );

    \I__8558\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35452\
        );

    \I__8557\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35447\
        );

    \I__8556\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35447\
        );

    \I__8555\ : InMux
    port map (
            O => \N__35514\,
            I => \N__35435\
        );

    \I__8554\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35435\
        );

    \I__8553\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35435\
        );

    \I__8552\ : InMux
    port map (
            O => \N__35509\,
            I => \N__35432\
        );

    \I__8551\ : InMux
    port map (
            O => \N__35508\,
            I => \N__35427\
        );

    \I__8550\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35427\
        );

    \I__8549\ : InMux
    port map (
            O => \N__35506\,
            I => \N__35424\
        );

    \I__8548\ : CascadeMux
    port map (
            O => \N__35505\,
            I => \N__35420\
        );

    \I__8547\ : InMux
    port map (
            O => \N__35504\,
            I => \N__35416\
        );

    \I__8546\ : CascadeMux
    port map (
            O => \N__35503\,
            I => \N__35412\
        );

    \I__8545\ : InMux
    port map (
            O => \N__35502\,
            I => \N__35409\
        );

    \I__8544\ : InMux
    port map (
            O => \N__35501\,
            I => \N__35406\
        );

    \I__8543\ : InMux
    port map (
            O => \N__35500\,
            I => \N__35403\
        );

    \I__8542\ : InMux
    port map (
            O => \N__35497\,
            I => \N__35398\
        );

    \I__8541\ : InMux
    port map (
            O => \N__35496\,
            I => \N__35398\
        );

    \I__8540\ : CascadeMux
    port map (
            O => \N__35495\,
            I => \N__35391\
        );

    \I__8539\ : InMux
    port map (
            O => \N__35494\,
            I => \N__35367\
        );

    \I__8538\ : InMux
    port map (
            O => \N__35493\,
            I => \N__35358\
        );

    \I__8537\ : InMux
    port map (
            O => \N__35492\,
            I => \N__35358\
        );

    \I__8536\ : InMux
    port map (
            O => \N__35491\,
            I => \N__35358\
        );

    \I__8535\ : InMux
    port map (
            O => \N__35490\,
            I => \N__35358\
        );

    \I__8534\ : InMux
    port map (
            O => \N__35489\,
            I => \N__35353\
        );

    \I__8533\ : InMux
    port map (
            O => \N__35488\,
            I => \N__35350\
        );

    \I__8532\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35347\
        );

    \I__8531\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35342\
        );

    \I__8530\ : InMux
    port map (
            O => \N__35485\,
            I => \N__35342\
        );

    \I__8529\ : InMux
    port map (
            O => \N__35484\,
            I => \N__35337\
        );

    \I__8528\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35337\
        );

    \I__8527\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35332\
        );

    \I__8526\ : InMux
    port map (
            O => \N__35481\,
            I => \N__35332\
        );

    \I__8525\ : InMux
    port map (
            O => \N__35480\,
            I => \N__35326\
        );

    \I__8524\ : InMux
    port map (
            O => \N__35479\,
            I => \N__35321\
        );

    \I__8523\ : InMux
    port map (
            O => \N__35478\,
            I => \N__35321\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__35475\,
            I => \N__35318\
        );

    \I__8521\ : InMux
    port map (
            O => \N__35474\,
            I => \N__35315\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__35469\,
            I => \N__35312\
        );

    \I__8519\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35305\
        );

    \I__8518\ : InMux
    port map (
            O => \N__35467\,
            I => \N__35305\
        );

    \I__8517\ : InMux
    port map (
            O => \N__35466\,
            I => \N__35305\
        );

    \I__8516\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35302\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__35460\,
            I => \N__35297\
        );

    \I__8514\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35288\
        );

    \I__8513\ : InMux
    port map (
            O => \N__35458\,
            I => \N__35288\
        );

    \I__8512\ : InMux
    port map (
            O => \N__35457\,
            I => \N__35288\
        );

    \I__8511\ : InMux
    port map (
            O => \N__35456\,
            I => \N__35288\
        );

    \I__8510\ : InMux
    port map (
            O => \N__35455\,
            I => \N__35285\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__35452\,
            I => \N__35280\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__35447\,
            I => \N__35280\
        );

    \I__8507\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35273\
        );

    \I__8506\ : InMux
    port map (
            O => \N__35445\,
            I => \N__35273\
        );

    \I__8505\ : CascadeMux
    port map (
            O => \N__35444\,
            I => \N__35269\
        );

    \I__8504\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35261\
        );

    \I__8503\ : InMux
    port map (
            O => \N__35442\,
            I => \N__35257\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__35435\,
            I => \N__35254\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__35432\,
            I => \N__35247\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__35427\,
            I => \N__35247\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__35424\,
            I => \N__35247\
        );

    \I__8498\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35242\
        );

    \I__8497\ : InMux
    port map (
            O => \N__35420\,
            I => \N__35242\
        );

    \I__8496\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35239\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__35416\,
            I => \N__35234\
        );

    \I__8494\ : InMux
    port map (
            O => \N__35415\,
            I => \N__35229\
        );

    \I__8493\ : InMux
    port map (
            O => \N__35412\,
            I => \N__35229\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__35409\,
            I => \N__35222\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__35406\,
            I => \N__35222\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__35403\,
            I => \N__35222\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__35398\,
            I => \N__35219\
        );

    \I__8488\ : InMux
    port map (
            O => \N__35397\,
            I => \N__35214\
        );

    \I__8487\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35214\
        );

    \I__8486\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35207\
        );

    \I__8485\ : InMux
    port map (
            O => \N__35394\,
            I => \N__35207\
        );

    \I__8484\ : InMux
    port map (
            O => \N__35391\,
            I => \N__35207\
        );

    \I__8483\ : InMux
    port map (
            O => \N__35390\,
            I => \N__35203\
        );

    \I__8482\ : InMux
    port map (
            O => \N__35389\,
            I => \N__35200\
        );

    \I__8481\ : InMux
    port map (
            O => \N__35388\,
            I => \N__35187\
        );

    \I__8480\ : InMux
    port map (
            O => \N__35387\,
            I => \N__35187\
        );

    \I__8479\ : InMux
    port map (
            O => \N__35386\,
            I => \N__35187\
        );

    \I__8478\ : InMux
    port map (
            O => \N__35385\,
            I => \N__35187\
        );

    \I__8477\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35187\
        );

    \I__8476\ : InMux
    port map (
            O => \N__35383\,
            I => \N__35180\
        );

    \I__8475\ : InMux
    port map (
            O => \N__35382\,
            I => \N__35180\
        );

    \I__8474\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35180\
        );

    \I__8473\ : InMux
    port map (
            O => \N__35380\,
            I => \N__35173\
        );

    \I__8472\ : InMux
    port map (
            O => \N__35379\,
            I => \N__35173\
        );

    \I__8471\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35173\
        );

    \I__8470\ : InMux
    port map (
            O => \N__35377\,
            I => \N__35170\
        );

    \I__8469\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35167\
        );

    \I__8468\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35164\
        );

    \I__8467\ : InMux
    port map (
            O => \N__35374\,
            I => \N__35159\
        );

    \I__8466\ : InMux
    port map (
            O => \N__35373\,
            I => \N__35159\
        );

    \I__8465\ : InMux
    port map (
            O => \N__35372\,
            I => \N__35152\
        );

    \I__8464\ : InMux
    port map (
            O => \N__35371\,
            I => \N__35152\
        );

    \I__8463\ : InMux
    port map (
            O => \N__35370\,
            I => \N__35152\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__35367\,
            I => \N__35147\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__35358\,
            I => \N__35147\
        );

    \I__8460\ : InMux
    port map (
            O => \N__35357\,
            I => \N__35142\
        );

    \I__8459\ : InMux
    port map (
            O => \N__35356\,
            I => \N__35142\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__35353\,
            I => \N__35137\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__35350\,
            I => \N__35137\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__35347\,
            I => \N__35128\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__35342\,
            I => \N__35128\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__35337\,
            I => \N__35128\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__35332\,
            I => \N__35128\
        );

    \I__8452\ : InMux
    port map (
            O => \N__35331\,
            I => \N__35124\
        );

    \I__8451\ : InMux
    port map (
            O => \N__35330\,
            I => \N__35121\
        );

    \I__8450\ : InMux
    port map (
            O => \N__35329\,
            I => \N__35118\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__35326\,
            I => \N__35115\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__35321\,
            I => \N__35110\
        );

    \I__8447\ : Span4Mux_s2_v
    port map (
            O => \N__35318\,
            I => \N__35110\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__35315\,
            I => \N__35103\
        );

    \I__8445\ : Span4Mux_v
    port map (
            O => \N__35312\,
            I => \N__35103\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__35305\,
            I => \N__35103\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__35302\,
            I => \N__35100\
        );

    \I__8442\ : InMux
    port map (
            O => \N__35301\,
            I => \N__35095\
        );

    \I__8441\ : InMux
    port map (
            O => \N__35300\,
            I => \N__35095\
        );

    \I__8440\ : Span4Mux_v
    port map (
            O => \N__35297\,
            I => \N__35090\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__35288\,
            I => \N__35090\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__35285\,
            I => \N__35085\
        );

    \I__8437\ : Span4Mux_v
    port map (
            O => \N__35280\,
            I => \N__35085\
        );

    \I__8436\ : InMux
    port map (
            O => \N__35279\,
            I => \N__35080\
        );

    \I__8435\ : InMux
    port map (
            O => \N__35278\,
            I => \N__35080\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__35273\,
            I => \N__35077\
        );

    \I__8433\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35070\
        );

    \I__8432\ : InMux
    port map (
            O => \N__35269\,
            I => \N__35070\
        );

    \I__8431\ : InMux
    port map (
            O => \N__35268\,
            I => \N__35070\
        );

    \I__8430\ : InMux
    port map (
            O => \N__35267\,
            I => \N__35067\
        );

    \I__8429\ : InMux
    port map (
            O => \N__35266\,
            I => \N__35064\
        );

    \I__8428\ : InMux
    port map (
            O => \N__35265\,
            I => \N__35061\
        );

    \I__8427\ : InMux
    port map (
            O => \N__35264\,
            I => \N__35058\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__35261\,
            I => \N__35054\
        );

    \I__8425\ : InMux
    port map (
            O => \N__35260\,
            I => \N__35051\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__35257\,
            I => \N__35044\
        );

    \I__8423\ : Span4Mux_s2_h
    port map (
            O => \N__35254\,
            I => \N__35044\
        );

    \I__8422\ : Span4Mux_v
    port map (
            O => \N__35247\,
            I => \N__35044\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__35242\,
            I => \N__35039\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__35239\,
            I => \N__35039\
        );

    \I__8419\ : InMux
    port map (
            O => \N__35238\,
            I => \N__35034\
        );

    \I__8418\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35034\
        );

    \I__8417\ : Span4Mux_h
    port map (
            O => \N__35234\,
            I => \N__35021\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__35229\,
            I => \N__35021\
        );

    \I__8415\ : Span4Mux_s3_v
    port map (
            O => \N__35222\,
            I => \N__35021\
        );

    \I__8414\ : Span4Mux_h
    port map (
            O => \N__35219\,
            I => \N__35021\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__35214\,
            I => \N__35021\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__35207\,
            I => \N__35021\
        );

    \I__8411\ : InMux
    port map (
            O => \N__35206\,
            I => \N__35018\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__35203\,
            I => \N__35015\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__35200\,
            I => \N__35012\
        );

    \I__8408\ : InMux
    port map (
            O => \N__35199\,
            I => \N__35009\
        );

    \I__8407\ : InMux
    port map (
            O => \N__35198\,
            I => \N__35006\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__35187\,
            I => \N__34999\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__35180\,
            I => \N__34999\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__35173\,
            I => \N__34999\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__35170\,
            I => \N__34986\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__35167\,
            I => \N__34986\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__35164\,
            I => \N__34986\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__35159\,
            I => \N__34986\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__35152\,
            I => \N__34986\
        );

    \I__8398\ : Span4Mux_v
    port map (
            O => \N__35147\,
            I => \N__34986\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__35142\,
            I => \N__34979\
        );

    \I__8396\ : Span4Mux_v
    port map (
            O => \N__35137\,
            I => \N__34979\
        );

    \I__8395\ : Span4Mux_v
    port map (
            O => \N__35128\,
            I => \N__34979\
        );

    \I__8394\ : InMux
    port map (
            O => \N__35127\,
            I => \N__34976\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__35124\,
            I => \N__34971\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__35121\,
            I => \N__34971\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__35118\,
            I => \N__34968\
        );

    \I__8390\ : Span4Mux_v
    port map (
            O => \N__35115\,
            I => \N__34965\
        );

    \I__8389\ : Span4Mux_v
    port map (
            O => \N__35110\,
            I => \N__34960\
        );

    \I__8388\ : Span4Mux_h
    port map (
            O => \N__35103\,
            I => \N__34960\
        );

    \I__8387\ : Span4Mux_s3_v
    port map (
            O => \N__35100\,
            I => \N__34949\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__35095\,
            I => \N__34949\
        );

    \I__8385\ : Span4Mux_s3_v
    port map (
            O => \N__35090\,
            I => \N__34949\
        );

    \I__8384\ : Span4Mux_v
    port map (
            O => \N__35085\,
            I => \N__34949\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__35080\,
            I => \N__34949\
        );

    \I__8382\ : Span4Mux_v
    port map (
            O => \N__35077\,
            I => \N__34942\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__35070\,
            I => \N__34942\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__35067\,
            I => \N__34942\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__35064\,
            I => \N__34935\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__35061\,
            I => \N__34935\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__35058\,
            I => \N__34935\
        );

    \I__8376\ : CascadeMux
    port map (
            O => \N__35057\,
            I => \N__34932\
        );

    \I__8375\ : Span4Mux_h
    port map (
            O => \N__35054\,
            I => \N__34927\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__35051\,
            I => \N__34927\
        );

    \I__8373\ : Span4Mux_h
    port map (
            O => \N__35044\,
            I => \N__34918\
        );

    \I__8372\ : Span4Mux_v
    port map (
            O => \N__35039\,
            I => \N__34918\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__35034\,
            I => \N__34918\
        );

    \I__8370\ : Span4Mux_v
    port map (
            O => \N__35021\,
            I => \N__34918\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__35018\,
            I => \N__34910\
        );

    \I__8368\ : Span4Mux_s2_v
    port map (
            O => \N__35015\,
            I => \N__34910\
        );

    \I__8367\ : Span4Mux_s2_v
    port map (
            O => \N__35012\,
            I => \N__34910\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__35009\,
            I => \N__34907\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__35006\,
            I => \N__34896\
        );

    \I__8364\ : Span4Mux_s2_v
    port map (
            O => \N__34999\,
            I => \N__34896\
        );

    \I__8363\ : Span4Mux_v
    port map (
            O => \N__34986\,
            I => \N__34896\
        );

    \I__8362\ : Span4Mux_h
    port map (
            O => \N__34979\,
            I => \N__34896\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__34976\,
            I => \N__34896\
        );

    \I__8360\ : Span12Mux_s10_v
    port map (
            O => \N__34971\,
            I => \N__34893\
        );

    \I__8359\ : Span4Mux_s3_v
    port map (
            O => \N__34968\,
            I => \N__34880\
        );

    \I__8358\ : Span4Mux_v
    port map (
            O => \N__34965\,
            I => \N__34880\
        );

    \I__8357\ : Span4Mux_v
    port map (
            O => \N__34960\,
            I => \N__34880\
        );

    \I__8356\ : Span4Mux_h
    port map (
            O => \N__34949\,
            I => \N__34880\
        );

    \I__8355\ : Span4Mux_s3_v
    port map (
            O => \N__34942\,
            I => \N__34880\
        );

    \I__8354\ : Span4Mux_s3_v
    port map (
            O => \N__34935\,
            I => \N__34880\
        );

    \I__8353\ : InMux
    port map (
            O => \N__34932\,
            I => \N__34877\
        );

    \I__8352\ : Span4Mux_v
    port map (
            O => \N__34927\,
            I => \N__34872\
        );

    \I__8351\ : Span4Mux_h
    port map (
            O => \N__34918\,
            I => \N__34872\
        );

    \I__8350\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34869\
        );

    \I__8349\ : Span4Mux_h
    port map (
            O => \N__34910\,
            I => \N__34862\
        );

    \I__8348\ : Span4Mux_v
    port map (
            O => \N__34907\,
            I => \N__34862\
        );

    \I__8347\ : Span4Mux_h
    port map (
            O => \N__34896\,
            I => \N__34862\
        );

    \I__8346\ : Odrv12
    port map (
            O => \N__34893\,
            I => \tok.T_6\
        );

    \I__8345\ : Odrv4
    port map (
            O => \N__34880\,
            I => \tok.T_6\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__34877\,
            I => \tok.T_6\
        );

    \I__8343\ : Odrv4
    port map (
            O => \N__34872\,
            I => \tok.T_6\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__34869\,
            I => \tok.T_6\
        );

    \I__8341\ : Odrv4
    port map (
            O => \N__34862\,
            I => \tok.T_6\
        );

    \I__8340\ : CascadeMux
    port map (
            O => \N__34849\,
            I => \tok.n186_adj_812_cascade_\
        );

    \I__8339\ : InMux
    port map (
            O => \N__34846\,
            I => \N__34835\
        );

    \I__8338\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34832\
        );

    \I__8337\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34827\
        );

    \I__8336\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34827\
        );

    \I__8335\ : InMux
    port map (
            O => \N__34842\,
            I => \N__34822\
        );

    \I__8334\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34822\
        );

    \I__8333\ : CascadeMux
    port map (
            O => \N__34840\,
            I => \N__34804\
        );

    \I__8332\ : CascadeMux
    port map (
            O => \N__34839\,
            I => \N__34787\
        );

    \I__8331\ : CascadeMux
    port map (
            O => \N__34838\,
            I => \N__34782\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__34835\,
            I => \N__34773\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__34832\,
            I => \N__34773\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__34827\,
            I => \N__34768\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__34822\,
            I => \N__34768\
        );

    \I__8326\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34765\
        );

    \I__8325\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34755\
        );

    \I__8324\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34743\
        );

    \I__8323\ : InMux
    port map (
            O => \N__34818\,
            I => \N__34743\
        );

    \I__8322\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34743\
        );

    \I__8321\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34736\
        );

    \I__8320\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34736\
        );

    \I__8319\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34736\
        );

    \I__8318\ : CascadeMux
    port map (
            O => \N__34813\,
            I => \N__34733\
        );

    \I__8317\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34730\
        );

    \I__8316\ : InMux
    port map (
            O => \N__34811\,
            I => \N__34727\
        );

    \I__8315\ : InMux
    port map (
            O => \N__34810\,
            I => \N__34724\
        );

    \I__8314\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34717\
        );

    \I__8313\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34717\
        );

    \I__8312\ : InMux
    port map (
            O => \N__34807\,
            I => \N__34714\
        );

    \I__8311\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34707\
        );

    \I__8310\ : CascadeMux
    port map (
            O => \N__34803\,
            I => \N__34701\
        );

    \I__8309\ : InMux
    port map (
            O => \N__34802\,
            I => \N__34690\
        );

    \I__8308\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34690\
        );

    \I__8307\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34690\
        );

    \I__8306\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34683\
        );

    \I__8305\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34683\
        );

    \I__8304\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34683\
        );

    \I__8303\ : CascadeMux
    port map (
            O => \N__34796\,
            I => \N__34677\
        );

    \I__8302\ : InMux
    port map (
            O => \N__34795\,
            I => \N__34672\
        );

    \I__8301\ : InMux
    port map (
            O => \N__34794\,
            I => \N__34665\
        );

    \I__8300\ : InMux
    port map (
            O => \N__34793\,
            I => \N__34665\
        );

    \I__8299\ : InMux
    port map (
            O => \N__34792\,
            I => \N__34665\
        );

    \I__8298\ : CascadeMux
    port map (
            O => \N__34791\,
            I => \N__34662\
        );

    \I__8297\ : InMux
    port map (
            O => \N__34790\,
            I => \N__34657\
        );

    \I__8296\ : InMux
    port map (
            O => \N__34787\,
            I => \N__34654\
        );

    \I__8295\ : InMux
    port map (
            O => \N__34786\,
            I => \N__34649\
        );

    \I__8294\ : InMux
    port map (
            O => \N__34785\,
            I => \N__34649\
        );

    \I__8293\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34644\
        );

    \I__8292\ : InMux
    port map (
            O => \N__34781\,
            I => \N__34644\
        );

    \I__8291\ : CascadeMux
    port map (
            O => \N__34780\,
            I => \N__34640\
        );

    \I__8290\ : InMux
    port map (
            O => \N__34779\,
            I => \N__34637\
        );

    \I__8289\ : InMux
    port map (
            O => \N__34778\,
            I => \N__34634\
        );

    \I__8288\ : Span4Mux_v
    port map (
            O => \N__34773\,
            I => \N__34627\
        );

    \I__8287\ : Span4Mux_v
    port map (
            O => \N__34768\,
            I => \N__34627\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34627\
        );

    \I__8285\ : InMux
    port map (
            O => \N__34764\,
            I => \N__34624\
        );

    \I__8284\ : InMux
    port map (
            O => \N__34763\,
            I => \N__34615\
        );

    \I__8283\ : InMux
    port map (
            O => \N__34762\,
            I => \N__34615\
        );

    \I__8282\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34615\
        );

    \I__8281\ : InMux
    port map (
            O => \N__34760\,
            I => \N__34615\
        );

    \I__8280\ : CascadeMux
    port map (
            O => \N__34759\,
            I => \N__34607\
        );

    \I__8279\ : CascadeMux
    port map (
            O => \N__34758\,
            I => \N__34603\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__34755\,
            I => \N__34600\
        );

    \I__8277\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34595\
        );

    \I__8276\ : InMux
    port map (
            O => \N__34753\,
            I => \N__34595\
        );

    \I__8275\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34590\
        );

    \I__8274\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34590\
        );

    \I__8273\ : InMux
    port map (
            O => \N__34750\,
            I => \N__34587\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__34743\,
            I => \N__34582\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__34736\,
            I => \N__34582\
        );

    \I__8270\ : InMux
    port map (
            O => \N__34733\,
            I => \N__34579\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__34730\,
            I => \N__34574\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__34727\,
            I => \N__34574\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__34724\,
            I => \N__34571\
        );

    \I__8266\ : InMux
    port map (
            O => \N__34723\,
            I => \N__34566\
        );

    \I__8265\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34566\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__34717\,
            I => \N__34561\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__34714\,
            I => \N__34561\
        );

    \I__8262\ : CascadeMux
    port map (
            O => \N__34713\,
            I => \N__34555\
        );

    \I__8261\ : CascadeMux
    port map (
            O => \N__34712\,
            I => \N__34552\
        );

    \I__8260\ : CascadeMux
    port map (
            O => \N__34711\,
            I => \N__34548\
        );

    \I__8259\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34544\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__34707\,
            I => \N__34541\
        );

    \I__8257\ : CascadeMux
    port map (
            O => \N__34706\,
            I => \N__34538\
        );

    \I__8256\ : InMux
    port map (
            O => \N__34705\,
            I => \N__34532\
        );

    \I__8255\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34529\
        );

    \I__8254\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34524\
        );

    \I__8253\ : InMux
    port map (
            O => \N__34700\,
            I => \N__34518\
        );

    \I__8252\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34518\
        );

    \I__8251\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34515\
        );

    \I__8250\ : InMux
    port map (
            O => \N__34697\,
            I => \N__34511\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__34690\,
            I => \N__34506\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__34683\,
            I => \N__34506\
        );

    \I__8247\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34497\
        );

    \I__8246\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34497\
        );

    \I__8245\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34497\
        );

    \I__8244\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34497\
        );

    \I__8243\ : InMux
    port map (
            O => \N__34676\,
            I => \N__34492\
        );

    \I__8242\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34492\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__34672\,
            I => \N__34487\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__34665\,
            I => \N__34487\
        );

    \I__8239\ : InMux
    port map (
            O => \N__34662\,
            I => \N__34484\
        );

    \I__8238\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34476\
        );

    \I__8237\ : InMux
    port map (
            O => \N__34660\,
            I => \N__34476\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__34657\,
            I => \N__34467\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__34654\,
            I => \N__34467\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__34649\,
            I => \N__34467\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__34644\,
            I => \N__34467\
        );

    \I__8232\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34462\
        );

    \I__8231\ : InMux
    port map (
            O => \N__34640\,
            I => \N__34462\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__34637\,
            I => \N__34451\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__34634\,
            I => \N__34451\
        );

    \I__8228\ : Span4Mux_h
    port map (
            O => \N__34627\,
            I => \N__34451\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__34624\,
            I => \N__34451\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__34615\,
            I => \N__34448\
        );

    \I__8225\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34443\
        );

    \I__8224\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34443\
        );

    \I__8223\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34436\
        );

    \I__8222\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34436\
        );

    \I__8221\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34436\
        );

    \I__8220\ : InMux
    port map (
            O => \N__34607\,
            I => \N__34429\
        );

    \I__8219\ : InMux
    port map (
            O => \N__34606\,
            I => \N__34429\
        );

    \I__8218\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34429\
        );

    \I__8217\ : Span4Mux_h
    port map (
            O => \N__34600\,
            I => \N__34425\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__34595\,
            I => \N__34420\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__34590\,
            I => \N__34420\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__34587\,
            I => \N__34415\
        );

    \I__8213\ : Span4Mux_v
    port map (
            O => \N__34582\,
            I => \N__34415\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__34579\,
            I => \N__34404\
        );

    \I__8211\ : Span4Mux_v
    port map (
            O => \N__34574\,
            I => \N__34404\
        );

    \I__8210\ : Span4Mux_s2_h
    port map (
            O => \N__34571\,
            I => \N__34404\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__34566\,
            I => \N__34404\
        );

    \I__8208\ : Span4Mux_s2_h
    port map (
            O => \N__34561\,
            I => \N__34404\
        );

    \I__8207\ : CascadeMux
    port map (
            O => \N__34560\,
            I => \N__34401\
        );

    \I__8206\ : CascadeMux
    port map (
            O => \N__34559\,
            I => \N__34398\
        );

    \I__8205\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34394\
        );

    \I__8204\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34391\
        );

    \I__8203\ : InMux
    port map (
            O => \N__34552\,
            I => \N__34384\
        );

    \I__8202\ : InMux
    port map (
            O => \N__34551\,
            I => \N__34384\
        );

    \I__8201\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34384\
        );

    \I__8200\ : InMux
    port map (
            O => \N__34547\,
            I => \N__34381\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34376\
        );

    \I__8198\ : Span4Mux_s3_v
    port map (
            O => \N__34541\,
            I => \N__34376\
        );

    \I__8197\ : InMux
    port map (
            O => \N__34538\,
            I => \N__34371\
        );

    \I__8196\ : InMux
    port map (
            O => \N__34537\,
            I => \N__34371\
        );

    \I__8195\ : InMux
    port map (
            O => \N__34536\,
            I => \N__34368\
        );

    \I__8194\ : InMux
    port map (
            O => \N__34535\,
            I => \N__34365\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__34532\,
            I => \N__34360\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__34529\,
            I => \N__34360\
        );

    \I__8191\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34355\
        );

    \I__8190\ : InMux
    port map (
            O => \N__34527\,
            I => \N__34355\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__34524\,
            I => \N__34352\
        );

    \I__8188\ : InMux
    port map (
            O => \N__34523\,
            I => \N__34349\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__34518\,
            I => \N__34344\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__34515\,
            I => \N__34344\
        );

    \I__8185\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34341\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__34511\,
            I => \N__34334\
        );

    \I__8183\ : Span4Mux_v
    port map (
            O => \N__34506\,
            I => \N__34334\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__34497\,
            I => \N__34334\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__34492\,
            I => \N__34331\
        );

    \I__8180\ : Span4Mux_s1_v
    port map (
            O => \N__34487\,
            I => \N__34326\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__34484\,
            I => \N__34326\
        );

    \I__8178\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34321\
        );

    \I__8177\ : InMux
    port map (
            O => \N__34482\,
            I => \N__34321\
        );

    \I__8176\ : InMux
    port map (
            O => \N__34481\,
            I => \N__34318\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__34476\,
            I => \N__34311\
        );

    \I__8174\ : Span4Mux_h
    port map (
            O => \N__34467\,
            I => \N__34311\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__34462\,
            I => \N__34311\
        );

    \I__8172\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34308\
        );

    \I__8171\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34305\
        );

    \I__8170\ : Span4Mux_v
    port map (
            O => \N__34451\,
            I => \N__34300\
        );

    \I__8169\ : Span4Mux_v
    port map (
            O => \N__34448\,
            I => \N__34300\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__34443\,
            I => \N__34293\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__34436\,
            I => \N__34293\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__34429\,
            I => \N__34293\
        );

    \I__8165\ : CascadeMux
    port map (
            O => \N__34428\,
            I => \N__34290\
        );

    \I__8164\ : Span4Mux_v
    port map (
            O => \N__34425\,
            I => \N__34281\
        );

    \I__8163\ : Span4Mux_v
    port map (
            O => \N__34420\,
            I => \N__34281\
        );

    \I__8162\ : Span4Mux_h
    port map (
            O => \N__34415\,
            I => \N__34281\
        );

    \I__8161\ : Span4Mux_h
    port map (
            O => \N__34404\,
            I => \N__34281\
        );

    \I__8160\ : InMux
    port map (
            O => \N__34401\,
            I => \N__34276\
        );

    \I__8159\ : InMux
    port map (
            O => \N__34398\,
            I => \N__34276\
        );

    \I__8158\ : InMux
    port map (
            O => \N__34397\,
            I => \N__34261\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__34394\,
            I => \N__34258\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__34391\,
            I => \N__34253\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__34384\,
            I => \N__34253\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__34381\,
            I => \N__34246\
        );

    \I__8153\ : Span4Mux_v
    port map (
            O => \N__34376\,
            I => \N__34246\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__34371\,
            I => \N__34246\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__34368\,
            I => \N__34237\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__34365\,
            I => \N__34237\
        );

    \I__8149\ : Span4Mux_v
    port map (
            O => \N__34360\,
            I => \N__34237\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__34355\,
            I => \N__34237\
        );

    \I__8147\ : Span4Mux_v
    port map (
            O => \N__34352\,
            I => \N__34226\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__34349\,
            I => \N__34226\
        );

    \I__8145\ : Span4Mux_s3_h
    port map (
            O => \N__34344\,
            I => \N__34226\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__34341\,
            I => \N__34226\
        );

    \I__8143\ : Span4Mux_v
    port map (
            O => \N__34334\,
            I => \N__34226\
        );

    \I__8142\ : Span4Mux_h
    port map (
            O => \N__34331\,
            I => \N__34219\
        );

    \I__8141\ : Span4Mux_v
    port map (
            O => \N__34326\,
            I => \N__34219\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__34321\,
            I => \N__34219\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__34318\,
            I => \N__34212\
        );

    \I__8138\ : Span4Mux_h
    port map (
            O => \N__34311\,
            I => \N__34212\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__34308\,
            I => \N__34212\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__34305\,
            I => \N__34205\
        );

    \I__8135\ : Span4Mux_h
    port map (
            O => \N__34300\,
            I => \N__34205\
        );

    \I__8134\ : Span4Mux_v
    port map (
            O => \N__34293\,
            I => \N__34205\
        );

    \I__8133\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34202\
        );

    \I__8132\ : Span4Mux_h
    port map (
            O => \N__34281\,
            I => \N__34197\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__34276\,
            I => \N__34197\
        );

    \I__8130\ : InMux
    port map (
            O => \N__34275\,
            I => \N__34190\
        );

    \I__8129\ : InMux
    port map (
            O => \N__34274\,
            I => \N__34190\
        );

    \I__8128\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34190\
        );

    \I__8127\ : InMux
    port map (
            O => \N__34272\,
            I => \N__34185\
        );

    \I__8126\ : InMux
    port map (
            O => \N__34271\,
            I => \N__34185\
        );

    \I__8125\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34176\
        );

    \I__8124\ : InMux
    port map (
            O => \N__34269\,
            I => \N__34176\
        );

    \I__8123\ : InMux
    port map (
            O => \N__34268\,
            I => \N__34176\
        );

    \I__8122\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34176\
        );

    \I__8121\ : InMux
    port map (
            O => \N__34266\,
            I => \N__34169\
        );

    \I__8120\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34169\
        );

    \I__8119\ : InMux
    port map (
            O => \N__34264\,
            I => \N__34169\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__34261\,
            I => \N__34156\
        );

    \I__8117\ : Span4Mux_s2_v
    port map (
            O => \N__34258\,
            I => \N__34156\
        );

    \I__8116\ : Span4Mux_v
    port map (
            O => \N__34253\,
            I => \N__34156\
        );

    \I__8115\ : Span4Mux_v
    port map (
            O => \N__34246\,
            I => \N__34156\
        );

    \I__8114\ : Span4Mux_v
    port map (
            O => \N__34237\,
            I => \N__34156\
        );

    \I__8113\ : Span4Mux_h
    port map (
            O => \N__34226\,
            I => \N__34156\
        );

    \I__8112\ : Span4Mux_h
    port map (
            O => \N__34219\,
            I => \N__34149\
        );

    \I__8111\ : Span4Mux_v
    port map (
            O => \N__34212\,
            I => \N__34149\
        );

    \I__8110\ : Span4Mux_h
    port map (
            O => \N__34205\,
            I => \N__34149\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__34202\,
            I => \N__34144\
        );

    \I__8108\ : Span4Mux_v
    port map (
            O => \N__34197\,
            I => \N__34144\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__34190\,
            I => \tok.T_3\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__34185\,
            I => \tok.T_3\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__34176\,
            I => \tok.T_3\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__34169\,
            I => \tok.T_3\
        );

    \I__8103\ : Odrv4
    port map (
            O => \N__34156\,
            I => \tok.T_3\
        );

    \I__8102\ : Odrv4
    port map (
            O => \N__34149\,
            I => \tok.T_3\
        );

    \I__8101\ : Odrv4
    port map (
            O => \N__34144\,
            I => \tok.T_3\
        );

    \I__8100\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34126\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__34126\,
            I => \N__34123\
        );

    \I__8098\ : Span4Mux_h
    port map (
            O => \N__34123\,
            I => \N__34120\
        );

    \I__8097\ : Span4Mux_h
    port map (
            O => \N__34120\,
            I => \N__34117\
        );

    \I__8096\ : Odrv4
    port map (
            O => \N__34117\,
            I => \tok.n338_adj_819\
        );

    \I__8095\ : CascadeMux
    port map (
            O => \N__34114\,
            I => \N__34109\
        );

    \I__8094\ : CascadeMux
    port map (
            O => \N__34113\,
            I => \N__34097\
        );

    \I__8093\ : CascadeMux
    port map (
            O => \N__34112\,
            I => \N__34089\
        );

    \I__8092\ : InMux
    port map (
            O => \N__34109\,
            I => \N__34084\
        );

    \I__8091\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34084\
        );

    \I__8090\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34072\
        );

    \I__8089\ : InMux
    port map (
            O => \N__34106\,
            I => \N__34064\
        );

    \I__8088\ : InMux
    port map (
            O => \N__34105\,
            I => \N__34064\
        );

    \I__8087\ : CascadeMux
    port map (
            O => \N__34104\,
            I => \N__34056\
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__34103\,
            I => \N__34049\
        );

    \I__8085\ : CascadeMux
    port map (
            O => \N__34102\,
            I => \N__34042\
        );

    \I__8084\ : CascadeMux
    port map (
            O => \N__34101\,
            I => \N__34037\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__34100\,
            I => \N__34032\
        );

    \I__8082\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34027\
        );

    \I__8081\ : CascadeMux
    port map (
            O => \N__34096\,
            I => \N__34023\
        );

    \I__8080\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34020\
        );

    \I__8079\ : InMux
    port map (
            O => \N__34094\,
            I => \N__34017\
        );

    \I__8078\ : InMux
    port map (
            O => \N__34093\,
            I => \N__34012\
        );

    \I__8077\ : InMux
    port map (
            O => \N__34092\,
            I => \N__34012\
        );

    \I__8076\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34009\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__34084\,
            I => \N__34006\
        );

    \I__8074\ : InMux
    port map (
            O => \N__34083\,
            I => \N__33996\
        );

    \I__8073\ : InMux
    port map (
            O => \N__34082\,
            I => \N__33996\
        );

    \I__8072\ : InMux
    port map (
            O => \N__34081\,
            I => \N__33996\
        );

    \I__8071\ : CascadeMux
    port map (
            O => \N__34080\,
            I => \N__33991\
        );

    \I__8070\ : CascadeMux
    port map (
            O => \N__34079\,
            I => \N__33988\
        );

    \I__8069\ : InMux
    port map (
            O => \N__34078\,
            I => \N__33981\
        );

    \I__8068\ : InMux
    port map (
            O => \N__34077\,
            I => \N__33981\
        );

    \I__8067\ : InMux
    port map (
            O => \N__34076\,
            I => \N__33974\
        );

    \I__8066\ : InMux
    port map (
            O => \N__34075\,
            I => \N__33974\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__34072\,
            I => \N__33971\
        );

    \I__8064\ : InMux
    port map (
            O => \N__34071\,
            I => \N__33968\
        );

    \I__8063\ : InMux
    port map (
            O => \N__34070\,
            I => \N__33963\
        );

    \I__8062\ : InMux
    port map (
            O => \N__34069\,
            I => \N__33963\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__34064\,
            I => \N__33960\
        );

    \I__8060\ : InMux
    port map (
            O => \N__34063\,
            I => \N__33953\
        );

    \I__8059\ : InMux
    port map (
            O => \N__34062\,
            I => \N__33953\
        );

    \I__8058\ : InMux
    port map (
            O => \N__34061\,
            I => \N__33953\
        );

    \I__8057\ : CascadeMux
    port map (
            O => \N__34060\,
            I => \N__33947\
        );

    \I__8056\ : InMux
    port map (
            O => \N__34059\,
            I => \N__33942\
        );

    \I__8055\ : InMux
    port map (
            O => \N__34056\,
            I => \N__33937\
        );

    \I__8054\ : InMux
    port map (
            O => \N__34055\,
            I => \N__33937\
        );

    \I__8053\ : InMux
    port map (
            O => \N__34054\,
            I => \N__33931\
        );

    \I__8052\ : InMux
    port map (
            O => \N__34053\,
            I => \N__33926\
        );

    \I__8051\ : InMux
    port map (
            O => \N__34052\,
            I => \N__33926\
        );

    \I__8050\ : InMux
    port map (
            O => \N__34049\,
            I => \N__33923\
        );

    \I__8049\ : InMux
    port map (
            O => \N__34048\,
            I => \N__33916\
        );

    \I__8048\ : InMux
    port map (
            O => \N__34047\,
            I => \N__33916\
        );

    \I__8047\ : InMux
    port map (
            O => \N__34046\,
            I => \N__33916\
        );

    \I__8046\ : InMux
    port map (
            O => \N__34045\,
            I => \N__33909\
        );

    \I__8045\ : InMux
    port map (
            O => \N__34042\,
            I => \N__33909\
        );

    \I__8044\ : InMux
    port map (
            O => \N__34041\,
            I => \N__33909\
        );

    \I__8043\ : InMux
    port map (
            O => \N__34040\,
            I => \N__33906\
        );

    \I__8042\ : InMux
    port map (
            O => \N__34037\,
            I => \N__33899\
        );

    \I__8041\ : InMux
    port map (
            O => \N__34036\,
            I => \N__33899\
        );

    \I__8040\ : InMux
    port map (
            O => \N__34035\,
            I => \N__33899\
        );

    \I__8039\ : InMux
    port map (
            O => \N__34032\,
            I => \N__33892\
        );

    \I__8038\ : InMux
    port map (
            O => \N__34031\,
            I => \N__33892\
        );

    \I__8037\ : InMux
    port map (
            O => \N__34030\,
            I => \N__33892\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__34027\,
            I => \N__33889\
        );

    \I__8035\ : InMux
    port map (
            O => \N__34026\,
            I => \N__33884\
        );

    \I__8034\ : InMux
    port map (
            O => \N__34023\,
            I => \N__33884\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__34020\,
            I => \N__33873\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__34017\,
            I => \N__33873\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__34012\,
            I => \N__33873\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__34009\,
            I => \N__33873\
        );

    \I__8029\ : Span4Mux_v
    port map (
            O => \N__34006\,
            I => \N__33873\
        );

    \I__8028\ : InMux
    port map (
            O => \N__34005\,
            I => \N__33868\
        );

    \I__8027\ : InMux
    port map (
            O => \N__34004\,
            I => \N__33863\
        );

    \I__8026\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33863\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__33996\,
            I => \N__33860\
        );

    \I__8024\ : InMux
    port map (
            O => \N__33995\,
            I => \N__33857\
        );

    \I__8023\ : InMux
    port map (
            O => \N__33994\,
            I => \N__33848\
        );

    \I__8022\ : InMux
    port map (
            O => \N__33991\,
            I => \N__33848\
        );

    \I__8021\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33848\
        );

    \I__8020\ : InMux
    port map (
            O => \N__33987\,
            I => \N__33848\
        );

    \I__8019\ : InMux
    port map (
            O => \N__33986\,
            I => \N__33845\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__33981\,
            I => \N__33842\
        );

    \I__8017\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33837\
        );

    \I__8016\ : InMux
    port map (
            O => \N__33979\,
            I => \N__33837\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__33974\,
            I => \N__33834\
        );

    \I__8014\ : Span4Mux_v
    port map (
            O => \N__33971\,
            I => \N__33827\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__33968\,
            I => \N__33827\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__33963\,
            I => \N__33827\
        );

    \I__8011\ : Span4Mux_v
    port map (
            O => \N__33960\,
            I => \N__33822\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__33953\,
            I => \N__33822\
        );

    \I__8009\ : InMux
    port map (
            O => \N__33952\,
            I => \N__33813\
        );

    \I__8008\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33813\
        );

    \I__8007\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33813\
        );

    \I__8006\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33813\
        );

    \I__8005\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33808\
        );

    \I__8004\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33808\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__33942\,
            I => \N__33803\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__33937\,
            I => \N__33803\
        );

    \I__8001\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33799\
        );

    \I__8000\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33792\
        );

    \I__7999\ : InMux
    port map (
            O => \N__33934\,
            I => \N__33792\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__33931\,
            I => \N__33789\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__33926\,
            I => \N__33786\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__33923\,
            I => \N__33779\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__33916\,
            I => \N__33779\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__33909\,
            I => \N__33779\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__33906\,
            I => \N__33770\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33770\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__33892\,
            I => \N__33770\
        );

    \I__7990\ : Span4Mux_v
    port map (
            O => \N__33889\,
            I => \N__33770\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__33884\,
            I => \N__33765\
        );

    \I__7988\ : Span4Mux_v
    port map (
            O => \N__33873\,
            I => \N__33765\
        );

    \I__7987\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33760\
        );

    \I__7986\ : InMux
    port map (
            O => \N__33871\,
            I => \N__33760\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__33868\,
            I => \N__33757\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__33863\,
            I => \N__33754\
        );

    \I__7983\ : Span4Mux_v
    port map (
            O => \N__33860\,
            I => \N__33751\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__33857\,
            I => \N__33746\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__33848\,
            I => \N__33746\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__33845\,
            I => \N__33733\
        );

    \I__7979\ : Span4Mux_s3_h
    port map (
            O => \N__33842\,
            I => \N__33733\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__33837\,
            I => \N__33733\
        );

    \I__7977\ : Span4Mux_v
    port map (
            O => \N__33834\,
            I => \N__33733\
        );

    \I__7976\ : Span4Mux_s3_v
    port map (
            O => \N__33827\,
            I => \N__33733\
        );

    \I__7975\ : Span4Mux_v
    port map (
            O => \N__33822\,
            I => \N__33733\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__33813\,
            I => \N__33730\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__33808\,
            I => \N__33727\
        );

    \I__7972\ : Span4Mux_v
    port map (
            O => \N__33803\,
            I => \N__33724\
        );

    \I__7971\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33721\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__33799\,
            I => \N__33718\
        );

    \I__7969\ : InMux
    port map (
            O => \N__33798\,
            I => \N__33715\
        );

    \I__7968\ : CascadeMux
    port map (
            O => \N__33797\,
            I => \N__33712\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__33792\,
            I => \N__33696\
        );

    \I__7966\ : Span4Mux_s2_v
    port map (
            O => \N__33789\,
            I => \N__33696\
        );

    \I__7965\ : Span4Mux_h
    port map (
            O => \N__33786\,
            I => \N__33696\
        );

    \I__7964\ : Span4Mux_s2_v
    port map (
            O => \N__33779\,
            I => \N__33696\
        );

    \I__7963\ : Span4Mux_v
    port map (
            O => \N__33770\,
            I => \N__33696\
        );

    \I__7962\ : Span4Mux_h
    port map (
            O => \N__33765\,
            I => \N__33696\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__33760\,
            I => \N__33696\
        );

    \I__7960\ : Span4Mux_h
    port map (
            O => \N__33757\,
            I => \N__33693\
        );

    \I__7959\ : Span4Mux_s3_v
    port map (
            O => \N__33754\,
            I => \N__33682\
        );

    \I__7958\ : Span4Mux_v
    port map (
            O => \N__33751\,
            I => \N__33682\
        );

    \I__7957\ : Span4Mux_s3_v
    port map (
            O => \N__33746\,
            I => \N__33682\
        );

    \I__7956\ : Span4Mux_h
    port map (
            O => \N__33733\,
            I => \N__33682\
        );

    \I__7955\ : Span4Mux_s3_v
    port map (
            O => \N__33730\,
            I => \N__33682\
        );

    \I__7954\ : Span4Mux_h
    port map (
            O => \N__33727\,
            I => \N__33675\
        );

    \I__7953\ : Span4Mux_h
    port map (
            O => \N__33724\,
            I => \N__33675\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__33721\,
            I => \N__33675\
        );

    \I__7951\ : Span4Mux_s3_v
    port map (
            O => \N__33718\,
            I => \N__33670\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__33715\,
            I => \N__33670\
        );

    \I__7949\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33667\
        );

    \I__7948\ : InMux
    port map (
            O => \N__33711\,
            I => \N__33664\
        );

    \I__7947\ : Span4Mux_h
    port map (
            O => \N__33696\,
            I => \N__33661\
        );

    \I__7946\ : Odrv4
    port map (
            O => \N__33693\,
            I => \tok.T_7\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__33682\,
            I => \tok.T_7\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__33675\,
            I => \tok.T_7\
        );

    \I__7943\ : Odrv4
    port map (
            O => \N__33670\,
            I => \tok.T_7\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__33667\,
            I => \tok.T_7\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__33664\,
            I => \tok.T_7\
        );

    \I__7940\ : Odrv4
    port map (
            O => \N__33661\,
            I => \tok.T_7\
        );

    \I__7939\ : CascadeMux
    port map (
            O => \N__33646\,
            I => \N__33639\
        );

    \I__7938\ : CascadeMux
    port map (
            O => \N__33645\,
            I => \N__33636\
        );

    \I__7937\ : InMux
    port map (
            O => \N__33644\,
            I => \N__33629\
        );

    \I__7936\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33626\
        );

    \I__7935\ : InMux
    port map (
            O => \N__33642\,
            I => \N__33622\
        );

    \I__7934\ : InMux
    port map (
            O => \N__33639\,
            I => \N__33619\
        );

    \I__7933\ : InMux
    port map (
            O => \N__33636\,
            I => \N__33616\
        );

    \I__7932\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33611\
        );

    \I__7931\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33611\
        );

    \I__7930\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33604\
        );

    \I__7929\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33601\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__33629\,
            I => \N__33598\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__33626\,
            I => \N__33594\
        );

    \I__7926\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33591\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__33622\,
            I => \N__33586\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__33619\,
            I => \N__33586\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__33616\,
            I => \N__33583\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__33611\,
            I => \N__33578\
        );

    \I__7921\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33571\
        );

    \I__7920\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33571\
        );

    \I__7919\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33571\
        );

    \I__7918\ : InMux
    port map (
            O => \N__33607\,
            I => \N__33568\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__33604\,
            I => \N__33565\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__33601\,
            I => \N__33558\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__33598\,
            I => \N__33555\
        );

    \I__7914\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33552\
        );

    \I__7913\ : Span4Mux_v
    port map (
            O => \N__33594\,
            I => \N__33547\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__33591\,
            I => \N__33547\
        );

    \I__7911\ : Span4Mux_v
    port map (
            O => \N__33586\,
            I => \N__33542\
        );

    \I__7910\ : Span4Mux_v
    port map (
            O => \N__33583\,
            I => \N__33542\
        );

    \I__7909\ : InMux
    port map (
            O => \N__33582\,
            I => \N__33539\
        );

    \I__7908\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33536\
        );

    \I__7907\ : Span4Mux_h
    port map (
            O => \N__33578\,
            I => \N__33533\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__33571\,
            I => \N__33530\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__33568\,
            I => \N__33525\
        );

    \I__7904\ : Span12Mux_s5_v
    port map (
            O => \N__33565\,
            I => \N__33525\
        );

    \I__7903\ : InMux
    port map (
            O => \N__33564\,
            I => \N__33516\
        );

    \I__7902\ : InMux
    port map (
            O => \N__33563\,
            I => \N__33516\
        );

    \I__7901\ : InMux
    port map (
            O => \N__33562\,
            I => \N__33516\
        );

    \I__7900\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33516\
        );

    \I__7899\ : Span4Mux_v
    port map (
            O => \N__33558\,
            I => \N__33505\
        );

    \I__7898\ : Span4Mux_h
    port map (
            O => \N__33555\,
            I => \N__33505\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__33552\,
            I => \N__33505\
        );

    \I__7896\ : Span4Mux_h
    port map (
            O => \N__33547\,
            I => \N__33505\
        );

    \I__7895\ : Span4Mux_h
    port map (
            O => \N__33542\,
            I => \N__33505\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__33539\,
            I => \tok.A_low_2\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__33536\,
            I => \tok.A_low_2\
        );

    \I__7892\ : Odrv4
    port map (
            O => \N__33533\,
            I => \tok.A_low_2\
        );

    \I__7891\ : Odrv12
    port map (
            O => \N__33530\,
            I => \tok.A_low_2\
        );

    \I__7890\ : Odrv12
    port map (
            O => \N__33525\,
            I => \tok.A_low_2\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__33516\,
            I => \tok.A_low_2\
        );

    \I__7888\ : Odrv4
    port map (
            O => \N__33505\,
            I => \tok.A_low_2\
        );

    \I__7887\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33486\
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__33489\,
            I => \N__33480\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__33486\,
            I => \N__33476\
        );

    \I__7884\ : InMux
    port map (
            O => \N__33485\,
            I => \N__33472\
        );

    \I__7883\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33468\
        );

    \I__7882\ : CascadeMux
    port map (
            O => \N__33483\,
            I => \N__33464\
        );

    \I__7881\ : InMux
    port map (
            O => \N__33480\,
            I => \N__33461\
        );

    \I__7880\ : InMux
    port map (
            O => \N__33479\,
            I => \N__33458\
        );

    \I__7879\ : Span4Mux_v
    port map (
            O => \N__33476\,
            I => \N__33455\
        );

    \I__7878\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33452\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__33472\,
            I => \N__33449\
        );

    \I__7876\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33446\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__33468\,
            I => \N__33442\
        );

    \I__7874\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33439\
        );

    \I__7873\ : InMux
    port map (
            O => \N__33464\,
            I => \N__33436\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__33461\,
            I => \N__33433\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__33458\,
            I => \N__33421\
        );

    \I__7870\ : Span4Mux_h
    port map (
            O => \N__33455\,
            I => \N__33421\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__33452\,
            I => \N__33421\
        );

    \I__7868\ : Span4Mux_v
    port map (
            O => \N__33449\,
            I => \N__33418\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__33446\,
            I => \N__33411\
        );

    \I__7866\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33408\
        );

    \I__7865\ : Span4Mux_s3_v
    port map (
            O => \N__33442\,
            I => \N__33405\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__33439\,
            I => \N__33400\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__33436\,
            I => \N__33400\
        );

    \I__7862\ : Span4Mux_v
    port map (
            O => \N__33433\,
            I => \N__33397\
        );

    \I__7861\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33394\
        );

    \I__7860\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33391\
        );

    \I__7859\ : InMux
    port map (
            O => \N__33430\,
            I => \N__33388\
        );

    \I__7858\ : InMux
    port map (
            O => \N__33429\,
            I => \N__33383\
        );

    \I__7857\ : InMux
    port map (
            O => \N__33428\,
            I => \N__33383\
        );

    \I__7856\ : Span4Mux_v
    port map (
            O => \N__33421\,
            I => \N__33378\
        );

    \I__7855\ : Span4Mux_v
    port map (
            O => \N__33418\,
            I => \N__33378\
        );

    \I__7854\ : InMux
    port map (
            O => \N__33417\,
            I => \N__33373\
        );

    \I__7853\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33373\
        );

    \I__7852\ : InMux
    port map (
            O => \N__33415\,
            I => \N__33368\
        );

    \I__7851\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33365\
        );

    \I__7850\ : Span4Mux_s3_v
    port map (
            O => \N__33411\,
            I => \N__33362\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__33408\,
            I => \N__33359\
        );

    \I__7848\ : Span4Mux_s3_h
    port map (
            O => \N__33405\,
            I => \N__33352\
        );

    \I__7847\ : Span4Mux_s3_h
    port map (
            O => \N__33400\,
            I => \N__33352\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__33397\,
            I => \N__33352\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__33394\,
            I => \N__33347\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__33391\,
            I => \N__33347\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__33388\,
            I => \N__33344\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__33383\,
            I => \N__33337\
        );

    \I__7841\ : Sp12to4
    port map (
            O => \N__33378\,
            I => \N__33337\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__33373\,
            I => \N__33337\
        );

    \I__7839\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33334\
        );

    \I__7838\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33331\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__33368\,
            I => \N__33326\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__33365\,
            I => \N__33326\
        );

    \I__7835\ : Span4Mux_h
    port map (
            O => \N__33362\,
            I => \N__33317\
        );

    \I__7834\ : Span4Mux_s2_h
    port map (
            O => \N__33359\,
            I => \N__33317\
        );

    \I__7833\ : Span4Mux_h
    port map (
            O => \N__33352\,
            I => \N__33317\
        );

    \I__7832\ : Span4Mux_s3_v
    port map (
            O => \N__33347\,
            I => \N__33317\
        );

    \I__7831\ : Span12Mux_s2_h
    port map (
            O => \N__33344\,
            I => \N__33312\
        );

    \I__7830\ : Span12Mux_s11_h
    port map (
            O => \N__33337\,
            I => \N__33312\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__33334\,
            I => \tok.n289\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__33331\,
            I => \tok.n289\
        );

    \I__7827\ : Odrv4
    port map (
            O => \N__33326\,
            I => \tok.n289\
        );

    \I__7826\ : Odrv4
    port map (
            O => \N__33317\,
            I => \tok.n289\
        );

    \I__7825\ : Odrv12
    port map (
            O => \N__33312\,
            I => \tok.n289\
        );

    \I__7824\ : CascadeMux
    port map (
            O => \N__33301\,
            I => \N__33284\
        );

    \I__7823\ : CascadeMux
    port map (
            O => \N__33300\,
            I => \N__33276\
        );

    \I__7822\ : CascadeMux
    port map (
            O => \N__33299\,
            I => \N__33260\
        );

    \I__7821\ : CascadeMux
    port map (
            O => \N__33298\,
            I => \N__33254\
        );

    \I__7820\ : CascadeMux
    port map (
            O => \N__33297\,
            I => \N__33245\
        );

    \I__7819\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33241\
        );

    \I__7818\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33237\
        );

    \I__7817\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33229\
        );

    \I__7816\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33224\
        );

    \I__7815\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33224\
        );

    \I__7814\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33220\
        );

    \I__7813\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33212\
        );

    \I__7812\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33212\
        );

    \I__7811\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33209\
        );

    \I__7810\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33206\
        );

    \I__7809\ : InMux
    port map (
            O => \N__33284\,
            I => \N__33199\
        );

    \I__7808\ : InMux
    port map (
            O => \N__33283\,
            I => \N__33199\
        );

    \I__7807\ : InMux
    port map (
            O => \N__33282\,
            I => \N__33199\
        );

    \I__7806\ : CascadeMux
    port map (
            O => \N__33281\,
            I => \N__33193\
        );

    \I__7805\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33187\
        );

    \I__7804\ : InMux
    port map (
            O => \N__33279\,
            I => \N__33176\
        );

    \I__7803\ : InMux
    port map (
            O => \N__33276\,
            I => \N__33176\
        );

    \I__7802\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33176\
        );

    \I__7801\ : InMux
    port map (
            O => \N__33274\,
            I => \N__33169\
        );

    \I__7800\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33169\
        );

    \I__7799\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33169\
        );

    \I__7798\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33154\
        );

    \I__7797\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33154\
        );

    \I__7796\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33154\
        );

    \I__7795\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33151\
        );

    \I__7794\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33148\
        );

    \I__7793\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33143\
        );

    \I__7792\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33143\
        );

    \I__7791\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33138\
        );

    \I__7790\ : InMux
    port map (
            O => \N__33263\,
            I => \N__33138\
        );

    \I__7789\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33130\
        );

    \I__7788\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33130\
        );

    \I__7787\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33125\
        );

    \I__7786\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33125\
        );

    \I__7785\ : InMux
    port map (
            O => \N__33254\,
            I => \N__33117\
        );

    \I__7784\ : InMux
    port map (
            O => \N__33253\,
            I => \N__33117\
        );

    \I__7783\ : InMux
    port map (
            O => \N__33252\,
            I => \N__33117\
        );

    \I__7782\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33110\
        );

    \I__7781\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33110\
        );

    \I__7780\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33110\
        );

    \I__7779\ : InMux
    port map (
            O => \N__33248\,
            I => \N__33103\
        );

    \I__7778\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33103\
        );

    \I__7777\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33103\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33094\
        );

    \I__7775\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33090\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__33237\,
            I => \N__33087\
        );

    \I__7773\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33084\
        );

    \I__7772\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33079\
        );

    \I__7771\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33079\
        );

    \I__7770\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33074\
        );

    \I__7769\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33074\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__33229\,
            I => \N__33069\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__33224\,
            I => \N__33069\
        );

    \I__7766\ : CascadeMux
    port map (
            O => \N__33223\,
            I => \N__33066\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__33220\,
            I => \N__33061\
        );

    \I__7764\ : InMux
    port map (
            O => \N__33219\,
            I => \N__33056\
        );

    \I__7763\ : InMux
    port map (
            O => \N__33218\,
            I => \N__33056\
        );

    \I__7762\ : InMux
    port map (
            O => \N__33217\,
            I => \N__33053\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__33212\,
            I => \N__33044\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__33209\,
            I => \N__33044\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__33206\,
            I => \N__33044\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__33199\,
            I => \N__33044\
        );

    \I__7757\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33041\
        );

    \I__7756\ : InMux
    port map (
            O => \N__33197\,
            I => \N__33032\
        );

    \I__7755\ : InMux
    port map (
            O => \N__33196\,
            I => \N__33032\
        );

    \I__7754\ : InMux
    port map (
            O => \N__33193\,
            I => \N__33032\
        );

    \I__7753\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33032\
        );

    \I__7752\ : InMux
    port map (
            O => \N__33191\,
            I => \N__33026\
        );

    \I__7751\ : InMux
    port map (
            O => \N__33190\,
            I => \N__33026\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__33187\,
            I => \N__33023\
        );

    \I__7749\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33015\
        );

    \I__7748\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33015\
        );

    \I__7747\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33015\
        );

    \I__7746\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33012\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__33176\,
            I => \N__33007\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__33169\,
            I => \N__33007\
        );

    \I__7743\ : InMux
    port map (
            O => \N__33168\,
            I => \N__33000\
        );

    \I__7742\ : InMux
    port map (
            O => \N__33167\,
            I => \N__33000\
        );

    \I__7741\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33000\
        );

    \I__7740\ : InMux
    port map (
            O => \N__33165\,
            I => \N__32995\
        );

    \I__7739\ : InMux
    port map (
            O => \N__33164\,
            I => \N__32995\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__33163\,
            I => \N__32992\
        );

    \I__7737\ : InMux
    port map (
            O => \N__33162\,
            I => \N__32989\
        );

    \I__7736\ : InMux
    port map (
            O => \N__33161\,
            I => \N__32986\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__33154\,
            I => \N__32983\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__33151\,
            I => \N__32978\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__33148\,
            I => \N__32978\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__33143\,
            I => \N__32973\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__33138\,
            I => \N__32973\
        );

    \I__7730\ : InMux
    port map (
            O => \N__33137\,
            I => \N__32968\
        );

    \I__7729\ : InMux
    port map (
            O => \N__33136\,
            I => \N__32968\
        );

    \I__7728\ : CascadeMux
    port map (
            O => \N__33135\,
            I => \N__32962\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__33130\,
            I => \N__32950\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__33125\,
            I => \N__32950\
        );

    \I__7725\ : InMux
    port map (
            O => \N__33124\,
            I => \N__32947\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__32944\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__33110\,
            I => \N__32941\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__33103\,
            I => \N__32938\
        );

    \I__7721\ : InMux
    port map (
            O => \N__33102\,
            I => \N__32935\
        );

    \I__7720\ : InMux
    port map (
            O => \N__33101\,
            I => \N__32932\
        );

    \I__7719\ : InMux
    port map (
            O => \N__33100\,
            I => \N__32929\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33099\,
            I => \N__32926\
        );

    \I__7717\ : InMux
    port map (
            O => \N__33098\,
            I => \N__32923\
        );

    \I__7716\ : InMux
    port map (
            O => \N__33097\,
            I => \N__32920\
        );

    \I__7715\ : Span4Mux_s3_v
    port map (
            O => \N__33094\,
            I => \N__32917\
        );

    \I__7714\ : InMux
    port map (
            O => \N__33093\,
            I => \N__32914\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__33090\,
            I => \N__32907\
        );

    \I__7712\ : Span4Mux_s3_v
    port map (
            O => \N__33087\,
            I => \N__32907\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__33084\,
            I => \N__32907\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__33079\,
            I => \N__32904\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__33074\,
            I => \N__32899\
        );

    \I__7708\ : Span4Mux_v
    port map (
            O => \N__33069\,
            I => \N__32899\
        );

    \I__7707\ : InMux
    port map (
            O => \N__33066\,
            I => \N__32892\
        );

    \I__7706\ : InMux
    port map (
            O => \N__33065\,
            I => \N__32892\
        );

    \I__7705\ : InMux
    port map (
            O => \N__33064\,
            I => \N__32892\
        );

    \I__7704\ : Span4Mux_v
    port map (
            O => \N__33061\,
            I => \N__32887\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__33056\,
            I => \N__32887\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__33053\,
            I => \N__32878\
        );

    \I__7701\ : Span4Mux_v
    port map (
            O => \N__33044\,
            I => \N__32878\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__33041\,
            I => \N__32878\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__33032\,
            I => \N__32878\
        );

    \I__7698\ : InMux
    port map (
            O => \N__33031\,
            I => \N__32874\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__33026\,
            I => \N__32869\
        );

    \I__7696\ : Span4Mux_v
    port map (
            O => \N__33023\,
            I => \N__32869\
        );

    \I__7695\ : InMux
    port map (
            O => \N__33022\,
            I => \N__32866\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__33015\,
            I => \N__32857\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__33012\,
            I => \N__32857\
        );

    \I__7692\ : Span4Mux_s3_v
    port map (
            O => \N__33007\,
            I => \N__32857\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__33000\,
            I => \N__32857\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__32995\,
            I => \N__32854\
        );

    \I__7689\ : InMux
    port map (
            O => \N__32992\,
            I => \N__32848\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__32989\,
            I => \N__32845\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__32986\,
            I => \N__32842\
        );

    \I__7686\ : Span4Mux_v
    port map (
            O => \N__32983\,
            I => \N__32833\
        );

    \I__7685\ : Span4Mux_s3_v
    port map (
            O => \N__32978\,
            I => \N__32833\
        );

    \I__7684\ : Span4Mux_h
    port map (
            O => \N__32973\,
            I => \N__32833\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__32968\,
            I => \N__32833\
        );

    \I__7682\ : InMux
    port map (
            O => \N__32967\,
            I => \N__32828\
        );

    \I__7681\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32828\
        );

    \I__7680\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32824\
        );

    \I__7679\ : InMux
    port map (
            O => \N__32962\,
            I => \N__32821\
        );

    \I__7678\ : InMux
    port map (
            O => \N__32961\,
            I => \N__32816\
        );

    \I__7677\ : InMux
    port map (
            O => \N__32960\,
            I => \N__32816\
        );

    \I__7676\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32811\
        );

    \I__7675\ : InMux
    port map (
            O => \N__32958\,
            I => \N__32811\
        );

    \I__7674\ : InMux
    port map (
            O => \N__32957\,
            I => \N__32804\
        );

    \I__7673\ : InMux
    port map (
            O => \N__32956\,
            I => \N__32804\
        );

    \I__7672\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32804\
        );

    \I__7671\ : Span4Mux_v
    port map (
            O => \N__32950\,
            I => \N__32799\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__32947\,
            I => \N__32799\
        );

    \I__7669\ : Span4Mux_v
    port map (
            O => \N__32944\,
            I => \N__32790\
        );

    \I__7668\ : Span4Mux_v
    port map (
            O => \N__32941\,
            I => \N__32790\
        );

    \I__7667\ : Span4Mux_s2_h
    port map (
            O => \N__32938\,
            I => \N__32790\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__32935\,
            I => \N__32790\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32782\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__32929\,
            I => \N__32775\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__32926\,
            I => \N__32766\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__32923\,
            I => \N__32766\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__32920\,
            I => \N__32766\
        );

    \I__7660\ : Span4Mux_v
    port map (
            O => \N__32917\,
            I => \N__32766\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__32914\,
            I => \N__32761\
        );

    \I__7658\ : Span4Mux_v
    port map (
            O => \N__32907\,
            I => \N__32761\
        );

    \I__7657\ : Span4Mux_v
    port map (
            O => \N__32904\,
            I => \N__32750\
        );

    \I__7656\ : Span4Mux_h
    port map (
            O => \N__32899\,
            I => \N__32750\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__32892\,
            I => \N__32750\
        );

    \I__7654\ : Span4Mux_s2_v
    port map (
            O => \N__32887\,
            I => \N__32750\
        );

    \I__7653\ : Span4Mux_v
    port map (
            O => \N__32878\,
            I => \N__32750\
        );

    \I__7652\ : InMux
    port map (
            O => \N__32877\,
            I => \N__32747\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__32874\,
            I => \N__32736\
        );

    \I__7650\ : Span4Mux_h
    port map (
            O => \N__32869\,
            I => \N__32736\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__32866\,
            I => \N__32736\
        );

    \I__7648\ : Span4Mux_v
    port map (
            O => \N__32857\,
            I => \N__32736\
        );

    \I__7647\ : Span4Mux_v
    port map (
            O => \N__32854\,
            I => \N__32736\
        );

    \I__7646\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32731\
        );

    \I__7645\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32731\
        );

    \I__7644\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32728\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__32848\,
            I => \N__32717\
        );

    \I__7642\ : Span4Mux_h
    port map (
            O => \N__32845\,
            I => \N__32717\
        );

    \I__7641\ : Span4Mux_s3_h
    port map (
            O => \N__32842\,
            I => \N__32717\
        );

    \I__7640\ : Span4Mux_h
    port map (
            O => \N__32833\,
            I => \N__32717\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__32828\,
            I => \N__32717\
        );

    \I__7638\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32714\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__32824\,
            I => \N__32711\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__32821\,
            I => \N__32708\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__32816\,
            I => \N__32701\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__32811\,
            I => \N__32701\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__32804\,
            I => \N__32701\
        );

    \I__7632\ : Span4Mux_s2_v
    port map (
            O => \N__32799\,
            I => \N__32696\
        );

    \I__7631\ : Span4Mux_v
    port map (
            O => \N__32790\,
            I => \N__32696\
        );

    \I__7630\ : InMux
    port map (
            O => \N__32789\,
            I => \N__32691\
        );

    \I__7629\ : InMux
    port map (
            O => \N__32788\,
            I => \N__32686\
        );

    \I__7628\ : InMux
    port map (
            O => \N__32787\,
            I => \N__32686\
        );

    \I__7627\ : InMux
    port map (
            O => \N__32786\,
            I => \N__32683\
        );

    \I__7626\ : InMux
    port map (
            O => \N__32785\,
            I => \N__32680\
        );

    \I__7625\ : Span12Mux_s11_v
    port map (
            O => \N__32782\,
            I => \N__32677\
        );

    \I__7624\ : InMux
    port map (
            O => \N__32781\,
            I => \N__32674\
        );

    \I__7623\ : InMux
    port map (
            O => \N__32780\,
            I => \N__32667\
        );

    \I__7622\ : InMux
    port map (
            O => \N__32779\,
            I => \N__32667\
        );

    \I__7621\ : InMux
    port map (
            O => \N__32778\,
            I => \N__32667\
        );

    \I__7620\ : Span4Mux_s2_v
    port map (
            O => \N__32775\,
            I => \N__32658\
        );

    \I__7619\ : Span4Mux_v
    port map (
            O => \N__32766\,
            I => \N__32658\
        );

    \I__7618\ : Span4Mux_v
    port map (
            O => \N__32761\,
            I => \N__32658\
        );

    \I__7617\ : Span4Mux_h
    port map (
            O => \N__32750\,
            I => \N__32658\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__32747\,
            I => \N__32651\
        );

    \I__7615\ : Span4Mux_h
    port map (
            O => \N__32736\,
            I => \N__32651\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__32731\,
            I => \N__32651\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__32728\,
            I => \N__32644\
        );

    \I__7612\ : Span4Mux_v
    port map (
            O => \N__32717\,
            I => \N__32644\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__32714\,
            I => \N__32644\
        );

    \I__7610\ : Span4Mux_s2_v
    port map (
            O => \N__32711\,
            I => \N__32635\
        );

    \I__7609\ : Span4Mux_s2_v
    port map (
            O => \N__32708\,
            I => \N__32635\
        );

    \I__7608\ : Span4Mux_v
    port map (
            O => \N__32701\,
            I => \N__32635\
        );

    \I__7607\ : Span4Mux_h
    port map (
            O => \N__32696\,
            I => \N__32635\
        );

    \I__7606\ : InMux
    port map (
            O => \N__32695\,
            I => \N__32630\
        );

    \I__7605\ : InMux
    port map (
            O => \N__32694\,
            I => \N__32630\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__32691\,
            I => \tok.T_1\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__32686\,
            I => \tok.T_1\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__32683\,
            I => \tok.T_1\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__32680\,
            I => \tok.T_1\
        );

    \I__7600\ : Odrv12
    port map (
            O => \N__32677\,
            I => \tok.T_1\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__32674\,
            I => \tok.T_1\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__32667\,
            I => \tok.T_1\
        );

    \I__7597\ : Odrv4
    port map (
            O => \N__32658\,
            I => \tok.T_1\
        );

    \I__7596\ : Odrv4
    port map (
            O => \N__32651\,
            I => \tok.T_1\
        );

    \I__7595\ : Odrv4
    port map (
            O => \N__32644\,
            I => \tok.T_1\
        );

    \I__7594\ : Odrv4
    port map (
            O => \N__32635\,
            I => \tok.T_1\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__32630\,
            I => \tok.T_1\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__32605\,
            I => \N__32602\
        );

    \I__7591\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32598\
        );

    \I__7590\ : InMux
    port map (
            O => \N__32601\,
            I => \N__32595\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__32598\,
            I => \N__32590\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__32595\,
            I => \N__32587\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__32594\,
            I => \N__32582\
        );

    \I__7586\ : CascadeMux
    port map (
            O => \N__32593\,
            I => \N__32578\
        );

    \I__7585\ : Span4Mux_h
    port map (
            O => \N__32590\,
            I => \N__32573\
        );

    \I__7584\ : Span4Mux_h
    port map (
            O => \N__32587\,
            I => \N__32573\
        );

    \I__7583\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32570\
        );

    \I__7582\ : InMux
    port map (
            O => \N__32585\,
            I => \N__32565\
        );

    \I__7581\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32565\
        );

    \I__7580\ : InMux
    port map (
            O => \N__32581\,
            I => \N__32560\
        );

    \I__7579\ : InMux
    port map (
            O => \N__32578\,
            I => \N__32560\
        );

    \I__7578\ : Odrv4
    port map (
            O => \N__32573\,
            I => \tok.n222\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__32570\,
            I => \tok.n222\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__32565\,
            I => \tok.n222\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__32560\,
            I => \tok.n222\
        );

    \I__7574\ : InMux
    port map (
            O => \N__32551\,
            I => \N__32544\
        );

    \I__7573\ : InMux
    port map (
            O => \N__32550\,
            I => \N__32541\
        );

    \I__7572\ : InMux
    port map (
            O => \N__32549\,
            I => \N__32538\
        );

    \I__7571\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32535\
        );

    \I__7570\ : InMux
    port map (
            O => \N__32547\,
            I => \N__32532\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__32544\,
            I => \N__32529\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__32541\,
            I => \N__32526\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__32538\,
            I => \N__32523\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__32535\,
            I => \N__32520\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__32532\,
            I => \N__32517\
        );

    \I__7564\ : Span4Mux_v
    port map (
            O => \N__32529\,
            I => \N__32514\
        );

    \I__7563\ : Span4Mux_v
    port map (
            O => \N__32526\,
            I => \N__32509\
        );

    \I__7562\ : Span4Mux_v
    port map (
            O => \N__32523\,
            I => \N__32509\
        );

    \I__7561\ : Span4Mux_s2_h
    port map (
            O => \N__32520\,
            I => \N__32506\
        );

    \I__7560\ : Span4Mux_v
    port map (
            O => \N__32517\,
            I => \N__32503\
        );

    \I__7559\ : Span4Mux_v
    port map (
            O => \N__32514\,
            I => \N__32498\
        );

    \I__7558\ : Span4Mux_h
    port map (
            O => \N__32509\,
            I => \N__32498\
        );

    \I__7557\ : Span4Mux_h
    port map (
            O => \N__32506\,
            I => \N__32495\
        );

    \I__7556\ : Span4Mux_h
    port map (
            O => \N__32503\,
            I => \N__32492\
        );

    \I__7555\ : Odrv4
    port map (
            O => \N__32498\,
            I => \tok.n838\
        );

    \I__7554\ : Odrv4
    port map (
            O => \N__32495\,
            I => \tok.n838\
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__32492\,
            I => \tok.n838\
        );

    \I__7552\ : CascadeMux
    port map (
            O => \N__32485\,
            I => \tok.n863_cascade_\
        );

    \I__7551\ : InMux
    port map (
            O => \N__32482\,
            I => \N__32479\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__32479\,
            I => \tok.n6472\
        );

    \I__7549\ : InMux
    port map (
            O => \N__32476\,
            I => \N__32473\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__32473\,
            I => \N__32466\
        );

    \I__7547\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32461\
        );

    \I__7546\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32461\
        );

    \I__7545\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32457\
        );

    \I__7544\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32454\
        );

    \I__7543\ : Span4Mux_v
    port map (
            O => \N__32466\,
            I => \N__32449\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__32461\,
            I => \N__32449\
        );

    \I__7541\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32446\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__32457\,
            I => \N__32443\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__32454\,
            I => \N__32438\
        );

    \I__7538\ : Span4Mux_v
    port map (
            O => \N__32449\,
            I => \N__32438\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__32446\,
            I => \N__32435\
        );

    \I__7536\ : Span4Mux_h
    port map (
            O => \N__32443\,
            I => \N__32426\
        );

    \I__7535\ : Span4Mux_h
    port map (
            O => \N__32438\,
            I => \N__32426\
        );

    \I__7534\ : Span4Mux_v
    port map (
            O => \N__32435\,
            I => \N__32426\
        );

    \I__7533\ : InMux
    port map (
            O => \N__32434\,
            I => \N__32421\
        );

    \I__7532\ : InMux
    port map (
            O => \N__32433\,
            I => \N__32421\
        );

    \I__7531\ : Span4Mux_h
    port map (
            O => \N__32426\,
            I => \N__32418\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__32421\,
            I => \N__32415\
        );

    \I__7529\ : Span4Mux_h
    port map (
            O => \N__32418\,
            I => \N__32412\
        );

    \I__7528\ : Odrv12
    port map (
            O => \N__32415\,
            I => \tok.n9_adj_677\
        );

    \I__7527\ : Odrv4
    port map (
            O => \N__32412\,
            I => \tok.n9_adj_677\
        );

    \I__7526\ : InMux
    port map (
            O => \N__32407\,
            I => \N__32404\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__32404\,
            I => \N__32401\
        );

    \I__7524\ : Span4Mux_v
    port map (
            O => \N__32401\,
            I => \N__32397\
        );

    \I__7523\ : InMux
    port map (
            O => \N__32400\,
            I => \N__32394\
        );

    \I__7522\ : Span4Mux_h
    port map (
            O => \N__32397\,
            I => \N__32391\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__32394\,
            I => \tok.n205\
        );

    \I__7520\ : Odrv4
    port map (
            O => \N__32391\,
            I => \tok.n205\
        );

    \I__7519\ : InMux
    port map (
            O => \N__32386\,
            I => \N__32383\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__32383\,
            I => \tok.n6477\
        );

    \I__7517\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32374\
        );

    \I__7516\ : InMux
    port map (
            O => \N__32379\,
            I => \N__32369\
        );

    \I__7515\ : InMux
    port map (
            O => \N__32378\,
            I => \N__32363\
        );

    \I__7514\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32363\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__32374\,
            I => \N__32360\
        );

    \I__7512\ : CascadeMux
    port map (
            O => \N__32373\,
            I => \N__32357\
        );

    \I__7511\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32351\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__32369\,
            I => \N__32348\
        );

    \I__7509\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32345\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__32363\,
            I => \N__32342\
        );

    \I__7507\ : Span4Mux_s3_v
    port map (
            O => \N__32360\,
            I => \N__32339\
        );

    \I__7506\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32336\
        );

    \I__7505\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32331\
        );

    \I__7504\ : InMux
    port map (
            O => \N__32355\,
            I => \N__32331\
        );

    \I__7503\ : InMux
    port map (
            O => \N__32354\,
            I => \N__32327\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__32351\,
            I => \N__32324\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__32348\,
            I => \N__32319\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__32345\,
            I => \N__32319\
        );

    \I__7499\ : Span4Mux_v
    port map (
            O => \N__32342\,
            I => \N__32316\
        );

    \I__7498\ : Span4Mux_v
    port map (
            O => \N__32339\,
            I => \N__32313\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__32336\,
            I => \N__32308\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__32331\,
            I => \N__32308\
        );

    \I__7495\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32305\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__32327\,
            I => \N__32302\
        );

    \I__7493\ : Span4Mux_v
    port map (
            O => \N__32324\,
            I => \N__32295\
        );

    \I__7492\ : Span4Mux_v
    port map (
            O => \N__32319\,
            I => \N__32295\
        );

    \I__7491\ : Span4Mux_h
    port map (
            O => \N__32316\,
            I => \N__32295\
        );

    \I__7490\ : Span4Mux_h
    port map (
            O => \N__32313\,
            I => \N__32290\
        );

    \I__7489\ : Span4Mux_h
    port map (
            O => \N__32308\,
            I => \N__32290\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__32305\,
            I => \tok.n43\
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__32302\,
            I => \tok.n43\
        );

    \I__7486\ : Odrv4
    port map (
            O => \N__32295\,
            I => \tok.n43\
        );

    \I__7485\ : Odrv4
    port map (
            O => \N__32290\,
            I => \tok.n43\
        );

    \I__7484\ : InMux
    port map (
            O => \N__32281\,
            I => \N__32278\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__32278\,
            I => \N__32275\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__32275\,
            I => \N__32271\
        );

    \I__7481\ : CascadeMux
    port map (
            O => \N__32274\,
            I => \N__32268\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__32271\,
            I => \N__32265\
        );

    \I__7479\ : InMux
    port map (
            O => \N__32268\,
            I => \N__32262\
        );

    \I__7478\ : Span4Mux_h
    port map (
            O => \N__32265\,
            I => \N__32259\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__32262\,
            I => \N__32256\
        );

    \I__7476\ : Odrv4
    port map (
            O => \N__32259\,
            I => \tok.n311\
        );

    \I__7475\ : Odrv12
    port map (
            O => \N__32256\,
            I => \tok.n311\
        );

    \I__7474\ : CascadeMux
    port map (
            O => \N__32251\,
            I => \N__32248\
        );

    \I__7473\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32244\
        );

    \I__7472\ : InMux
    port map (
            O => \N__32247\,
            I => \N__32241\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__32244\,
            I => \N__32236\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__32241\,
            I => \N__32236\
        );

    \I__7469\ : Odrv12
    port map (
            O => \N__32236\,
            I => \tok.n190_adj_797\
        );

    \I__7468\ : InMux
    port map (
            O => \N__32233\,
            I => \N__32227\
        );

    \I__7467\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32224\
        );

    \I__7466\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32221\
        );

    \I__7465\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32217\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__32227\,
            I => \N__32214\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__32224\,
            I => \N__32211\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__32221\,
            I => \N__32207\
        );

    \I__7461\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32204\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__32217\,
            I => \N__32201\
        );

    \I__7459\ : Span4Mux_h
    port map (
            O => \N__32214\,
            I => \N__32197\
        );

    \I__7458\ : Span4Mux_v
    port map (
            O => \N__32211\,
            I => \N__32194\
        );

    \I__7457\ : InMux
    port map (
            O => \N__32210\,
            I => \N__32191\
        );

    \I__7456\ : Span4Mux_h
    port map (
            O => \N__32207\,
            I => \N__32183\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__32204\,
            I => \N__32183\
        );

    \I__7454\ : Span4Mux_h
    port map (
            O => \N__32201\,
            I => \N__32180\
        );

    \I__7453\ : InMux
    port map (
            O => \N__32200\,
            I => \N__32177\
        );

    \I__7452\ : Span4Mux_v
    port map (
            O => \N__32197\,
            I => \N__32170\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__32194\,
            I => \N__32170\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__32191\,
            I => \N__32170\
        );

    \I__7449\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32164\
        );

    \I__7448\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32164\
        );

    \I__7447\ : InMux
    port map (
            O => \N__32188\,
            I => \N__32161\
        );

    \I__7446\ : Span4Mux_h
    port map (
            O => \N__32183\,
            I => \N__32154\
        );

    \I__7445\ : Span4Mux_h
    port map (
            O => \N__32180\,
            I => \N__32154\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__32177\,
            I => \N__32154\
        );

    \I__7443\ : Span4Mux_h
    port map (
            O => \N__32170\,
            I => \N__32151\
        );

    \I__7442\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32148\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__32164\,
            I => \N__32145\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__32161\,
            I => \tok.n44\
        );

    \I__7439\ : Odrv4
    port map (
            O => \N__32154\,
            I => \tok.n44\
        );

    \I__7438\ : Odrv4
    port map (
            O => \N__32151\,
            I => \tok.n44\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__32148\,
            I => \tok.n44\
        );

    \I__7436\ : Odrv12
    port map (
            O => \N__32145\,
            I => \tok.n44\
        );

    \I__7435\ : CascadeMux
    port map (
            O => \N__32134\,
            I => \N__32128\
        );

    \I__7434\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32101\
        );

    \I__7433\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32101\
        );

    \I__7432\ : CascadeMux
    port map (
            O => \N__32131\,
            I => \N__32088\
        );

    \I__7431\ : InMux
    port map (
            O => \N__32128\,
            I => \N__32084\
        );

    \I__7430\ : InMux
    port map (
            O => \N__32127\,
            I => \N__32081\
        );

    \I__7429\ : CascadeMux
    port map (
            O => \N__32126\,
            I => \N__32072\
        );

    \I__7428\ : InMux
    port map (
            O => \N__32125\,
            I => \N__32066\
        );

    \I__7427\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32066\
        );

    \I__7426\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32060\
        );

    \I__7425\ : InMux
    port map (
            O => \N__32122\,
            I => \N__32056\
        );

    \I__7424\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32053\
        );

    \I__7423\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32046\
        );

    \I__7422\ : InMux
    port map (
            O => \N__32119\,
            I => \N__32046\
        );

    \I__7421\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32046\
        );

    \I__7420\ : CascadeMux
    port map (
            O => \N__32117\,
            I => \N__32038\
        );

    \I__7419\ : CascadeMux
    port map (
            O => \N__32116\,
            I => \N__32035\
        );

    \I__7418\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32030\
        );

    \I__7417\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32025\
        );

    \I__7416\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32025\
        );

    \I__7415\ : CascadeMux
    port map (
            O => \N__32112\,
            I => \N__32015\
        );

    \I__7414\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32012\
        );

    \I__7413\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32005\
        );

    \I__7412\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32005\
        );

    \I__7411\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32005\
        );

    \I__7410\ : InMux
    port map (
            O => \N__32107\,
            I => \N__32002\
        );

    \I__7409\ : InMux
    port map (
            O => \N__32106\,
            I => \N__31999\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__32101\,
            I => \N__31996\
        );

    \I__7407\ : InMux
    port map (
            O => \N__32100\,
            I => \N__31989\
        );

    \I__7406\ : InMux
    port map (
            O => \N__32099\,
            I => \N__31989\
        );

    \I__7405\ : InMux
    port map (
            O => \N__32098\,
            I => \N__31989\
        );

    \I__7404\ : InMux
    port map (
            O => \N__32097\,
            I => \N__31982\
        );

    \I__7403\ : InMux
    port map (
            O => \N__32096\,
            I => \N__31982\
        );

    \I__7402\ : InMux
    port map (
            O => \N__32095\,
            I => \N__31982\
        );

    \I__7401\ : CascadeMux
    port map (
            O => \N__32094\,
            I => \N__31975\
        );

    \I__7400\ : InMux
    port map (
            O => \N__32093\,
            I => \N__31968\
        );

    \I__7399\ : InMux
    port map (
            O => \N__32092\,
            I => \N__31968\
        );

    \I__7398\ : InMux
    port map (
            O => \N__32091\,
            I => \N__31961\
        );

    \I__7397\ : InMux
    port map (
            O => \N__32088\,
            I => \N__31961\
        );

    \I__7396\ : InMux
    port map (
            O => \N__32087\,
            I => \N__31961\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__32084\,
            I => \N__31950\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__32081\,
            I => \N__31950\
        );

    \I__7393\ : InMux
    port map (
            O => \N__32080\,
            I => \N__31945\
        );

    \I__7392\ : InMux
    port map (
            O => \N__32079\,
            I => \N__31945\
        );

    \I__7391\ : InMux
    port map (
            O => \N__32078\,
            I => \N__31928\
        );

    \I__7390\ : InMux
    port map (
            O => \N__32077\,
            I => \N__31923\
        );

    \I__7389\ : InMux
    port map (
            O => \N__32076\,
            I => \N__31923\
        );

    \I__7388\ : CascadeMux
    port map (
            O => \N__32075\,
            I => \N__31909\
        );

    \I__7387\ : InMux
    port map (
            O => \N__32072\,
            I => \N__31902\
        );

    \I__7386\ : InMux
    port map (
            O => \N__32071\,
            I => \N__31899\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__32066\,
            I => \N__31893\
        );

    \I__7384\ : InMux
    port map (
            O => \N__32065\,
            I => \N__31886\
        );

    \I__7383\ : InMux
    port map (
            O => \N__32064\,
            I => \N__31886\
        );

    \I__7382\ : InMux
    port map (
            O => \N__32063\,
            I => \N__31886\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__32060\,
            I => \N__31881\
        );

    \I__7380\ : InMux
    port map (
            O => \N__32059\,
            I => \N__31872\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__32056\,
            I => \N__31865\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__32053\,
            I => \N__31865\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__32046\,
            I => \N__31865\
        );

    \I__7376\ : InMux
    port map (
            O => \N__32045\,
            I => \N__31858\
        );

    \I__7375\ : InMux
    port map (
            O => \N__32044\,
            I => \N__31858\
        );

    \I__7374\ : InMux
    port map (
            O => \N__32043\,
            I => \N__31858\
        );

    \I__7373\ : InMux
    port map (
            O => \N__32042\,
            I => \N__31855\
        );

    \I__7372\ : InMux
    port map (
            O => \N__32041\,
            I => \N__31844\
        );

    \I__7371\ : InMux
    port map (
            O => \N__32038\,
            I => \N__31844\
        );

    \I__7370\ : InMux
    port map (
            O => \N__32035\,
            I => \N__31844\
        );

    \I__7369\ : InMux
    port map (
            O => \N__32034\,
            I => \N__31844\
        );

    \I__7368\ : InMux
    port map (
            O => \N__32033\,
            I => \N__31844\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__32030\,
            I => \N__31839\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__32025\,
            I => \N__31839\
        );

    \I__7365\ : InMux
    port map (
            O => \N__32024\,
            I => \N__31834\
        );

    \I__7364\ : InMux
    port map (
            O => \N__32023\,
            I => \N__31834\
        );

    \I__7363\ : InMux
    port map (
            O => \N__32022\,
            I => \N__31829\
        );

    \I__7362\ : InMux
    port map (
            O => \N__32021\,
            I => \N__31829\
        );

    \I__7361\ : InMux
    port map (
            O => \N__32020\,
            I => \N__31823\
        );

    \I__7360\ : InMux
    port map (
            O => \N__32019\,
            I => \N__31818\
        );

    \I__7359\ : InMux
    port map (
            O => \N__32018\,
            I => \N__31818\
        );

    \I__7358\ : InMux
    port map (
            O => \N__32015\,
            I => \N__31815\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__32012\,
            I => \N__31810\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__32005\,
            I => \N__31810\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__32002\,
            I => \N__31801\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__31999\,
            I => \N__31801\
        );

    \I__7353\ : Span4Mux_s2_h
    port map (
            O => \N__31996\,
            I => \N__31801\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__31989\,
            I => \N__31801\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31798\
        );

    \I__7350\ : InMux
    port map (
            O => \N__31981\,
            I => \N__31789\
        );

    \I__7349\ : InMux
    port map (
            O => \N__31980\,
            I => \N__31789\
        );

    \I__7348\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31789\
        );

    \I__7347\ : InMux
    port map (
            O => \N__31978\,
            I => \N__31789\
        );

    \I__7346\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31782\
        );

    \I__7345\ : InMux
    port map (
            O => \N__31974\,
            I => \N__31782\
        );

    \I__7344\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31782\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__31968\,
            I => \N__31779\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__31961\,
            I => \N__31776\
        );

    \I__7341\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31769\
        );

    \I__7340\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31769\
        );

    \I__7339\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31769\
        );

    \I__7338\ : CascadeMux
    port map (
            O => \N__31957\,
            I => \N__31766\
        );

    \I__7337\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31762\
        );

    \I__7336\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31759\
        );

    \I__7335\ : Span4Mux_s2_h
    port map (
            O => \N__31950\,
            I => \N__31756\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__31945\,
            I => \N__31753\
        );

    \I__7333\ : InMux
    port map (
            O => \N__31944\,
            I => \N__31746\
        );

    \I__7332\ : InMux
    port map (
            O => \N__31943\,
            I => \N__31746\
        );

    \I__7331\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31746\
        );

    \I__7330\ : InMux
    port map (
            O => \N__31941\,
            I => \N__31738\
        );

    \I__7329\ : InMux
    port map (
            O => \N__31940\,
            I => \N__31738\
        );

    \I__7328\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31735\
        );

    \I__7327\ : InMux
    port map (
            O => \N__31938\,
            I => \N__31730\
        );

    \I__7326\ : InMux
    port map (
            O => \N__31937\,
            I => \N__31730\
        );

    \I__7325\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31725\
        );

    \I__7324\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31725\
        );

    \I__7323\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31720\
        );

    \I__7322\ : InMux
    port map (
            O => \N__31933\,
            I => \N__31720\
        );

    \I__7321\ : InMux
    port map (
            O => \N__31932\,
            I => \N__31715\
        );

    \I__7320\ : InMux
    port map (
            O => \N__31931\,
            I => \N__31715\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__31928\,
            I => \N__31712\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__31923\,
            I => \N__31709\
        );

    \I__7317\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31704\
        );

    \I__7316\ : InMux
    port map (
            O => \N__31921\,
            I => \N__31704\
        );

    \I__7315\ : InMux
    port map (
            O => \N__31920\,
            I => \N__31699\
        );

    \I__7314\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31699\
        );

    \I__7313\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31694\
        );

    \I__7312\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31694\
        );

    \I__7311\ : InMux
    port map (
            O => \N__31916\,
            I => \N__31691\
        );

    \I__7310\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31682\
        );

    \I__7309\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31682\
        );

    \I__7308\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31682\
        );

    \I__7307\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31682\
        );

    \I__7306\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31679\
        );

    \I__7305\ : InMux
    port map (
            O => \N__31908\,
            I => \N__31676\
        );

    \I__7304\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31673\
        );

    \I__7303\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31666\
        );

    \I__7302\ : InMux
    port map (
            O => \N__31905\,
            I => \N__31666\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__31902\,
            I => \N__31661\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__31899\,
            I => \N__31661\
        );

    \I__7299\ : InMux
    port map (
            O => \N__31898\,
            I => \N__31658\
        );

    \I__7298\ : InMux
    port map (
            O => \N__31897\,
            I => \N__31653\
        );

    \I__7297\ : InMux
    port map (
            O => \N__31896\,
            I => \N__31653\
        );

    \I__7296\ : Span4Mux_v
    port map (
            O => \N__31893\,
            I => \N__31650\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__31886\,
            I => \N__31647\
        );

    \I__7294\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31642\
        );

    \I__7293\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31642\
        );

    \I__7292\ : Span4Mux_v
    port map (
            O => \N__31881\,
            I => \N__31639\
        );

    \I__7291\ : InMux
    port map (
            O => \N__31880\,
            I => \N__31634\
        );

    \I__7290\ : InMux
    port map (
            O => \N__31879\,
            I => \N__31634\
        );

    \I__7289\ : InMux
    port map (
            O => \N__31878\,
            I => \N__31625\
        );

    \I__7288\ : InMux
    port map (
            O => \N__31877\,
            I => \N__31625\
        );

    \I__7287\ : InMux
    port map (
            O => \N__31876\,
            I => \N__31625\
        );

    \I__7286\ : InMux
    port map (
            O => \N__31875\,
            I => \N__31625\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__31872\,
            I => \N__31618\
        );

    \I__7284\ : Span4Mux_h
    port map (
            O => \N__31865\,
            I => \N__31618\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__31858\,
            I => \N__31618\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__31855\,
            I => \N__31611\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__31844\,
            I => \N__31611\
        );

    \I__7280\ : Span4Mux_s2_h
    port map (
            O => \N__31839\,
            I => \N__31611\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__31834\,
            I => \N__31606\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__31829\,
            I => \N__31606\
        );

    \I__7277\ : InMux
    port map (
            O => \N__31828\,
            I => \N__31601\
        );

    \I__7276\ : InMux
    port map (
            O => \N__31827\,
            I => \N__31601\
        );

    \I__7275\ : InMux
    port map (
            O => \N__31826\,
            I => \N__31598\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__31823\,
            I => \N__31593\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__31818\,
            I => \N__31593\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__31815\,
            I => \N__31582\
        );

    \I__7271\ : Span4Mux_h
    port map (
            O => \N__31810\,
            I => \N__31582\
        );

    \I__7270\ : Span4Mux_h
    port map (
            O => \N__31801\,
            I => \N__31582\
        );

    \I__7269\ : Span4Mux_v
    port map (
            O => \N__31798\,
            I => \N__31582\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__31789\,
            I => \N__31582\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__31782\,
            I => \N__31573\
        );

    \I__7266\ : Span4Mux_v
    port map (
            O => \N__31779\,
            I => \N__31573\
        );

    \I__7265\ : Span4Mux_s2_h
    port map (
            O => \N__31776\,
            I => \N__31573\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__31769\,
            I => \N__31573\
        );

    \I__7263\ : InMux
    port map (
            O => \N__31766\,
            I => \N__31569\
        );

    \I__7262\ : InMux
    port map (
            O => \N__31765\,
            I => \N__31566\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__31762\,
            I => \N__31555\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__31759\,
            I => \N__31555\
        );

    \I__7259\ : Span4Mux_v
    port map (
            O => \N__31756\,
            I => \N__31555\
        );

    \I__7258\ : Span4Mux_s3_v
    port map (
            O => \N__31753\,
            I => \N__31555\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__31746\,
            I => \N__31555\
        );

    \I__7256\ : InMux
    port map (
            O => \N__31745\,
            I => \N__31550\
        );

    \I__7255\ : InMux
    port map (
            O => \N__31744\,
            I => \N__31550\
        );

    \I__7254\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31542\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__31738\,
            I => \N__31539\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__31735\,
            I => \N__31535\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__31730\,
            I => \N__31528\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__31725\,
            I => \N__31528\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__31720\,
            I => \N__31528\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__31715\,
            I => \N__31525\
        );

    \I__7247\ : Span4Mux_s3_h
    port map (
            O => \N__31712\,
            I => \N__31520\
        );

    \I__7246\ : Span4Mux_v
    port map (
            O => \N__31709\,
            I => \N__31520\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__31704\,
            I => \N__31513\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__31699\,
            I => \N__31513\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__31694\,
            I => \N__31513\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__31691\,
            I => \N__31510\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__31682\,
            I => \N__31507\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__31679\,
            I => \N__31504\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__31676\,
            I => \N__31499\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__31673\,
            I => \N__31499\
        );

    \I__7237\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31494\
        );

    \I__7236\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31494\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__31666\,
            I => \N__31487\
        );

    \I__7234\ : Span4Mux_v
    port map (
            O => \N__31661\,
            I => \N__31487\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__31658\,
            I => \N__31487\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__31653\,
            I => \N__31476\
        );

    \I__7231\ : Span4Mux_v
    port map (
            O => \N__31650\,
            I => \N__31476\
        );

    \I__7230\ : Span4Mux_s2_v
    port map (
            O => \N__31647\,
            I => \N__31476\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__31642\,
            I => \N__31476\
        );

    \I__7228\ : Span4Mux_v
    port map (
            O => \N__31639\,
            I => \N__31476\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__31634\,
            I => \N__31471\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__31625\,
            I => \N__31471\
        );

    \I__7225\ : Span4Mux_v
    port map (
            O => \N__31618\,
            I => \N__31463\
        );

    \I__7224\ : Span4Mux_h
    port map (
            O => \N__31611\,
            I => \N__31463\
        );

    \I__7223\ : Span4Mux_h
    port map (
            O => \N__31606\,
            I => \N__31458\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__31601\,
            I => \N__31458\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__31598\,
            I => \N__31455\
        );

    \I__7220\ : Span4Mux_v
    port map (
            O => \N__31593\,
            I => \N__31448\
        );

    \I__7219\ : Span4Mux_v
    port map (
            O => \N__31582\,
            I => \N__31448\
        );

    \I__7218\ : Span4Mux_h
    port map (
            O => \N__31573\,
            I => \N__31448\
        );

    \I__7217\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31445\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__31569\,
            I => \N__31436\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__31566\,
            I => \N__31436\
        );

    \I__7214\ : Sp12to4
    port map (
            O => \N__31555\,
            I => \N__31436\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__31550\,
            I => \N__31436\
        );

    \I__7212\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31431\
        );

    \I__7211\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31431\
        );

    \I__7210\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31428\
        );

    \I__7209\ : InMux
    port map (
            O => \N__31546\,
            I => \N__31423\
        );

    \I__7208\ : InMux
    port map (
            O => \N__31545\,
            I => \N__31423\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__31542\,
            I => \N__31420\
        );

    \I__7206\ : Span4Mux_v
    port map (
            O => \N__31539\,
            I => \N__31417\
        );

    \I__7205\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31414\
        );

    \I__7204\ : Span12Mux_s3_h
    port map (
            O => \N__31535\,
            I => \N__31409\
        );

    \I__7203\ : Span12Mux_s10_h
    port map (
            O => \N__31528\,
            I => \N__31409\
        );

    \I__7202\ : Span4Mux_v
    port map (
            O => \N__31525\,
            I => \N__31398\
        );

    \I__7201\ : Span4Mux_h
    port map (
            O => \N__31520\,
            I => \N__31398\
        );

    \I__7200\ : Span4Mux_v
    port map (
            O => \N__31513\,
            I => \N__31398\
        );

    \I__7199\ : Span4Mux_s2_v
    port map (
            O => \N__31510\,
            I => \N__31398\
        );

    \I__7198\ : Span4Mux_v
    port map (
            O => \N__31507\,
            I => \N__31398\
        );

    \I__7197\ : Span4Mux_v
    port map (
            O => \N__31504\,
            I => \N__31389\
        );

    \I__7196\ : Span4Mux_v
    port map (
            O => \N__31499\,
            I => \N__31389\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__31494\,
            I => \N__31389\
        );

    \I__7194\ : Span4Mux_h
    port map (
            O => \N__31487\,
            I => \N__31389\
        );

    \I__7193\ : Sp12to4
    port map (
            O => \N__31476\,
            I => \N__31384\
        );

    \I__7192\ : Span12Mux_s11_v
    port map (
            O => \N__31471\,
            I => \N__31384\
        );

    \I__7191\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31377\
        );

    \I__7190\ : InMux
    port map (
            O => \N__31469\,
            I => \N__31377\
        );

    \I__7189\ : InMux
    port map (
            O => \N__31468\,
            I => \N__31377\
        );

    \I__7188\ : Span4Mux_h
    port map (
            O => \N__31463\,
            I => \N__31372\
        );

    \I__7187\ : Span4Mux_v
    port map (
            O => \N__31458\,
            I => \N__31372\
        );

    \I__7186\ : Span4Mux_v
    port map (
            O => \N__31455\,
            I => \N__31365\
        );

    \I__7185\ : Span4Mux_h
    port map (
            O => \N__31448\,
            I => \N__31365\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__31445\,
            I => \N__31365\
        );

    \I__7183\ : Span12Mux_s10_h
    port map (
            O => \N__31436\,
            I => \N__31362\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__31431\,
            I => \tok.T_2\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__31428\,
            I => \tok.T_2\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__31423\,
            I => \tok.T_2\
        );

    \I__7179\ : Odrv4
    port map (
            O => \N__31420\,
            I => \tok.T_2\
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__31417\,
            I => \tok.T_2\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__31414\,
            I => \tok.T_2\
        );

    \I__7176\ : Odrv12
    port map (
            O => \N__31409\,
            I => \tok.T_2\
        );

    \I__7175\ : Odrv4
    port map (
            O => \N__31398\,
            I => \tok.T_2\
        );

    \I__7174\ : Odrv4
    port map (
            O => \N__31389\,
            I => \tok.T_2\
        );

    \I__7173\ : Odrv12
    port map (
            O => \N__31384\,
            I => \tok.T_2\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__31377\,
            I => \tok.T_2\
        );

    \I__7171\ : Odrv4
    port map (
            O => \N__31372\,
            I => \tok.T_2\
        );

    \I__7170\ : Odrv4
    port map (
            O => \N__31365\,
            I => \tok.T_2\
        );

    \I__7169\ : Odrv12
    port map (
            O => \N__31362\,
            I => \tok.T_2\
        );

    \I__7168\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31291\
        );

    \I__7167\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31291\
        );

    \I__7166\ : InMux
    port map (
            O => \N__31331\,
            I => \N__31286\
        );

    \I__7165\ : InMux
    port map (
            O => \N__31330\,
            I => \N__31286\
        );

    \I__7164\ : InMux
    port map (
            O => \N__31329\,
            I => \N__31276\
        );

    \I__7163\ : InMux
    port map (
            O => \N__31328\,
            I => \N__31276\
        );

    \I__7162\ : InMux
    port map (
            O => \N__31327\,
            I => \N__31276\
        );

    \I__7161\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31276\
        );

    \I__7160\ : InMux
    port map (
            O => \N__31325\,
            I => \N__31271\
        );

    \I__7159\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31271\
        );

    \I__7158\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31262\
        );

    \I__7157\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31262\
        );

    \I__7156\ : InMux
    port map (
            O => \N__31321\,
            I => \N__31262\
        );

    \I__7155\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31262\
        );

    \I__7154\ : InMux
    port map (
            O => \N__31319\,
            I => \N__31253\
        );

    \I__7153\ : InMux
    port map (
            O => \N__31318\,
            I => \N__31253\
        );

    \I__7152\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31253\
        );

    \I__7151\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31253\
        );

    \I__7150\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31244\
        );

    \I__7149\ : InMux
    port map (
            O => \N__31314\,
            I => \N__31244\
        );

    \I__7148\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31241\
        );

    \I__7147\ : InMux
    port map (
            O => \N__31312\,
            I => \N__31232\
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__31311\,
            I => \N__31217\
        );

    \I__7145\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31203\
        );

    \I__7144\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31196\
        );

    \I__7143\ : InMux
    port map (
            O => \N__31308\,
            I => \N__31196\
        );

    \I__7142\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31196\
        );

    \I__7141\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31189\
        );

    \I__7140\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31189\
        );

    \I__7139\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31189\
        );

    \I__7138\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31182\
        );

    \I__7137\ : InMux
    port map (
            O => \N__31302\,
            I => \N__31182\
        );

    \I__7136\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31175\
        );

    \I__7135\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31175\
        );

    \I__7134\ : InMux
    port map (
            O => \N__31299\,
            I => \N__31175\
        );

    \I__7133\ : InMux
    port map (
            O => \N__31298\,
            I => \N__31168\
        );

    \I__7132\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31168\
        );

    \I__7131\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31156\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__31291\,
            I => \N__31151\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__31286\,
            I => \N__31151\
        );

    \I__7128\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31148\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__31276\,
            I => \N__31145\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__31271\,
            I => \N__31138\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__31262\,
            I => \N__31138\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__31253\,
            I => \N__31138\
        );

    \I__7123\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31131\
        );

    \I__7122\ : InMux
    port map (
            O => \N__31251\,
            I => \N__31131\
        );

    \I__7121\ : InMux
    port map (
            O => \N__31250\,
            I => \N__31131\
        );

    \I__7120\ : InMux
    port map (
            O => \N__31249\,
            I => \N__31127\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__31244\,
            I => \N__31122\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__31241\,
            I => \N__31122\
        );

    \I__7117\ : InMux
    port map (
            O => \N__31240\,
            I => \N__31113\
        );

    \I__7116\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31113\
        );

    \I__7115\ : InMux
    port map (
            O => \N__31238\,
            I => \N__31113\
        );

    \I__7114\ : InMux
    port map (
            O => \N__31237\,
            I => \N__31113\
        );

    \I__7113\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31105\
        );

    \I__7112\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31105\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__31232\,
            I => \N__31102\
        );

    \I__7110\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31097\
        );

    \I__7109\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31097\
        );

    \I__7108\ : InMux
    port map (
            O => \N__31229\,
            I => \N__31083\
        );

    \I__7107\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31080\
        );

    \I__7106\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31073\
        );

    \I__7105\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31073\
        );

    \I__7104\ : InMux
    port map (
            O => \N__31225\,
            I => \N__31073\
        );

    \I__7103\ : InMux
    port map (
            O => \N__31224\,
            I => \N__31065\
        );

    \I__7102\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31058\
        );

    \I__7101\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31058\
        );

    \I__7100\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31058\
        );

    \I__7099\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31051\
        );

    \I__7098\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31051\
        );

    \I__7097\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31051\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__31215\,
            I => \N__31045\
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__31214\,
            I => \N__31042\
        );

    \I__7094\ : InMux
    port map (
            O => \N__31213\,
            I => \N__31036\
        );

    \I__7093\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31036\
        );

    \I__7092\ : InMux
    port map (
            O => \N__31211\,
            I => \N__31031\
        );

    \I__7091\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31031\
        );

    \I__7090\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31022\
        );

    \I__7089\ : InMux
    port map (
            O => \N__31208\,
            I => \N__31022\
        );

    \I__7088\ : InMux
    port map (
            O => \N__31207\,
            I => \N__31022\
        );

    \I__7087\ : InMux
    port map (
            O => \N__31206\,
            I => \N__31022\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__31203\,
            I => \N__31019\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__31196\,
            I => \N__31016\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__31189\,
            I => \N__31013\
        );

    \I__7083\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31008\
        );

    \I__7082\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31008\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__31182\,
            I => \N__31003\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__31175\,
            I => \N__31003\
        );

    \I__7079\ : InMux
    port map (
            O => \N__31174\,
            I => \N__30998\
        );

    \I__7078\ : InMux
    port map (
            O => \N__31173\,
            I => \N__30998\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__30995\
        );

    \I__7076\ : InMux
    port map (
            O => \N__31167\,
            I => \N__30986\
        );

    \I__7075\ : InMux
    port map (
            O => \N__31166\,
            I => \N__30986\
        );

    \I__7074\ : InMux
    port map (
            O => \N__31165\,
            I => \N__30986\
        );

    \I__7073\ : InMux
    port map (
            O => \N__31164\,
            I => \N__30986\
        );

    \I__7072\ : InMux
    port map (
            O => \N__31163\,
            I => \N__30975\
        );

    \I__7071\ : InMux
    port map (
            O => \N__31162\,
            I => \N__30975\
        );

    \I__7070\ : InMux
    port map (
            O => \N__31161\,
            I => \N__30975\
        );

    \I__7069\ : InMux
    port map (
            O => \N__31160\,
            I => \N__30975\
        );

    \I__7068\ : InMux
    port map (
            O => \N__31159\,
            I => \N__30975\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__31156\,
            I => \N__30967\
        );

    \I__7066\ : Span4Mux_s3_v
    port map (
            O => \N__31151\,
            I => \N__30956\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__31148\,
            I => \N__30956\
        );

    \I__7064\ : Span4Mux_h
    port map (
            O => \N__31145\,
            I => \N__30956\
        );

    \I__7063\ : Span4Mux_h
    port map (
            O => \N__31138\,
            I => \N__30956\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__31131\,
            I => \N__30956\
        );

    \I__7061\ : InMux
    port map (
            O => \N__31130\,
            I => \N__30951\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__31127\,
            I => \N__30948\
        );

    \I__7059\ : Span4Mux_s3_h
    port map (
            O => \N__31122\,
            I => \N__30943\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__31113\,
            I => \N__30943\
        );

    \I__7057\ : InMux
    port map (
            O => \N__31112\,
            I => \N__30940\
        );

    \I__7056\ : CascadeMux
    port map (
            O => \N__31111\,
            I => \N__30934\
        );

    \I__7055\ : InMux
    port map (
            O => \N__31110\,
            I => \N__30931\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__31105\,
            I => \N__30926\
        );

    \I__7053\ : Span4Mux_v
    port map (
            O => \N__31102\,
            I => \N__30926\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__31097\,
            I => \N__30923\
        );

    \I__7051\ : InMux
    port map (
            O => \N__31096\,
            I => \N__30916\
        );

    \I__7050\ : InMux
    port map (
            O => \N__31095\,
            I => \N__30916\
        );

    \I__7049\ : InMux
    port map (
            O => \N__31094\,
            I => \N__30916\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31093\,
            I => \N__30913\
        );

    \I__7047\ : InMux
    port map (
            O => \N__31092\,
            I => \N__30908\
        );

    \I__7046\ : InMux
    port map (
            O => \N__31091\,
            I => \N__30908\
        );

    \I__7045\ : InMux
    port map (
            O => \N__31090\,
            I => \N__30901\
        );

    \I__7044\ : InMux
    port map (
            O => \N__31089\,
            I => \N__30901\
        );

    \I__7043\ : InMux
    port map (
            O => \N__31088\,
            I => \N__30898\
        );

    \I__7042\ : InMux
    port map (
            O => \N__31087\,
            I => \N__30893\
        );

    \I__7041\ : InMux
    port map (
            O => \N__31086\,
            I => \N__30893\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__31083\,
            I => \N__30886\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__31080\,
            I => \N__30886\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__30886\
        );

    \I__7037\ : InMux
    port map (
            O => \N__31072\,
            I => \N__30881\
        );

    \I__7036\ : InMux
    port map (
            O => \N__31071\,
            I => \N__30881\
        );

    \I__7035\ : InMux
    port map (
            O => \N__31070\,
            I => \N__30874\
        );

    \I__7034\ : InMux
    port map (
            O => \N__31069\,
            I => \N__30874\
        );

    \I__7033\ : InMux
    port map (
            O => \N__31068\,
            I => \N__30874\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__31065\,
            I => \N__30867\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__31058\,
            I => \N__30867\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__31051\,
            I => \N__30867\
        );

    \I__7029\ : InMux
    port map (
            O => \N__31050\,
            I => \N__30860\
        );

    \I__7028\ : InMux
    port map (
            O => \N__31049\,
            I => \N__30860\
        );

    \I__7027\ : InMux
    port map (
            O => \N__31048\,
            I => \N__30860\
        );

    \I__7026\ : InMux
    port map (
            O => \N__31045\,
            I => \N__30854\
        );

    \I__7025\ : InMux
    port map (
            O => \N__31042\,
            I => \N__30851\
        );

    \I__7024\ : InMux
    port map (
            O => \N__31041\,
            I => \N__30848\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__31036\,
            I => \N__30843\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__31031\,
            I => \N__30843\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__31022\,
            I => \N__30832\
        );

    \I__7020\ : Span4Mux_v
    port map (
            O => \N__31019\,
            I => \N__30832\
        );

    \I__7019\ : Span4Mux_v
    port map (
            O => \N__31016\,
            I => \N__30832\
        );

    \I__7018\ : Span4Mux_s1_h
    port map (
            O => \N__31013\,
            I => \N__30832\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__31008\,
            I => \N__30832\
        );

    \I__7016\ : Span4Mux_h
    port map (
            O => \N__31003\,
            I => \N__30821\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__30998\,
            I => \N__30821\
        );

    \I__7014\ : Span4Mux_v
    port map (
            O => \N__30995\,
            I => \N__30821\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__30986\,
            I => \N__30821\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__30975\,
            I => \N__30821\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__30974\,
            I => \N__30818\
        );

    \I__7010\ : InMux
    port map (
            O => \N__30973\,
            I => \N__30815\
        );

    \I__7009\ : InMux
    port map (
            O => \N__30972\,
            I => \N__30808\
        );

    \I__7008\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30808\
        );

    \I__7007\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30808\
        );

    \I__7006\ : Span4Mux_s3_v
    port map (
            O => \N__30967\,
            I => \N__30803\
        );

    \I__7005\ : Span4Mux_h
    port map (
            O => \N__30956\,
            I => \N__30803\
        );

    \I__7004\ : InMux
    port map (
            O => \N__30955\,
            I => \N__30798\
        );

    \I__7003\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30798\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__30951\,
            I => \N__30789\
        );

    \I__7001\ : Span4Mux_v
    port map (
            O => \N__30948\,
            I => \N__30789\
        );

    \I__7000\ : Span4Mux_h
    port map (
            O => \N__30943\,
            I => \N__30789\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__30940\,
            I => \N__30789\
        );

    \I__6998\ : InMux
    port map (
            O => \N__30939\,
            I => \N__30778\
        );

    \I__6997\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30778\
        );

    \I__6996\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30778\
        );

    \I__6995\ : InMux
    port map (
            O => \N__30934\,
            I => \N__30775\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__30931\,
            I => \N__30764\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__30926\,
            I => \N__30764\
        );

    \I__6992\ : Span4Mux_v
    port map (
            O => \N__30923\,
            I => \N__30764\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30764\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__30913\,
            I => \N__30764\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__30908\,
            I => \N__30761\
        );

    \I__6988\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30756\
        );

    \I__6987\ : InMux
    port map (
            O => \N__30906\,
            I => \N__30756\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__30901\,
            I => \N__30747\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__30898\,
            I => \N__30747\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__30893\,
            I => \N__30747\
        );

    \I__6983\ : Span4Mux_v
    port map (
            O => \N__30886\,
            I => \N__30747\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__30881\,
            I => \N__30738\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__30874\,
            I => \N__30738\
        );

    \I__6980\ : Span4Mux_v
    port map (
            O => \N__30867\,
            I => \N__30738\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__30860\,
            I => \N__30738\
        );

    \I__6978\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30733\
        );

    \I__6977\ : InMux
    port map (
            O => \N__30858\,
            I => \N__30733\
        );

    \I__6976\ : CascadeMux
    port map (
            O => \N__30857\,
            I => \N__30730\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__30854\,
            I => \N__30722\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__30851\,
            I => \N__30722\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__30848\,
            I => \N__30711\
        );

    \I__6972\ : Span4Mux_v
    port map (
            O => \N__30843\,
            I => \N__30704\
        );

    \I__6971\ : Span4Mux_h
    port map (
            O => \N__30832\,
            I => \N__30704\
        );

    \I__6970\ : Span4Mux_v
    port map (
            O => \N__30821\,
            I => \N__30704\
        );

    \I__6969\ : InMux
    port map (
            O => \N__30818\,
            I => \N__30701\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__30815\,
            I => \N__30694\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__30808\,
            I => \N__30694\
        );

    \I__6966\ : Span4Mux_v
    port map (
            O => \N__30803\,
            I => \N__30694\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__30798\,
            I => \N__30689\
        );

    \I__6964\ : Span4Mux_v
    port map (
            O => \N__30789\,
            I => \N__30689\
        );

    \I__6963\ : InMux
    port map (
            O => \N__30788\,
            I => \N__30682\
        );

    \I__6962\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30682\
        );

    \I__6961\ : InMux
    port map (
            O => \N__30786\,
            I => \N__30682\
        );

    \I__6960\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30679\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30676\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__30775\,
            I => \N__30673\
        );

    \I__6957\ : Span4Mux_h
    port map (
            O => \N__30764\,
            I => \N__30668\
        );

    \I__6956\ : Span4Mux_s3_h
    port map (
            O => \N__30761\,
            I => \N__30668\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30659\
        );

    \I__6954\ : Span4Mux_h
    port map (
            O => \N__30747\,
            I => \N__30659\
        );

    \I__6953\ : Span4Mux_v
    port map (
            O => \N__30738\,
            I => \N__30659\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__30733\,
            I => \N__30659\
        );

    \I__6951\ : InMux
    port map (
            O => \N__30730\,
            I => \N__30656\
        );

    \I__6950\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30649\
        );

    \I__6949\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30649\
        );

    \I__6948\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30649\
        );

    \I__6947\ : Span4Mux_s3_h
    port map (
            O => \N__30722\,
            I => \N__30646\
        );

    \I__6946\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30641\
        );

    \I__6945\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30641\
        );

    \I__6944\ : InMux
    port map (
            O => \N__30719\,
            I => \N__30636\
        );

    \I__6943\ : InMux
    port map (
            O => \N__30718\,
            I => \N__30636\
        );

    \I__6942\ : InMux
    port map (
            O => \N__30717\,
            I => \N__30629\
        );

    \I__6941\ : InMux
    port map (
            O => \N__30716\,
            I => \N__30629\
        );

    \I__6940\ : InMux
    port map (
            O => \N__30715\,
            I => \N__30629\
        );

    \I__6939\ : InMux
    port map (
            O => \N__30714\,
            I => \N__30626\
        );

    \I__6938\ : Span4Mux_v
    port map (
            O => \N__30711\,
            I => \N__30621\
        );

    \I__6937\ : Span4Mux_h
    port map (
            O => \N__30704\,
            I => \N__30621\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__30701\,
            I => \N__30614\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__30694\,
            I => \N__30614\
        );

    \I__6934\ : Span4Mux_h
    port map (
            O => \N__30689\,
            I => \N__30614\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__30682\,
            I => \N__30607\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__30679\,
            I => \N__30607\
        );

    \I__6931\ : Span12Mux_s11_v
    port map (
            O => \N__30676\,
            I => \N__30607\
        );

    \I__6930\ : Span4Mux_v
    port map (
            O => \N__30673\,
            I => \N__30598\
        );

    \I__6929\ : Span4Mux_v
    port map (
            O => \N__30668\,
            I => \N__30598\
        );

    \I__6928\ : Span4Mux_h
    port map (
            O => \N__30659\,
            I => \N__30598\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__30656\,
            I => \N__30598\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__30649\,
            I => \tok.T_0\
        );

    \I__6925\ : Odrv4
    port map (
            O => \N__30646\,
            I => \tok.T_0\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__30641\,
            I => \tok.T_0\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__30636\,
            I => \tok.T_0\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__30629\,
            I => \tok.T_0\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__30626\,
            I => \tok.T_0\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__30621\,
            I => \tok.T_0\
        );

    \I__6919\ : Odrv4
    port map (
            O => \N__30614\,
            I => \tok.T_0\
        );

    \I__6918\ : Odrv12
    port map (
            O => \N__30607\,
            I => \tok.T_0\
        );

    \I__6917\ : Odrv4
    port map (
            O => \N__30598\,
            I => \tok.T_0\
        );

    \I__6916\ : CascadeMux
    port map (
            O => \N__30577\,
            I => \N__30574\
        );

    \I__6915\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30571\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__30571\,
            I => \tok.n168_adj_690\
        );

    \I__6913\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30565\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__30565\,
            I => \N__30562\
        );

    \I__6911\ : Span4Mux_s3_h
    port map (
            O => \N__30562\,
            I => \N__30559\
        );

    \I__6910\ : Span4Mux_h
    port map (
            O => \N__30559\,
            I => \N__30556\
        );

    \I__6909\ : Odrv4
    port map (
            O => \N__30556\,
            I => \tok.n6525\
        );

    \I__6908\ : CascadeMux
    port map (
            O => \N__30553\,
            I => \tok.n6526_cascade_\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__30550\,
            I => \tok.n186_adj_777_cascade_\
        );

    \I__6906\ : CascadeMux
    port map (
            O => \N__30547\,
            I => \N__30544\
        );

    \I__6905\ : InMux
    port map (
            O => \N__30544\,
            I => \N__30541\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__30541\,
            I => \N__30538\
        );

    \I__6903\ : Odrv12
    port map (
            O => \N__30538\,
            I => \tok.n338_adj_787\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__30535\,
            I => \N__30528\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__30534\,
            I => \N__30521\
        );

    \I__6900\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30518\
        );

    \I__6899\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30515\
        );

    \I__6898\ : InMux
    port map (
            O => \N__30531\,
            I => \N__30512\
        );

    \I__6897\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30504\
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__30527\,
            I => \N__30500\
        );

    \I__6895\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30496\
        );

    \I__6894\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30493\
        );

    \I__6893\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30488\
        );

    \I__6892\ : InMux
    port map (
            O => \N__30521\,
            I => \N__30488\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__30518\,
            I => \N__30482\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__30515\,
            I => \N__30482\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__30512\,
            I => \N__30479\
        );

    \I__6888\ : InMux
    port map (
            O => \N__30511\,
            I => \N__30475\
        );

    \I__6887\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30470\
        );

    \I__6886\ : InMux
    port map (
            O => \N__30509\,
            I => \N__30470\
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__30508\,
            I => \N__30467\
        );

    \I__6884\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30464\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__30504\,
            I => \N__30461\
        );

    \I__6882\ : InMux
    port map (
            O => \N__30503\,
            I => \N__30458\
        );

    \I__6881\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30455\
        );

    \I__6880\ : CascadeMux
    port map (
            O => \N__30499\,
            I => \N__30452\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__30496\,
            I => \N__30449\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__30493\,
            I => \N__30446\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__30488\,
            I => \N__30443\
        );

    \I__6876\ : InMux
    port map (
            O => \N__30487\,
            I => \N__30440\
        );

    \I__6875\ : Span4Mux_s3_v
    port map (
            O => \N__30482\,
            I => \N__30435\
        );

    \I__6874\ : Span4Mux_h
    port map (
            O => \N__30479\,
            I => \N__30435\
        );

    \I__6873\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30432\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__30475\,
            I => \N__30429\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__30470\,
            I => \N__30426\
        );

    \I__6870\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30423\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__30464\,
            I => \N__30414\
        );

    \I__6868\ : Span4Mux_v
    port map (
            O => \N__30461\,
            I => \N__30414\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__30458\,
            I => \N__30414\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__30455\,
            I => \N__30414\
        );

    \I__6865\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30411\
        );

    \I__6864\ : Span4Mux_v
    port map (
            O => \N__30449\,
            I => \N__30407\
        );

    \I__6863\ : Span4Mux_v
    port map (
            O => \N__30446\,
            I => \N__30404\
        );

    \I__6862\ : Span4Mux_s3_v
    port map (
            O => \N__30443\,
            I => \N__30395\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__30440\,
            I => \N__30395\
        );

    \I__6860\ : Span4Mux_h
    port map (
            O => \N__30435\,
            I => \N__30395\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__30432\,
            I => \N__30395\
        );

    \I__6858\ : Span4Mux_v
    port map (
            O => \N__30429\,
            I => \N__30382\
        );

    \I__6857\ : Span4Mux_v
    port map (
            O => \N__30426\,
            I => \N__30382\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__30423\,
            I => \N__30382\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__30414\,
            I => \N__30382\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__30411\,
            I => \N__30379\
        );

    \I__6853\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30376\
        );

    \I__6852\ : Span4Mux_h
    port map (
            O => \N__30407\,
            I => \N__30369\
        );

    \I__6851\ : Span4Mux_h
    port map (
            O => \N__30404\,
            I => \N__30369\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__30395\,
            I => \N__30369\
        );

    \I__6849\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30360\
        );

    \I__6848\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30360\
        );

    \I__6847\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30360\
        );

    \I__6846\ : InMux
    port map (
            O => \N__30391\,
            I => \N__30360\
        );

    \I__6845\ : Span4Mux_h
    port map (
            O => \N__30382\,
            I => \N__30357\
        );

    \I__6844\ : Odrv12
    port map (
            O => \N__30379\,
            I => \tok.A_low_0\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__30376\,
            I => \tok.A_low_0\
        );

    \I__6842\ : Odrv4
    port map (
            O => \N__30369\,
            I => \tok.A_low_0\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__30360\,
            I => \tok.A_low_0\
        );

    \I__6840\ : Odrv4
    port map (
            O => \N__30357\,
            I => \tok.A_low_0\
        );

    \I__6839\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30339\
        );

    \I__6838\ : CascadeMux
    port map (
            O => \N__30345\,
            I => \N__30336\
        );

    \I__6837\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30333\
        );

    \I__6836\ : InMux
    port map (
            O => \N__30343\,
            I => \N__30330\
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__30342\,
            I => \N__30315\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__30339\,
            I => \N__30309\
        );

    \I__6833\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30306\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__30333\,
            I => \N__30303\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__30330\,
            I => \N__30300\
        );

    \I__6830\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30293\
        );

    \I__6829\ : InMux
    port map (
            O => \N__30328\,
            I => \N__30293\
        );

    \I__6828\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30293\
        );

    \I__6827\ : InMux
    port map (
            O => \N__30326\,
            I => \N__30286\
        );

    \I__6826\ : InMux
    port map (
            O => \N__30325\,
            I => \N__30286\
        );

    \I__6825\ : InMux
    port map (
            O => \N__30324\,
            I => \N__30286\
        );

    \I__6824\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30283\
        );

    \I__6823\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30280\
        );

    \I__6822\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30277\
        );

    \I__6821\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30274\
        );

    \I__6820\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30271\
        );

    \I__6819\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30268\
        );

    \I__6818\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30265\
        );

    \I__6817\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30260\
        );

    \I__6816\ : InMux
    port map (
            O => \N__30313\,
            I => \N__30260\
        );

    \I__6815\ : CascadeMux
    port map (
            O => \N__30312\,
            I => \N__30255\
        );

    \I__6814\ : Span4Mux_s2_h
    port map (
            O => \N__30309\,
            I => \N__30250\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__30306\,
            I => \N__30250\
        );

    \I__6812\ : Span4Mux_s3_h
    port map (
            O => \N__30303\,
            I => \N__30247\
        );

    \I__6811\ : Span4Mux_s3_h
    port map (
            O => \N__30300\,
            I => \N__30240\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__30293\,
            I => \N__30240\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__30286\,
            I => \N__30240\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__30283\,
            I => \N__30237\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__30280\,
            I => \N__30232\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__30277\,
            I => \N__30232\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__30274\,
            I => \N__30227\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__30271\,
            I => \N__30227\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__30268\,
            I => \N__30222\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__30265\,
            I => \N__30222\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__30260\,
            I => \N__30219\
        );

    \I__6800\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30214\
        );

    \I__6799\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30214\
        );

    \I__6798\ : InMux
    port map (
            O => \N__30255\,
            I => \N__30211\
        );

    \I__6797\ : Span4Mux_h
    port map (
            O => \N__30250\,
            I => \N__30206\
        );

    \I__6796\ : Span4Mux_h
    port map (
            O => \N__30247\,
            I => \N__30206\
        );

    \I__6795\ : Span4Mux_h
    port map (
            O => \N__30240\,
            I => \N__30203\
        );

    \I__6794\ : Span4Mux_v
    port map (
            O => \N__30237\,
            I => \N__30194\
        );

    \I__6793\ : Span4Mux_h
    port map (
            O => \N__30232\,
            I => \N__30194\
        );

    \I__6792\ : Span4Mux_v
    port map (
            O => \N__30227\,
            I => \N__30194\
        );

    \I__6791\ : Span4Mux_v
    port map (
            O => \N__30222\,
            I => \N__30194\
        );

    \I__6790\ : Odrv12
    port map (
            O => \N__30219\,
            I => \tok.A_low_5\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__30214\,
            I => \tok.A_low_5\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__30211\,
            I => \tok.A_low_5\
        );

    \I__6787\ : Odrv4
    port map (
            O => \N__30206\,
            I => \tok.A_low_5\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__30203\,
            I => \tok.A_low_5\
        );

    \I__6785\ : Odrv4
    port map (
            O => \N__30194\,
            I => \tok.A_low_5\
        );

    \I__6784\ : CascadeMux
    port map (
            O => \N__30181\,
            I => \tok.n866_cascade_\
        );

    \I__6783\ : InMux
    port map (
            O => \N__30178\,
            I => \N__30175\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__30175\,
            I => \tok.n6520\
        );

    \I__6781\ : CascadeMux
    port map (
            O => \N__30172\,
            I => \tok.n10_cascade_\
        );

    \I__6780\ : SRMux
    port map (
            O => \N__30169\,
            I => \N__30166\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__30166\,
            I => \N__30163\
        );

    \I__6778\ : Span4Mux_h
    port map (
            O => \N__30163\,
            I => \N__30160\
        );

    \I__6777\ : Span4Mux_h
    port map (
            O => \N__30160\,
            I => \N__30157\
        );

    \I__6776\ : Span4Mux_s2_v
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__6775\ : Span4Mux_v
    port map (
            O => \N__30154\,
            I => \N__30151\
        );

    \I__6774\ : Odrv4
    port map (
            O => \N__30151\,
            I => \tok.write_flag\
        );

    \I__6773\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30135\
        );

    \I__6772\ : InMux
    port map (
            O => \N__30147\,
            I => \N__30135\
        );

    \I__6771\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30135\
        );

    \I__6770\ : InMux
    port map (
            O => \N__30145\,
            I => \N__30131\
        );

    \I__6769\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30124\
        );

    \I__6768\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30124\
        );

    \I__6767\ : InMux
    port map (
            O => \N__30142\,
            I => \N__30124\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__30135\,
            I => \N__30121\
        );

    \I__6765\ : InMux
    port map (
            O => \N__30134\,
            I => \N__30118\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__30131\,
            I => \N__30113\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__30124\,
            I => \N__30113\
        );

    \I__6762\ : Span4Mux_v
    port map (
            O => \N__30121\,
            I => \N__30110\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__30118\,
            I => \N__30105\
        );

    \I__6760\ : Span4Mux_h
    port map (
            O => \N__30113\,
            I => \N__30105\
        );

    \I__6759\ : Sp12to4
    port map (
            O => \N__30110\,
            I => \N__30102\
        );

    \I__6758\ : Span4Mux_v
    port map (
            O => \N__30105\,
            I => \N__30099\
        );

    \I__6757\ : Odrv12
    port map (
            O => \N__30102\,
            I => \tok.n14\
        );

    \I__6756\ : Odrv4
    port map (
            O => \N__30099\,
            I => \tok.n14\
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__30094\,
            I => \tok.uart.n10_cascade_\
        );

    \I__6754\ : CascadeMux
    port map (
            O => \N__30091\,
            I => \n23_cascade_\
        );

    \I__6753\ : CascadeMux
    port map (
            O => \N__30088\,
            I => \tok.n168_adj_710_cascade_\
        );

    \I__6752\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30080\
        );

    \I__6751\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30075\
        );

    \I__6750\ : InMux
    port map (
            O => \N__30083\,
            I => \N__30075\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__30080\,
            I => \N__30067\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__30075\,
            I => \N__30067\
        );

    \I__6747\ : CascadeMux
    port map (
            O => \N__30074\,
            I => \N__30059\
        );

    \I__6746\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30055\
        );

    \I__6745\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30050\
        );

    \I__6744\ : Span4Mux_h
    port map (
            O => \N__30067\,
            I => \N__30047\
        );

    \I__6743\ : CascadeMux
    port map (
            O => \N__30066\,
            I => \N__30044\
        );

    \I__6742\ : CascadeMux
    port map (
            O => \N__30065\,
            I => \N__30039\
        );

    \I__6741\ : InMux
    port map (
            O => \N__30064\,
            I => \N__30035\
        );

    \I__6740\ : InMux
    port map (
            O => \N__30063\,
            I => \N__30032\
        );

    \I__6739\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30029\
        );

    \I__6738\ : InMux
    port map (
            O => \N__30059\,
            I => \N__30023\
        );

    \I__6737\ : InMux
    port map (
            O => \N__30058\,
            I => \N__30020\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__30055\,
            I => \N__30017\
        );

    \I__6735\ : InMux
    port map (
            O => \N__30054\,
            I => \N__30014\
        );

    \I__6734\ : CascadeMux
    port map (
            O => \N__30053\,
            I => \N__30011\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__30050\,
            I => \N__30005\
        );

    \I__6732\ : IoSpan4Mux
    port map (
            O => \N__30047\,
            I => \N__30005\
        );

    \I__6731\ : InMux
    port map (
            O => \N__30044\,
            I => \N__30000\
        );

    \I__6730\ : InMux
    port map (
            O => \N__30043\,
            I => \N__30000\
        );

    \I__6729\ : InMux
    port map (
            O => \N__30042\,
            I => \N__29997\
        );

    \I__6728\ : InMux
    port map (
            O => \N__30039\,
            I => \N__29994\
        );

    \I__6727\ : InMux
    port map (
            O => \N__30038\,
            I => \N__29991\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__30035\,
            I => \N__29988\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__30032\,
            I => \N__29985\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__30029\,
            I => \N__29982\
        );

    \I__6723\ : InMux
    port map (
            O => \N__30028\,
            I => \N__29977\
        );

    \I__6722\ : InMux
    port map (
            O => \N__30027\,
            I => \N__29977\
        );

    \I__6721\ : InMux
    port map (
            O => \N__30026\,
            I => \N__29974\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__30023\,
            I => \N__29971\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__30020\,
            I => \N__29968\
        );

    \I__6718\ : Span4Mux_s3_v
    port map (
            O => \N__30017\,
            I => \N__29963\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__30014\,
            I => \N__29963\
        );

    \I__6716\ : InMux
    port map (
            O => \N__30011\,
            I => \N__29960\
        );

    \I__6715\ : InMux
    port map (
            O => \N__30010\,
            I => \N__29957\
        );

    \I__6714\ : Span4Mux_s2_v
    port map (
            O => \N__30005\,
            I => \N__29948\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__30000\,
            I => \N__29948\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__29997\,
            I => \N__29948\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__29994\,
            I => \N__29948\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__29991\,
            I => \N__29945\
        );

    \I__6709\ : Span4Mux_v
    port map (
            O => \N__29988\,
            I => \N__29942\
        );

    \I__6708\ : Span4Mux_v
    port map (
            O => \N__29985\,
            I => \N__29939\
        );

    \I__6707\ : Span4Mux_v
    port map (
            O => \N__29982\,
            I => \N__29932\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__29977\,
            I => \N__29932\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__29974\,
            I => \N__29932\
        );

    \I__6704\ : Span4Mux_s2_v
    port map (
            O => \N__29971\,
            I => \N__29926\
        );

    \I__6703\ : Span4Mux_h
    port map (
            O => \N__29968\,
            I => \N__29926\
        );

    \I__6702\ : Span4Mux_v
    port map (
            O => \N__29963\,
            I => \N__29917\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__29960\,
            I => \N__29917\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__29957\,
            I => \N__29917\
        );

    \I__6699\ : Span4Mux_v
    port map (
            O => \N__29948\,
            I => \N__29917\
        );

    \I__6698\ : Span12Mux_s8_v
    port map (
            O => \N__29945\,
            I => \N__29912\
        );

    \I__6697\ : Sp12to4
    port map (
            O => \N__29942\,
            I => \N__29912\
        );

    \I__6696\ : Span4Mux_v
    port map (
            O => \N__29939\,
            I => \N__29907\
        );

    \I__6695\ : Span4Mux_v
    port map (
            O => \N__29932\,
            I => \N__29907\
        );

    \I__6694\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29904\
        );

    \I__6693\ : Span4Mux_v
    port map (
            O => \N__29926\,
            I => \N__29899\
        );

    \I__6692\ : Span4Mux_h
    port map (
            O => \N__29917\,
            I => \N__29899\
        );

    \I__6691\ : Odrv12
    port map (
            O => \N__29912\,
            I => \tok.A_low_6\
        );

    \I__6690\ : Odrv4
    port map (
            O => \N__29907\,
            I => \tok.A_low_6\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__29904\,
            I => \tok.A_low_6\
        );

    \I__6688\ : Odrv4
    port map (
            O => \N__29899\,
            I => \tok.A_low_6\
        );

    \I__6687\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29887\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__29887\,
            I => \tok.n6502\
        );

    \I__6685\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29878\
        );

    \I__6684\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29878\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__29878\,
            I => uart_rx_data_6
        );

    \I__6682\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29865\
        );

    \I__6681\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29865\
        );

    \I__6680\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29856\
        );

    \I__6679\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29856\
        );

    \I__6678\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29856\
        );

    \I__6677\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29856\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__29865\,
            I => \tok.depth_1\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__29856\,
            I => \tok.depth_1\
        );

    \I__6674\ : CascadeMux
    port map (
            O => \N__29851\,
            I => \N__29848\
        );

    \I__6673\ : InMux
    port map (
            O => \N__29848\,
            I => \N__29842\
        );

    \I__6672\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29842\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__29842\,
            I => \tok.n741\
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__29839\,
            I => \N__29835\
        );

    \I__6669\ : CascadeMux
    port map (
            O => \N__29838\,
            I => \N__29832\
        );

    \I__6668\ : InMux
    port map (
            O => \N__29835\,
            I => \N__29827\
        );

    \I__6667\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29827\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__29827\,
            I => \N__29824\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__29824\,
            I => \N__29821\
        );

    \I__6664\ : Odrv4
    port map (
            O => \N__29821\,
            I => \tok.n806\
        );

    \I__6663\ : CascadeMux
    port map (
            O => \N__29818\,
            I => \N__29815\
        );

    \I__6662\ : InMux
    port map (
            O => \N__29815\,
            I => \N__29806\
        );

    \I__6661\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29806\
        );

    \I__6660\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29803\
        );

    \I__6659\ : CascadeMux
    port map (
            O => \N__29812\,
            I => \N__29799\
        );

    \I__6658\ : CascadeMux
    port map (
            O => \N__29811\,
            I => \N__29795\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__29806\,
            I => \N__29789\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__29803\,
            I => \N__29789\
        );

    \I__6655\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29784\
        );

    \I__6654\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29784\
        );

    \I__6653\ : InMux
    port map (
            O => \N__29798\,
            I => \N__29777\
        );

    \I__6652\ : InMux
    port map (
            O => \N__29795\,
            I => \N__29777\
        );

    \I__6651\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29777\
        );

    \I__6650\ : Odrv4
    port map (
            O => \N__29789\,
            I => \tok.depth_0\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__29784\,
            I => \tok.depth_0\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__29777\,
            I => \tok.depth_0\
        );

    \I__6647\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29767\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__29767\,
            I => \tok.n6213\
        );

    \I__6645\ : CascadeMux
    port map (
            O => \N__29764\,
            I => \tok.n806_cascade_\
        );

    \I__6644\ : CascadeMux
    port map (
            O => \N__29761\,
            I => \N__29754\
        );

    \I__6643\ : CascadeMux
    port map (
            O => \N__29760\,
            I => \N__29750\
        );

    \I__6642\ : InMux
    port map (
            O => \N__29759\,
            I => \N__29747\
        );

    \I__6641\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29744\
        );

    \I__6640\ : InMux
    port map (
            O => \N__29757\,
            I => \N__29741\
        );

    \I__6639\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29734\
        );

    \I__6638\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29734\
        );

    \I__6637\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29734\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__29747\,
            I => \tok.depth_3\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__29744\,
            I => \tok.depth_3\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__29741\,
            I => \tok.depth_3\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__29734\,
            I => \tok.depth_3\
        );

    \I__6632\ : CascadeMux
    port map (
            O => \N__29725\,
            I => \N__29720\
        );

    \I__6631\ : CascadeMux
    port map (
            O => \N__29724\,
            I => \N__29715\
        );

    \I__6630\ : CascadeMux
    port map (
            O => \N__29723\,
            I => \N__29712\
        );

    \I__6629\ : InMux
    port map (
            O => \N__29720\,
            I => \N__29707\
        );

    \I__6628\ : InMux
    port map (
            O => \N__29719\,
            I => \N__29703\
        );

    \I__6627\ : InMux
    port map (
            O => \N__29718\,
            I => \N__29700\
        );

    \I__6626\ : InMux
    port map (
            O => \N__29715\,
            I => \N__29697\
        );

    \I__6625\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29694\
        );

    \I__6624\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29691\
        );

    \I__6623\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29688\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__29707\,
            I => \N__29685\
        );

    \I__6621\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29682\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__29703\,
            I => \N__29677\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__29700\,
            I => \N__29677\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__29697\,
            I => \N__29674\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__29694\,
            I => \N__29671\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__29691\,
            I => \N__29668\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__29688\,
            I => \N__29661\
        );

    \I__6614\ : Span4Mux_h
    port map (
            O => \N__29685\,
            I => \N__29661\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__29682\,
            I => \N__29661\
        );

    \I__6612\ : Span4Mux_v
    port map (
            O => \N__29677\,
            I => \N__29658\
        );

    \I__6611\ : Span4Mux_v
    port map (
            O => \N__29674\,
            I => \N__29653\
        );

    \I__6610\ : Span4Mux_v
    port map (
            O => \N__29671\,
            I => \N__29653\
        );

    \I__6609\ : Span4Mux_h
    port map (
            O => \N__29668\,
            I => \N__29650\
        );

    \I__6608\ : Span4Mux_h
    port map (
            O => \N__29661\,
            I => \N__29647\
        );

    \I__6607\ : Span4Mux_h
    port map (
            O => \N__29658\,
            I => \N__29644\
        );

    \I__6606\ : Span4Mux_h
    port map (
            O => \N__29653\,
            I => \N__29641\
        );

    \I__6605\ : Span4Mux_v
    port map (
            O => \N__29650\,
            I => \N__29634\
        );

    \I__6604\ : Span4Mux_v
    port map (
            O => \N__29647\,
            I => \N__29634\
        );

    \I__6603\ : Span4Mux_h
    port map (
            O => \N__29644\,
            I => \N__29634\
        );

    \I__6602\ : Odrv4
    port map (
            O => \N__29641\,
            I => \tok.n748\
        );

    \I__6601\ : Odrv4
    port map (
            O => \N__29634\,
            I => \tok.n748\
        );

    \I__6600\ : InMux
    port map (
            O => \N__29629\,
            I => \N__29623\
        );

    \I__6599\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29614\
        );

    \I__6598\ : InMux
    port map (
            O => \N__29627\,
            I => \N__29611\
        );

    \I__6597\ : InMux
    port map (
            O => \N__29626\,
            I => \N__29608\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__29623\,
            I => \N__29605\
        );

    \I__6595\ : InMux
    port map (
            O => \N__29622\,
            I => \N__29600\
        );

    \I__6594\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29600\
        );

    \I__6593\ : InMux
    port map (
            O => \N__29620\,
            I => \N__29597\
        );

    \I__6592\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29592\
        );

    \I__6591\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29587\
        );

    \I__6590\ : InMux
    port map (
            O => \N__29617\,
            I => \N__29587\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__29614\,
            I => \N__29584\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__29611\,
            I => \N__29581\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__29608\,
            I => \N__29578\
        );

    \I__6586\ : Span4Mux_v
    port map (
            O => \N__29605\,
            I => \N__29572\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__29600\,
            I => \N__29572\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__29597\,
            I => \N__29569\
        );

    \I__6583\ : CascadeMux
    port map (
            O => \N__29596\,
            I => \N__29566\
        );

    \I__6582\ : InMux
    port map (
            O => \N__29595\,
            I => \N__29563\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__29592\,
            I => \N__29559\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__29587\,
            I => \N__29556\
        );

    \I__6579\ : Span4Mux_h
    port map (
            O => \N__29584\,
            I => \N__29553\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__29581\,
            I => \N__29550\
        );

    \I__6577\ : Span4Mux_v
    port map (
            O => \N__29578\,
            I => \N__29544\
        );

    \I__6576\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29541\
        );

    \I__6575\ : Span4Mux_v
    port map (
            O => \N__29572\,
            I => \N__29536\
        );

    \I__6574\ : Span4Mux_s3_h
    port map (
            O => \N__29569\,
            I => \N__29536\
        );

    \I__6573\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29533\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__29563\,
            I => \N__29530\
        );

    \I__6571\ : CascadeMux
    port map (
            O => \N__29562\,
            I => \N__29526\
        );

    \I__6570\ : Span4Mux_v
    port map (
            O => \N__29559\,
            I => \N__29521\
        );

    \I__6569\ : Span4Mux_v
    port map (
            O => \N__29556\,
            I => \N__29521\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__29553\,
            I => \N__29516\
        );

    \I__6567\ : Span4Mux_h
    port map (
            O => \N__29550\,
            I => \N__29516\
        );

    \I__6566\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29509\
        );

    \I__6565\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29509\
        );

    \I__6564\ : InMux
    port map (
            O => \N__29547\,
            I => \N__29509\
        );

    \I__6563\ : Span4Mux_h
    port map (
            O => \N__29544\,
            I => \N__29504\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29504\
        );

    \I__6561\ : Span4Mux_h
    port map (
            O => \N__29536\,
            I => \N__29501\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__29533\,
            I => \N__29496\
        );

    \I__6559\ : Span12Mux_s7_h
    port map (
            O => \N__29530\,
            I => \N__29496\
        );

    \I__6558\ : InMux
    port map (
            O => \N__29529\,
            I => \N__29491\
        );

    \I__6557\ : InMux
    port map (
            O => \N__29526\,
            I => \N__29491\
        );

    \I__6556\ : Odrv4
    port map (
            O => \N__29521\,
            I => \tok.n47\
        );

    \I__6555\ : Odrv4
    port map (
            O => \N__29516\,
            I => \tok.n47\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__29509\,
            I => \tok.n47\
        );

    \I__6553\ : Odrv4
    port map (
            O => \N__29504\,
            I => \tok.n47\
        );

    \I__6552\ : Odrv4
    port map (
            O => \N__29501\,
            I => \tok.n47\
        );

    \I__6551\ : Odrv12
    port map (
            O => \N__29496\,
            I => \tok.n47\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__29491\,
            I => \tok.n47\
        );

    \I__6549\ : CascadeMux
    port map (
            O => \N__29476\,
            I => \N__29473\
        );

    \I__6548\ : InMux
    port map (
            O => \N__29473\,
            I => \N__29470\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__29470\,
            I => \N__29467\
        );

    \I__6546\ : Span12Mux_s9_h
    port map (
            O => \N__29467\,
            I => \N__29464\
        );

    \I__6545\ : Odrv12
    port map (
            O => \N__29464\,
            I => \tok.n6615\
        );

    \I__6544\ : CascadeMux
    port map (
            O => \N__29461\,
            I => \tok.n158_cascade_\
        );

    \I__6543\ : InMux
    port map (
            O => \N__29458\,
            I => \N__29455\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__29455\,
            I => \N__29452\
        );

    \I__6541\ : Odrv4
    port map (
            O => \N__29452\,
            I => \tok.n6627\
        );

    \I__6540\ : InMux
    port map (
            O => \N__29449\,
            I => \N__29440\
        );

    \I__6539\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29440\
        );

    \I__6538\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29440\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29437\
        );

    \I__6536\ : Span4Mux_h
    port map (
            O => \N__29437\,
            I => \N__29434\
        );

    \I__6535\ : Span4Mux_h
    port map (
            O => \N__29434\,
            I => \N__29431\
        );

    \I__6534\ : Odrv4
    port map (
            O => \N__29431\,
            I => \tok.uart_stall_N_46\
        );

    \I__6533\ : InMux
    port map (
            O => \N__29428\,
            I => \N__29425\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__29425\,
            I => \tok.n9\
        );

    \I__6531\ : CascadeMux
    port map (
            O => \N__29422\,
            I => \N__29419\
        );

    \I__6530\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29416\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__29416\,
            I => \tok.n10\
        );

    \I__6528\ : InMux
    port map (
            O => \N__29413\,
            I => \N__29409\
        );

    \I__6527\ : CascadeMux
    port map (
            O => \N__29412\,
            I => \N__29405\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__29409\,
            I => \N__29402\
        );

    \I__6525\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29397\
        );

    \I__6524\ : InMux
    port map (
            O => \N__29405\,
            I => \N__29392\
        );

    \I__6523\ : Span12Mux_h
    port map (
            O => \N__29402\,
            I => \N__29389\
        );

    \I__6522\ : InMux
    port map (
            O => \N__29401\,
            I => \N__29384\
        );

    \I__6521\ : InMux
    port map (
            O => \N__29400\,
            I => \N__29384\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__29397\,
            I => \N__29381\
        );

    \I__6519\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29376\
        );

    \I__6518\ : InMux
    port map (
            O => \N__29395\,
            I => \N__29376\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__29392\,
            I => \N__29373\
        );

    \I__6516\ : Odrv12
    port map (
            O => \N__29389\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__29384\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__29381\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__29376\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__29373\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__6511\ : CascadeMux
    port map (
            O => \N__29362\,
            I => \tok.A_stk_delta_1__N_4_cascade_\
        );

    \I__6510\ : CascadeMux
    port map (
            O => \N__29359\,
            I => \N__29356\
        );

    \I__6509\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29347\
        );

    \I__6508\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29347\
        );

    \I__6507\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29347\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__29347\,
            I => \N__29341\
        );

    \I__6505\ : InMux
    port map (
            O => \N__29346\,
            I => \N__29334\
        );

    \I__6504\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29334\
        );

    \I__6503\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29334\
        );

    \I__6502\ : Span4Mux_s1_h
    port map (
            O => \N__29341\,
            I => \N__29331\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__29334\,
            I => \N__29328\
        );

    \I__6500\ : Odrv4
    port map (
            O => \N__29331\,
            I => \tok.n1\
        );

    \I__6499\ : Odrv12
    port map (
            O => \N__29328\,
            I => \tok.n1\
        );

    \I__6498\ : CascadeMux
    port map (
            O => \N__29323\,
            I => \tok.n4_adj_702_cascade_\
        );

    \I__6497\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29317\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__29317\,
            I => \tok.n52\
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__29314\,
            I => \tok.n51_cascade_\
        );

    \I__6494\ : InMux
    port map (
            O => \N__29311\,
            I => \N__29308\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__29308\,
            I => \tok.n50\
        );

    \I__6492\ : InMux
    port map (
            O => \N__29305\,
            I => \N__29302\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__29302\,
            I => \tok.n8_adj_854\
        );

    \I__6490\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29290\
        );

    \I__6489\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29290\
        );

    \I__6488\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29290\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__29290\,
            I => \tok.n174\
        );

    \I__6486\ : InMux
    port map (
            O => \N__29287\,
            I => \N__29282\
        );

    \I__6485\ : InMux
    port map (
            O => \N__29286\,
            I => \N__29277\
        );

    \I__6484\ : InMux
    port map (
            O => \N__29285\,
            I => \N__29277\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__29282\,
            I => \tok.n4_adj_702\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__29277\,
            I => \tok.n4_adj_702\
        );

    \I__6481\ : SRMux
    port map (
            O => \N__29272\,
            I => \N__29266\
        );

    \I__6480\ : SRMux
    port map (
            O => \N__29271\,
            I => \N__29263\
        );

    \I__6479\ : SRMux
    port map (
            O => \N__29270\,
            I => \N__29256\
        );

    \I__6478\ : SRMux
    port map (
            O => \N__29269\,
            I => \N__29251\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__29266\,
            I => \N__29246\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__29263\,
            I => \N__29246\
        );

    \I__6475\ : SRMux
    port map (
            O => \N__29262\,
            I => \N__29243\
        );

    \I__6474\ : SRMux
    port map (
            O => \N__29261\,
            I => \N__29238\
        );

    \I__6473\ : SRMux
    port map (
            O => \N__29260\,
            I => \N__29234\
        );

    \I__6472\ : SRMux
    port map (
            O => \N__29259\,
            I => \N__29231\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__29256\,
            I => \N__29227\
        );

    \I__6470\ : SRMux
    port map (
            O => \N__29255\,
            I => \N__29224\
        );

    \I__6469\ : SRMux
    port map (
            O => \N__29254\,
            I => \N__29221\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29217\
        );

    \I__6467\ : Span4Mux_s1_v
    port map (
            O => \N__29246\,
            I => \N__29211\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__29243\,
            I => \N__29211\
        );

    \I__6465\ : SRMux
    port map (
            O => \N__29242\,
            I => \N__29208\
        );

    \I__6464\ : SRMux
    port map (
            O => \N__29241\,
            I => \N__29205\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__29238\,
            I => \N__29201\
        );

    \I__6462\ : SRMux
    port map (
            O => \N__29237\,
            I => \N__29198\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__29234\,
            I => \N__29195\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__29231\,
            I => \N__29192\
        );

    \I__6459\ : SRMux
    port map (
            O => \N__29230\,
            I => \N__29189\
        );

    \I__6458\ : Span4Mux_v
    port map (
            O => \N__29227\,
            I => \N__29184\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__29224\,
            I => \N__29184\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__29221\,
            I => \N__29181\
        );

    \I__6455\ : SRMux
    port map (
            O => \N__29220\,
            I => \N__29176\
        );

    \I__6454\ : Span4Mux_v
    port map (
            O => \N__29217\,
            I => \N__29173\
        );

    \I__6453\ : SRMux
    port map (
            O => \N__29216\,
            I => \N__29170\
        );

    \I__6452\ : Span4Mux_v
    port map (
            O => \N__29211\,
            I => \N__29163\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__29208\,
            I => \N__29163\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__29205\,
            I => \N__29160\
        );

    \I__6449\ : SRMux
    port map (
            O => \N__29204\,
            I => \N__29157\
        );

    \I__6448\ : Span4Mux_v
    port map (
            O => \N__29201\,
            I => \N__29152\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__29198\,
            I => \N__29152\
        );

    \I__6446\ : Span4Mux_h
    port map (
            O => \N__29195\,
            I => \N__29149\
        );

    \I__6445\ : Span4Mux_v
    port map (
            O => \N__29192\,
            I => \N__29144\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__29189\,
            I => \N__29144\
        );

    \I__6443\ : Span4Mux_v
    port map (
            O => \N__29184\,
            I => \N__29141\
        );

    \I__6442\ : Span4Mux_v
    port map (
            O => \N__29181\,
            I => \N__29138\
        );

    \I__6441\ : SRMux
    port map (
            O => \N__29180\,
            I => \N__29135\
        );

    \I__6440\ : SRMux
    port map (
            O => \N__29179\,
            I => \N__29132\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__29176\,
            I => \N__29129\
        );

    \I__6438\ : Span4Mux_v
    port map (
            O => \N__29173\,
            I => \N__29124\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__29170\,
            I => \N__29124\
        );

    \I__6436\ : SRMux
    port map (
            O => \N__29169\,
            I => \N__29121\
        );

    \I__6435\ : SRMux
    port map (
            O => \N__29168\,
            I => \N__29118\
        );

    \I__6434\ : Span4Mux_v
    port map (
            O => \N__29163\,
            I => \N__29113\
        );

    \I__6433\ : Span4Mux_h
    port map (
            O => \N__29160\,
            I => \N__29108\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__29157\,
            I => \N__29108\
        );

    \I__6431\ : Span4Mux_h
    port map (
            O => \N__29152\,
            I => \N__29105\
        );

    \I__6430\ : Span4Mux_v
    port map (
            O => \N__29149\,
            I => \N__29100\
        );

    \I__6429\ : Span4Mux_h
    port map (
            O => \N__29144\,
            I => \N__29100\
        );

    \I__6428\ : IoSpan4Mux
    port map (
            O => \N__29141\,
            I => \N__29097\
        );

    \I__6427\ : Span4Mux_h
    port map (
            O => \N__29138\,
            I => \N__29092\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__29135\,
            I => \N__29092\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__29132\,
            I => \N__29089\
        );

    \I__6424\ : Span4Mux_v
    port map (
            O => \N__29129\,
            I => \N__29086\
        );

    \I__6423\ : Span4Mux_v
    port map (
            O => \N__29124\,
            I => \N__29081\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__29121\,
            I => \N__29081\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__29118\,
            I => \N__29078\
        );

    \I__6420\ : SRMux
    port map (
            O => \N__29117\,
            I => \N__29075\
        );

    \I__6419\ : SRMux
    port map (
            O => \N__29116\,
            I => \N__29072\
        );

    \I__6418\ : Span4Mux_h
    port map (
            O => \N__29113\,
            I => \N__29067\
        );

    \I__6417\ : Span4Mux_v
    port map (
            O => \N__29108\,
            I => \N__29067\
        );

    \I__6416\ : Span4Mux_h
    port map (
            O => \N__29105\,
            I => \N__29062\
        );

    \I__6415\ : Span4Mux_h
    port map (
            O => \N__29100\,
            I => \N__29062\
        );

    \I__6414\ : Span4Mux_s0_v
    port map (
            O => \N__29097\,
            I => \N__29057\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__29092\,
            I => \N__29057\
        );

    \I__6412\ : Span4Mux_v
    port map (
            O => \N__29089\,
            I => \N__29054\
        );

    \I__6411\ : Span4Mux_h
    port map (
            O => \N__29086\,
            I => \N__29049\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__29081\,
            I => \N__29049\
        );

    \I__6409\ : Span4Mux_h
    port map (
            O => \N__29078\,
            I => \N__29046\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__29075\,
            I => \N__29043\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__29072\,
            I => \N__29040\
        );

    \I__6406\ : Span4Mux_v
    port map (
            O => \N__29067\,
            I => \N__29037\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__29062\,
            I => \N__29034\
        );

    \I__6404\ : Span4Mux_h
    port map (
            O => \N__29057\,
            I => \N__29029\
        );

    \I__6403\ : Span4Mux_h
    port map (
            O => \N__29054\,
            I => \N__29029\
        );

    \I__6402\ : Span4Mux_h
    port map (
            O => \N__29049\,
            I => \N__29024\
        );

    \I__6401\ : Span4Mux_v
    port map (
            O => \N__29046\,
            I => \N__29024\
        );

    \I__6400\ : Span12Mux_h
    port map (
            O => \N__29043\,
            I => \N__29019\
        );

    \I__6399\ : Sp12to4
    port map (
            O => \N__29040\,
            I => \N__29019\
        );

    \I__6398\ : Odrv4
    port map (
            O => \N__29037\,
            I => \tok.reset_N_2\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__29034\,
            I => \tok.reset_N_2\
        );

    \I__6396\ : Odrv4
    port map (
            O => \N__29029\,
            I => \tok.reset_N_2\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__29024\,
            I => \tok.reset_N_2\
        );

    \I__6394\ : Odrv12
    port map (
            O => \N__29019\,
            I => \tok.reset_N_2\
        );

    \I__6393\ : InMux
    port map (
            O => \N__29008\,
            I => \N__29005\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__29005\,
            I => \N__29002\
        );

    \I__6391\ : Odrv4
    port map (
            O => \N__29002\,
            I => \tok.n256_adj_749\
        );

    \I__6390\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28996\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__28996\,
            I => \tok.n367\
        );

    \I__6388\ : InMux
    port map (
            O => \N__28993\,
            I => \N__28990\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__28990\,
            I => \N__28987\
        );

    \I__6386\ : Span12Mux_s8_h
    port map (
            O => \N__28987\,
            I => \N__28984\
        );

    \I__6385\ : Odrv12
    port map (
            O => \N__28984\,
            I => \tok.n215_adj_750\
        );

    \I__6384\ : CascadeMux
    port map (
            O => \N__28981\,
            I => \N__28974\
        );

    \I__6383\ : InMux
    port map (
            O => \N__28980\,
            I => \N__28966\
        );

    \I__6382\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28966\
        );

    \I__6381\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28959\
        );

    \I__6380\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28959\
        );

    \I__6379\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28959\
        );

    \I__6378\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28956\
        );

    \I__6377\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28953\
        );

    \I__6376\ : InMux
    port map (
            O => \N__28971\,
            I => \N__28950\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__28966\,
            I => \tok.depth_2\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__28959\,
            I => \tok.depth_2\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__28956\,
            I => \tok.depth_2\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__28953\,
            I => \tok.depth_2\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__28950\,
            I => \tok.depth_2\
        );

    \I__6370\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28936\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__28936\,
            I => \N__28932\
        );

    \I__6368\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28929\
        );

    \I__6367\ : Span4Mux_h
    port map (
            O => \N__28932\,
            I => \N__28926\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__28929\,
            I => \tok.tail_47\
        );

    \I__6365\ : Odrv4
    port map (
            O => \N__28926\,
            I => \tok.tail_47\
        );

    \I__6364\ : CEMux
    port map (
            O => \N__28921\,
            I => \N__28914\
        );

    \I__6363\ : CEMux
    port map (
            O => \N__28920\,
            I => \N__28911\
        );

    \I__6362\ : CEMux
    port map (
            O => \N__28919\,
            I => \N__28906\
        );

    \I__6361\ : CEMux
    port map (
            O => \N__28918\,
            I => \N__28902\
        );

    \I__6360\ : CEMux
    port map (
            O => \N__28917\,
            I => \N__28899\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__28914\,
            I => \N__28896\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__28911\,
            I => \N__28893\
        );

    \I__6357\ : CEMux
    port map (
            O => \N__28910\,
            I => \N__28890\
        );

    \I__6356\ : CEMux
    port map (
            O => \N__28909\,
            I => \N__28886\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__28906\,
            I => \N__28883\
        );

    \I__6354\ : CEMux
    port map (
            O => \N__28905\,
            I => \N__28880\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__28902\,
            I => \N__28877\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__28899\,
            I => \N__28874\
        );

    \I__6351\ : Span4Mux_h
    port map (
            O => \N__28896\,
            I => \N__28866\
        );

    \I__6350\ : Span4Mux_s2_v
    port map (
            O => \N__28893\,
            I => \N__28866\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__28890\,
            I => \N__28866\
        );

    \I__6348\ : CEMux
    port map (
            O => \N__28889\,
            I => \N__28863\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__28886\,
            I => \N__28859\
        );

    \I__6346\ : Span4Mux_s2_v
    port map (
            O => \N__28883\,
            I => \N__28856\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__28880\,
            I => \N__28853\
        );

    \I__6344\ : Span4Mux_s2_v
    port map (
            O => \N__28877\,
            I => \N__28850\
        );

    \I__6343\ : Span4Mux_v
    port map (
            O => \N__28874\,
            I => \N__28847\
        );

    \I__6342\ : CEMux
    port map (
            O => \N__28873\,
            I => \N__28844\
        );

    \I__6341\ : Span4Mux_s2_h
    port map (
            O => \N__28866\,
            I => \N__28839\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__28863\,
            I => \N__28839\
        );

    \I__6339\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28836\
        );

    \I__6338\ : Span4Mux_s2_v
    port map (
            O => \N__28859\,
            I => \N__28827\
        );

    \I__6337\ : Span4Mux_h
    port map (
            O => \N__28856\,
            I => \N__28822\
        );

    \I__6336\ : Span4Mux_s2_v
    port map (
            O => \N__28853\,
            I => \N__28822\
        );

    \I__6335\ : Span4Mux_h
    port map (
            O => \N__28850\,
            I => \N__28817\
        );

    \I__6334\ : Span4Mux_s0_h
    port map (
            O => \N__28847\,
            I => \N__28817\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__28844\,
            I => \N__28812\
        );

    \I__6332\ : Sp12to4
    port map (
            O => \N__28839\,
            I => \N__28812\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__28836\,
            I => \N__28809\
        );

    \I__6330\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28806\
        );

    \I__6329\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28795\
        );

    \I__6328\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28795\
        );

    \I__6327\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28795\
        );

    \I__6326\ : InMux
    port map (
            O => \N__28831\,
            I => \N__28795\
        );

    \I__6325\ : InMux
    port map (
            O => \N__28830\,
            I => \N__28795\
        );

    \I__6324\ : Odrv4
    port map (
            O => \N__28827\,
            I => \rd_7__N_373\
        );

    \I__6323\ : Odrv4
    port map (
            O => \N__28822\,
            I => \rd_7__N_373\
        );

    \I__6322\ : Odrv4
    port map (
            O => \N__28817\,
            I => \rd_7__N_373\
        );

    \I__6321\ : Odrv12
    port map (
            O => \N__28812\,
            I => \rd_7__N_373\
        );

    \I__6320\ : Odrv4
    port map (
            O => \N__28809\,
            I => \rd_7__N_373\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__28806\,
            I => \rd_7__N_373\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__28795\,
            I => \rd_7__N_373\
        );

    \I__6317\ : CascadeMux
    port map (
            O => \N__28780\,
            I => \N__28777\
        );

    \I__6316\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28773\
        );

    \I__6315\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28770\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__28773\,
            I => \N__28767\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__28770\,
            I => \N__28764\
        );

    \I__6312\ : Span4Mux_s2_h
    port map (
            O => \N__28767\,
            I => \N__28761\
        );

    \I__6311\ : Span4Mux_s1_h
    port map (
            O => \N__28764\,
            I => \N__28758\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__28761\,
            I => \tok.tail_55\
        );

    \I__6309\ : Odrv4
    port map (
            O => \N__28758\,
            I => \tok.tail_55\
        );

    \I__6308\ : InMux
    port map (
            O => \N__28753\,
            I => \N__28720\
        );

    \I__6307\ : InMux
    port map (
            O => \N__28752\,
            I => \N__28720\
        );

    \I__6306\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28720\
        );

    \I__6305\ : InMux
    port map (
            O => \N__28750\,
            I => \N__28720\
        );

    \I__6304\ : InMux
    port map (
            O => \N__28749\,
            I => \N__28720\
        );

    \I__6303\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28720\
        );

    \I__6302\ : InMux
    port map (
            O => \N__28747\,
            I => \N__28707\
        );

    \I__6301\ : InMux
    port map (
            O => \N__28746\,
            I => \N__28707\
        );

    \I__6300\ : InMux
    port map (
            O => \N__28745\,
            I => \N__28707\
        );

    \I__6299\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28707\
        );

    \I__6298\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28707\
        );

    \I__6297\ : InMux
    port map (
            O => \N__28742\,
            I => \N__28707\
        );

    \I__6296\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28694\
        );

    \I__6295\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28694\
        );

    \I__6294\ : InMux
    port map (
            O => \N__28739\,
            I => \N__28694\
        );

    \I__6293\ : InMux
    port map (
            O => \N__28738\,
            I => \N__28694\
        );

    \I__6292\ : InMux
    port map (
            O => \N__28737\,
            I => \N__28694\
        );

    \I__6291\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28694\
        );

    \I__6290\ : InMux
    port map (
            O => \N__28735\,
            I => \N__28686\
        );

    \I__6289\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28681\
        );

    \I__6288\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28681\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__28720\,
            I => \N__28671\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__28707\,
            I => \N__28666\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__28694\,
            I => \N__28666\
        );

    \I__6284\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28649\
        );

    \I__6283\ : InMux
    port map (
            O => \N__28692\,
            I => \N__28649\
        );

    \I__6282\ : InMux
    port map (
            O => \N__28691\,
            I => \N__28649\
        );

    \I__6281\ : InMux
    port map (
            O => \N__28690\,
            I => \N__28649\
        );

    \I__6280\ : InMux
    port map (
            O => \N__28689\,
            I => \N__28649\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__28686\,
            I => \N__28646\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__28681\,
            I => \N__28643\
        );

    \I__6277\ : InMux
    port map (
            O => \N__28680\,
            I => \N__28630\
        );

    \I__6276\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28630\
        );

    \I__6275\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28630\
        );

    \I__6274\ : InMux
    port map (
            O => \N__28677\,
            I => \N__28630\
        );

    \I__6273\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28630\
        );

    \I__6272\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28630\
        );

    \I__6271\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28603\
        );

    \I__6270\ : Span4Mux_s2_v
    port map (
            O => \N__28671\,
            I => \N__28600\
        );

    \I__6269\ : Span4Mux_h
    port map (
            O => \N__28666\,
            I => \N__28597\
        );

    \I__6268\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28584\
        );

    \I__6267\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28584\
        );

    \I__6266\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28584\
        );

    \I__6265\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28584\
        );

    \I__6264\ : InMux
    port map (
            O => \N__28661\,
            I => \N__28584\
        );

    \I__6263\ : InMux
    port map (
            O => \N__28660\,
            I => \N__28584\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__28649\,
            I => \N__28581\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__28646\,
            I => \N__28574\
        );

    \I__6260\ : Span4Mux_s2_v
    port map (
            O => \N__28643\,
            I => \N__28574\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__28630\,
            I => \N__28574\
        );

    \I__6258\ : InMux
    port map (
            O => \N__28629\,
            I => \N__28559\
        );

    \I__6257\ : InMux
    port map (
            O => \N__28628\,
            I => \N__28559\
        );

    \I__6256\ : InMux
    port map (
            O => \N__28627\,
            I => \N__28559\
        );

    \I__6255\ : InMux
    port map (
            O => \N__28626\,
            I => \N__28559\
        );

    \I__6254\ : InMux
    port map (
            O => \N__28625\,
            I => \N__28559\
        );

    \I__6253\ : InMux
    port map (
            O => \N__28624\,
            I => \N__28559\
        );

    \I__6252\ : InMux
    port map (
            O => \N__28623\,
            I => \N__28559\
        );

    \I__6251\ : InMux
    port map (
            O => \N__28622\,
            I => \N__28546\
        );

    \I__6250\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28546\
        );

    \I__6249\ : InMux
    port map (
            O => \N__28620\,
            I => \N__28546\
        );

    \I__6248\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28546\
        );

    \I__6247\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28546\
        );

    \I__6246\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28546\
        );

    \I__6245\ : InMux
    port map (
            O => \N__28616\,
            I => \N__28533\
        );

    \I__6244\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28533\
        );

    \I__6243\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28533\
        );

    \I__6242\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28533\
        );

    \I__6241\ : InMux
    port map (
            O => \N__28612\,
            I => \N__28533\
        );

    \I__6240\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28533\
        );

    \I__6239\ : InMux
    port map (
            O => \N__28610\,
            I => \N__28522\
        );

    \I__6238\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28522\
        );

    \I__6237\ : InMux
    port map (
            O => \N__28608\,
            I => \N__28522\
        );

    \I__6236\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28522\
        );

    \I__6235\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28522\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__28603\,
            I => \C_stk_delta_1\
        );

    \I__6233\ : Odrv4
    port map (
            O => \N__28600\,
            I => \C_stk_delta_1\
        );

    \I__6232\ : Odrv4
    port map (
            O => \N__28597\,
            I => \C_stk_delta_1\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__28584\,
            I => \C_stk_delta_1\
        );

    \I__6230\ : Odrv4
    port map (
            O => \N__28581\,
            I => \C_stk_delta_1\
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__28574\,
            I => \C_stk_delta_1\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__28559\,
            I => \C_stk_delta_1\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__28546\,
            I => \C_stk_delta_1\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__28533\,
            I => \C_stk_delta_1\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__28522\,
            I => \C_stk_delta_1\
        );

    \I__6224\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28498\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__28498\,
            I => \N__28495\
        );

    \I__6222\ : Span4Mux_s1_v
    port map (
            O => \N__28495\,
            I => \N__28491\
        );

    \I__6221\ : InMux
    port map (
            O => \N__28494\,
            I => \N__28488\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__28491\,
            I => \tok.tail_63\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__28488\,
            I => \tok.tail_63\
        );

    \I__6218\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28480\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__28480\,
            I => \N__28469\
        );

    \I__6216\ : InMux
    port map (
            O => \N__28479\,
            I => \N__28458\
        );

    \I__6215\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28458\
        );

    \I__6214\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28458\
        );

    \I__6213\ : InMux
    port map (
            O => \N__28476\,
            I => \N__28458\
        );

    \I__6212\ : InMux
    port map (
            O => \N__28475\,
            I => \N__28458\
        );

    \I__6211\ : InMux
    port map (
            O => \N__28474\,
            I => \N__28455\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__28473\,
            I => \N__28452\
        );

    \I__6209\ : InMux
    port map (
            O => \N__28472\,
            I => \N__28444\
        );

    \I__6208\ : Span4Mux_h
    port map (
            O => \N__28469\,
            I => \N__28441\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__28458\,
            I => \N__28438\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__28455\,
            I => \N__28435\
        );

    \I__6205\ : InMux
    port map (
            O => \N__28452\,
            I => \N__28426\
        );

    \I__6204\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28426\
        );

    \I__6203\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28426\
        );

    \I__6202\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28426\
        );

    \I__6201\ : InMux
    port map (
            O => \N__28448\,
            I => \N__28419\
        );

    \I__6200\ : InMux
    port map (
            O => \N__28447\,
            I => \N__28419\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__28444\,
            I => \N__28416\
        );

    \I__6198\ : Sp12to4
    port map (
            O => \N__28441\,
            I => \N__28413\
        );

    \I__6197\ : Span4Mux_s3_v
    port map (
            O => \N__28438\,
            I => \N__28410\
        );

    \I__6196\ : Span4Mux_v
    port map (
            O => \N__28435\,
            I => \N__28405\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__28426\,
            I => \N__28405\
        );

    \I__6194\ : InMux
    port map (
            O => \N__28425\,
            I => \N__28402\
        );

    \I__6193\ : InMux
    port map (
            O => \N__28424\,
            I => \N__28399\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__28419\,
            I => \N__28396\
        );

    \I__6191\ : Odrv12
    port map (
            O => \N__28416\,
            I => n15
        );

    \I__6190\ : Odrv12
    port map (
            O => \N__28413\,
            I => n15
        );

    \I__6189\ : Odrv4
    port map (
            O => \N__28410\,
            I => n15
        );

    \I__6188\ : Odrv4
    port map (
            O => \N__28405\,
            I => n15
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__28402\,
            I => n15
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__28399\,
            I => n15
        );

    \I__6185\ : Odrv4
    port map (
            O => \N__28396\,
            I => n15
        );

    \I__6184\ : InMux
    port map (
            O => \N__28381\,
            I => \N__28377\
        );

    \I__6183\ : InMux
    port map (
            O => \N__28380\,
            I => \N__28374\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__28377\,
            I => \N__28370\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__28374\,
            I => \N__28367\
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__28373\,
            I => \N__28364\
        );

    \I__6179\ : Span4Mux_s3_h
    port map (
            O => \N__28370\,
            I => \N__28360\
        );

    \I__6178\ : Span4Mux_s2_h
    port map (
            O => \N__28367\,
            I => \N__28357\
        );

    \I__6177\ : InMux
    port map (
            O => \N__28364\,
            I => \N__28352\
        );

    \I__6176\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28352\
        );

    \I__6175\ : Span4Mux_h
    port map (
            O => \N__28360\,
            I => \N__28349\
        );

    \I__6174\ : Span4Mux_h
    port map (
            O => \N__28357\,
            I => \N__28344\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__28352\,
            I => \N__28344\
        );

    \I__6172\ : Odrv4
    port map (
            O => \N__28349\,
            I => \tok.tc_plus_1_7\
        );

    \I__6171\ : Odrv4
    port map (
            O => \N__28344\,
            I => \tok.tc_plus_1_7\
        );

    \I__6170\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28335\
        );

    \I__6169\ : InMux
    port map (
            O => \N__28338\,
            I => \N__28331\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__28335\,
            I => \N__28325\
        );

    \I__6167\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28322\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__28331\,
            I => \N__28319\
        );

    \I__6165\ : CascadeMux
    port map (
            O => \N__28330\,
            I => \N__28316\
        );

    \I__6164\ : InMux
    port map (
            O => \N__28329\,
            I => \N__28313\
        );

    \I__6163\ : InMux
    port map (
            O => \N__28328\,
            I => \N__28310\
        );

    \I__6162\ : Span4Mux_v
    port map (
            O => \N__28325\,
            I => \N__28307\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__28322\,
            I => \N__28302\
        );

    \I__6160\ : Span4Mux_h
    port map (
            O => \N__28319\,
            I => \N__28302\
        );

    \I__6159\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28299\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__28313\,
            I => \N__28294\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__28310\,
            I => \N__28291\
        );

    \I__6156\ : Span4Mux_h
    port map (
            O => \N__28307\,
            I => \N__28286\
        );

    \I__6155\ : Span4Mux_v
    port map (
            O => \N__28302\,
            I => \N__28286\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__28299\,
            I => \N__28283\
        );

    \I__6153\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28280\
        );

    \I__6152\ : InMux
    port map (
            O => \N__28297\,
            I => \N__28277\
        );

    \I__6151\ : Span4Mux_v
    port map (
            O => \N__28294\,
            I => \N__28274\
        );

    \I__6150\ : Span4Mux_v
    port map (
            O => \N__28291\,
            I => \N__28271\
        );

    \I__6149\ : Span4Mux_h
    port map (
            O => \N__28286\,
            I => \N__28266\
        );

    \I__6148\ : Span4Mux_v
    port map (
            O => \N__28283\,
            I => \N__28266\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__28280\,
            I => \N__28263\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__28277\,
            I => \N__28258\
        );

    \I__6145\ : Span4Mux_v
    port map (
            O => \N__28274\,
            I => \N__28258\
        );

    \I__6144\ : Span4Mux_v
    port map (
            O => \N__28271\,
            I => \N__28253\
        );

    \I__6143\ : Span4Mux_v
    port map (
            O => \N__28266\,
            I => \N__28253\
        );

    \I__6142\ : Span12Mux_v
    port map (
            O => \N__28263\,
            I => \N__28250\
        );

    \I__6141\ : Odrv4
    port map (
            O => \N__28258\,
            I => \tok.S_7\
        );

    \I__6140\ : Odrv4
    port map (
            O => \N__28253\,
            I => \tok.S_7\
        );

    \I__6139\ : Odrv12
    port map (
            O => \N__28250\,
            I => \tok.S_7\
        );

    \I__6138\ : InMux
    port map (
            O => \N__28243\,
            I => \N__28240\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28237\
        );

    \I__6136\ : Span4Mux_v
    port map (
            O => \N__28237\,
            I => \N__28234\
        );

    \I__6135\ : Sp12to4
    port map (
            O => \N__28234\,
            I => \N__28231\
        );

    \I__6134\ : Span12Mux_h
    port map (
            O => \N__28231\,
            I => \N__28228\
        );

    \I__6133\ : Odrv12
    port map (
            O => \N__28228\,
            I => \tok.table_wr_data_7\
        );

    \I__6132\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28222\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__28222\,
            I => \N__28218\
        );

    \I__6130\ : InMux
    port map (
            O => \N__28221\,
            I => \N__28215\
        );

    \I__6129\ : Span4Mux_h
    port map (
            O => \N__28218\,
            I => \N__28212\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__28215\,
            I => uart_rx_data_4
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__28212\,
            I => uart_rx_data_4
        );

    \I__6126\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28204\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28200\
        );

    \I__6124\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28197\
        );

    \I__6123\ : Span4Mux_h
    port map (
            O => \N__28200\,
            I => \N__28194\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__28197\,
            I => uart_rx_data_2
        );

    \I__6121\ : Odrv4
    port map (
            O => \N__28194\,
            I => uart_rx_data_2
        );

    \I__6120\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28185\
        );

    \I__6119\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28182\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__28185\,
            I => \N__28179\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__28182\,
            I => uart_rx_data_1
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__28179\,
            I => uart_rx_data_1
        );

    \I__6115\ : InMux
    port map (
            O => \N__28174\,
            I => \N__28169\
        );

    \I__6114\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28164\
        );

    \I__6113\ : InMux
    port map (
            O => \N__28172\,
            I => \N__28164\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__28169\,
            I => capture_2
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__28164\,
            I => capture_2
        );

    \I__6110\ : CascadeMux
    port map (
            O => \N__28159\,
            I => \N__28155\
        );

    \I__6109\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28152\
        );

    \I__6108\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28149\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__28152\,
            I => \tok.tail_54\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__28149\,
            I => \tok.tail_54\
        );

    \I__6105\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28138\
        );

    \I__6104\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28138\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__28138\,
            I => \tok.C_stk.tail_38\
        );

    \I__6102\ : InMux
    port map (
            O => \N__28135\,
            I => \N__28131\
        );

    \I__6101\ : InMux
    port map (
            O => \N__28134\,
            I => \N__28128\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__28131\,
            I => \tok.tail_46\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__28128\,
            I => \tok.tail_46\
        );

    \I__6098\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28119\
        );

    \I__6097\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28113\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28110\
        );

    \I__6095\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28107\
        );

    \I__6094\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28104\
        );

    \I__6093\ : InMux
    port map (
            O => \N__28116\,
            I => \N__28099\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__28113\,
            I => \N__28095\
        );

    \I__6091\ : Span4Mux_s3_v
    port map (
            O => \N__28110\,
            I => \N__28088\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__28107\,
            I => \N__28088\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__28104\,
            I => \N__28088\
        );

    \I__6088\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28085\
        );

    \I__6087\ : InMux
    port map (
            O => \N__28102\,
            I => \N__28082\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__28099\,
            I => \N__28079\
        );

    \I__6085\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28076\
        );

    \I__6084\ : Span4Mux_s3_v
    port map (
            O => \N__28095\,
            I => \N__28071\
        );

    \I__6083\ : Span4Mux_h
    port map (
            O => \N__28088\,
            I => \N__28071\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__28085\,
            I => \N__28066\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__28082\,
            I => \N__28066\
        );

    \I__6080\ : Span4Mux_s0_v
    port map (
            O => \N__28079\,
            I => \N__28061\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__28076\,
            I => \N__28061\
        );

    \I__6078\ : Odrv4
    port map (
            O => \N__28071\,
            I => \tok.C_stk.n449\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__28066\,
            I => \tok.C_stk.n449\
        );

    \I__6076\ : Odrv4
    port map (
            O => \N__28061\,
            I => \tok.C_stk.n449\
        );

    \I__6075\ : InMux
    port map (
            O => \N__28054\,
            I => \N__28044\
        );

    \I__6074\ : InMux
    port map (
            O => \N__28053\,
            I => \N__28041\
        );

    \I__6073\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28038\
        );

    \I__6072\ : InMux
    port map (
            O => \N__28051\,
            I => \N__28035\
        );

    \I__6071\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28032\
        );

    \I__6070\ : InMux
    port map (
            O => \N__28049\,
            I => \N__28029\
        );

    \I__6069\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28026\
        );

    \I__6068\ : InMux
    port map (
            O => \N__28047\,
            I => \N__28023\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__28044\,
            I => \N__28020\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__28041\,
            I => \N__28015\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__28038\,
            I => \N__28015\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__28035\,
            I => \N__28010\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__28032\,
            I => \N__28010\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__28029\,
            I => \N__28005\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__28026\,
            I => \N__28005\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__28023\,
            I => \N__28001\
        );

    \I__6059\ : Span4Mux_s3_v
    port map (
            O => \N__28020\,
            I => \N__27996\
        );

    \I__6058\ : Span4Mux_h
    port map (
            O => \N__28015\,
            I => \N__27996\
        );

    \I__6057\ : Span4Mux_s2_v
    port map (
            O => \N__28010\,
            I => \N__27991\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__28005\,
            I => \N__27991\
        );

    \I__6055\ : InMux
    port map (
            O => \N__28004\,
            I => \N__27988\
        );

    \I__6054\ : Odrv12
    port map (
            O => \N__28001\,
            I => \tok.n273\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__27996\,
            I => \tok.n273\
        );

    \I__6052\ : Odrv4
    port map (
            O => \N__27991\,
            I => \tok.n273\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__27988\,
            I => \tok.n273\
        );

    \I__6050\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27974\
        );

    \I__6049\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27971\
        );

    \I__6048\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27967\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__27974\,
            I => \N__27964\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__27971\,
            I => \N__27961\
        );

    \I__6045\ : InMux
    port map (
            O => \N__27970\,
            I => \N__27958\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__27967\,
            I => \N__27955\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__27964\,
            I => tc_7
        );

    \I__6042\ : Odrv12
    port map (
            O => \N__27961\,
            I => tc_7
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__27958\,
            I => tc_7
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__27955\,
            I => tc_7
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__27946\,
            I => \tok.C_stk.n6227_cascade_\
        );

    \I__6038\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27937\
        );

    \I__6037\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27934\
        );

    \I__6036\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27930\
        );

    \I__6035\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27926\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27918\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__27934\,
            I => \N__27918\
        );

    \I__6032\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27915\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__27930\,
            I => \N__27912\
        );

    \I__6030\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27909\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27906\
        );

    \I__6028\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27903\
        );

    \I__6027\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27900\
        );

    \I__6026\ : InMux
    port map (
            O => \N__27923\,
            I => \N__27897\
        );

    \I__6025\ : Span4Mux_v
    port map (
            O => \N__27918\,
            I => \N__27894\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__27915\,
            I => \N__27891\
        );

    \I__6023\ : Span4Mux_v
    port map (
            O => \N__27912\,
            I => \N__27888\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__27909\,
            I => \N__27885\
        );

    \I__6021\ : Span4Mux_s1_v
    port map (
            O => \N__27906\,
            I => \N__27880\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__27903\,
            I => \N__27880\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__27900\,
            I => \N__27877\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__27897\,
            I => \N__27874\
        );

    \I__6017\ : Odrv4
    port map (
            O => \N__27894\,
            I => \tok.n15\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__27891\,
            I => \tok.n15\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__27888\,
            I => \tok.n15\
        );

    \I__6014\ : Odrv12
    port map (
            O => \N__27885\,
            I => \tok.n15\
        );

    \I__6013\ : Odrv4
    port map (
            O => \N__27880\,
            I => \tok.n15\
        );

    \I__6012\ : Odrv4
    port map (
            O => \N__27877\,
            I => \tok.n15\
        );

    \I__6011\ : Odrv12
    port map (
            O => \N__27874\,
            I => \tok.n15\
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__27859\,
            I => \N__27855\
        );

    \I__6009\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27846\
        );

    \I__6008\ : InMux
    port map (
            O => \N__27855\,
            I => \N__27846\
        );

    \I__6007\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27846\
        );

    \I__6006\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27843\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__27846\,
            I => \N__27840\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__27843\,
            I => \tok.c_stk_r_7\
        );

    \I__6003\ : Odrv12
    port map (
            O => \N__27840\,
            I => \tok.c_stk_r_7\
        );

    \I__6002\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27829\
        );

    \I__6001\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27829\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__27829\,
            I => \tok.C_stk.tail_7\
        );

    \I__5999\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27820\
        );

    \I__5998\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27820\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__27820\,
            I => \tok.tail_15\
        );

    \I__5996\ : CascadeMux
    port map (
            O => \N__27817\,
            I => \N__27814\
        );

    \I__5995\ : InMux
    port map (
            O => \N__27814\,
            I => \N__27808\
        );

    \I__5994\ : InMux
    port map (
            O => \N__27813\,
            I => \N__27808\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__27808\,
            I => \tok.C_stk.tail_23\
        );

    \I__5992\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27799\
        );

    \I__5991\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27799\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__27799\,
            I => \tok.tail_31\
        );

    \I__5989\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27790\
        );

    \I__5988\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27790\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__27790\,
            I => \tok.C_stk.tail_39\
        );

    \I__5986\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27784\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__27784\,
            I => reset_c
        );

    \I__5984\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27778\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__27778\,
            I => \N__27774\
        );

    \I__5982\ : CascadeMux
    port map (
            O => \N__27777\,
            I => \N__27771\
        );

    \I__5981\ : Span4Mux_h
    port map (
            O => \N__27774\,
            I => \N__27768\
        );

    \I__5980\ : InMux
    port map (
            O => \N__27771\,
            I => \N__27765\
        );

    \I__5979\ : Odrv4
    port map (
            O => \N__27768\,
            I => \tok.tail_50\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__27765\,
            I => \tok.tail_50\
        );

    \I__5977\ : InMux
    port map (
            O => \N__27760\,
            I => \N__27756\
        );

    \I__5976\ : InMux
    port map (
            O => \N__27759\,
            I => \N__27753\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__27756\,
            I => \tok.tail_58\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__27753\,
            I => \tok.tail_58\
        );

    \I__5973\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27745\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__27745\,
            I => \N__27742\
        );

    \I__5971\ : Span4Mux_s2_h
    port map (
            O => \N__27742\,
            I => \N__27739\
        );

    \I__5970\ : Span4Mux_h
    port map (
            O => \N__27739\,
            I => \N__27733\
        );

    \I__5969\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27730\
        );

    \I__5968\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27725\
        );

    \I__5967\ : InMux
    port map (
            O => \N__27736\,
            I => \N__27725\
        );

    \I__5966\ : Odrv4
    port map (
            O => \N__27733\,
            I => \tok.tc_plus_1_6\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__27730\,
            I => \tok.tc_plus_1_6\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__27725\,
            I => \tok.tc_plus_1_6\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__27718\,
            I => \tok.C_stk.n6233_cascade_\
        );

    \I__5962\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27712\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__27712\,
            I => \N__27708\
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__27711\,
            I => \N__27703\
        );

    \I__5959\ : Span4Mux_h
    port map (
            O => \N__27708\,
            I => \N__27700\
        );

    \I__5958\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27695\
        );

    \I__5957\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27695\
        );

    \I__5956\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27692\
        );

    \I__5955\ : Odrv4
    port map (
            O => \N__27700\,
            I => tc_6
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__27695\,
            I => tc_6
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__27692\,
            I => tc_6
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__27685\,
            I => \N__27681\
        );

    \I__5951\ : InMux
    port map (
            O => \N__27684\,
            I => \N__27673\
        );

    \I__5950\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27673\
        );

    \I__5949\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27673\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__27673\,
            I => \N__27669\
        );

    \I__5947\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27666\
        );

    \I__5946\ : Span4Mux_h
    port map (
            O => \N__27669\,
            I => \N__27663\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__27666\,
            I => \tok.c_stk_r_6\
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__27663\,
            I => \tok.c_stk_r_6\
        );

    \I__5943\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27652\
        );

    \I__5942\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27652\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__27652\,
            I => \tok.C_stk.tail_6\
        );

    \I__5940\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27643\
        );

    \I__5939\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27643\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__27643\,
            I => \tok.tail_14\
        );

    \I__5937\ : CascadeMux
    port map (
            O => \N__27640\,
            I => \N__27637\
        );

    \I__5936\ : InMux
    port map (
            O => \N__27637\,
            I => \N__27631\
        );

    \I__5935\ : InMux
    port map (
            O => \N__27636\,
            I => \N__27631\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__27631\,
            I => \tok.C_stk.tail_22\
        );

    \I__5933\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27622\
        );

    \I__5932\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27622\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__27622\,
            I => \tok.tail_30\
        );

    \I__5930\ : InMux
    port map (
            O => \N__27619\,
            I => \N__27616\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__27616\,
            I => \tok.n6641\
        );

    \I__5928\ : CascadeMux
    port map (
            O => \N__27613\,
            I => \tok.n266_cascade_\
        );

    \I__5927\ : InMux
    port map (
            O => \N__27610\,
            I => \N__27604\
        );

    \I__5926\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27604\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__27604\,
            I => \N__27601\
        );

    \I__5924\ : Span4Mux_v
    port map (
            O => \N__27601\,
            I => \N__27598\
        );

    \I__5923\ : Sp12to4
    port map (
            O => \N__27598\,
            I => \N__27595\
        );

    \I__5922\ : Odrv12
    port map (
            O => \N__27595\,
            I => \tok.n5_adj_713\
        );

    \I__5921\ : InMux
    port map (
            O => \N__27592\,
            I => \N__27589\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__27589\,
            I => \N__27586\
        );

    \I__5919\ : Span4Mux_h
    port map (
            O => \N__27586\,
            I => \N__27583\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__27583\,
            I => \tok.n256\
        );

    \I__5917\ : CascadeMux
    port map (
            O => \N__27580\,
            I => \tok.n4_adj_718_cascade_\
        );

    \I__5916\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27574\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__27574\,
            I => \N__27571\
        );

    \I__5914\ : Span4Mux_h
    port map (
            O => \N__27571\,
            I => \N__27568\
        );

    \I__5913\ : Span4Mux_v
    port map (
            O => \N__27568\,
            I => \N__27565\
        );

    \I__5912\ : Odrv4
    port map (
            O => \N__27565\,
            I => \tok.n221\
        );

    \I__5911\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27555\
        );

    \I__5910\ : CascadeMux
    port map (
            O => \N__27561\,
            I => \N__27548\
        );

    \I__5909\ : InMux
    port map (
            O => \N__27560\,
            I => \N__27545\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__27559\,
            I => \N__27537\
        );

    \I__5907\ : CascadeMux
    port map (
            O => \N__27558\,
            I => \N__27533\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__27555\,
            I => \N__27530\
        );

    \I__5905\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27525\
        );

    \I__5904\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27525\
        );

    \I__5903\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27520\
        );

    \I__5902\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27515\
        );

    \I__5901\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27515\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27511\
        );

    \I__5899\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27506\
        );

    \I__5898\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27501\
        );

    \I__5897\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27501\
        );

    \I__5896\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27498\
        );

    \I__5895\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27493\
        );

    \I__5894\ : InMux
    port map (
            O => \N__27537\,
            I => \N__27493\
        );

    \I__5893\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27490\
        );

    \I__5892\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27487\
        );

    \I__5891\ : Span4Mux_s3_v
    port map (
            O => \N__27530\,
            I => \N__27482\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__27525\,
            I => \N__27482\
        );

    \I__5889\ : InMux
    port map (
            O => \N__27524\,
            I => \N__27477\
        );

    \I__5888\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27477\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27472\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__27515\,
            I => \N__27472\
        );

    \I__5885\ : InMux
    port map (
            O => \N__27514\,
            I => \N__27468\
        );

    \I__5884\ : Sp12to4
    port map (
            O => \N__27511\,
            I => \N__27465\
        );

    \I__5883\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27462\
        );

    \I__5882\ : CascadeMux
    port map (
            O => \N__27509\,
            I => \N__27458\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__27506\,
            I => \N__27452\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__27501\,
            I => \N__27452\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__27498\,
            I => \N__27449\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__27493\,
            I => \N__27442\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__27490\,
            I => \N__27442\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__27487\,
            I => \N__27442\
        );

    \I__5875\ : Span4Mux_v
    port map (
            O => \N__27482\,
            I => \N__27435\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__27477\,
            I => \N__27435\
        );

    \I__5873\ : Span4Mux_v
    port map (
            O => \N__27472\,
            I => \N__27435\
        );

    \I__5872\ : InMux
    port map (
            O => \N__27471\,
            I => \N__27432\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__27468\,
            I => \N__27425\
        );

    \I__5870\ : Span12Mux_s6_v
    port map (
            O => \N__27465\,
            I => \N__27425\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__27462\,
            I => \N__27425\
        );

    \I__5868\ : InMux
    port map (
            O => \N__27461\,
            I => \N__27418\
        );

    \I__5867\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27418\
        );

    \I__5866\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27418\
        );

    \I__5865\ : Span4Mux_v
    port map (
            O => \N__27452\,
            I => \N__27409\
        );

    \I__5864\ : Span4Mux_v
    port map (
            O => \N__27449\,
            I => \N__27409\
        );

    \I__5863\ : Span4Mux_v
    port map (
            O => \N__27442\,
            I => \N__27409\
        );

    \I__5862\ : Span4Mux_h
    port map (
            O => \N__27435\,
            I => \N__27409\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__27432\,
            I => \tok.A_low_1\
        );

    \I__5860\ : Odrv12
    port map (
            O => \N__27425\,
            I => \tok.A_low_1\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__27418\,
            I => \tok.A_low_1\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__27409\,
            I => \tok.A_low_1\
        );

    \I__5857\ : InMux
    port map (
            O => \N__27400\,
            I => \N__27397\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__27397\,
            I => \tok.n2637\
        );

    \I__5855\ : CascadeMux
    port map (
            O => \N__27394\,
            I => \N__27383\
        );

    \I__5854\ : InMux
    port map (
            O => \N__27393\,
            I => \N__27379\
        );

    \I__5853\ : CascadeMux
    port map (
            O => \N__27392\,
            I => \N__27375\
        );

    \I__5852\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27371\
        );

    \I__5851\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27367\
        );

    \I__5850\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27364\
        );

    \I__5849\ : InMux
    port map (
            O => \N__27388\,
            I => \N__27359\
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__27387\,
            I => \N__27354\
        );

    \I__5847\ : InMux
    port map (
            O => \N__27386\,
            I => \N__27350\
        );

    \I__5846\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27347\
        );

    \I__5845\ : InMux
    port map (
            O => \N__27382\,
            I => \N__27343\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__27379\,
            I => \N__27340\
        );

    \I__5843\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27337\
        );

    \I__5842\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27334\
        );

    \I__5841\ : InMux
    port map (
            O => \N__27374\,
            I => \N__27331\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__27371\,
            I => \N__27328\
        );

    \I__5839\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27325\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__27367\,
            I => \N__27320\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__27364\,
            I => \N__27320\
        );

    \I__5836\ : InMux
    port map (
            O => \N__27363\,
            I => \N__27317\
        );

    \I__5835\ : InMux
    port map (
            O => \N__27362\,
            I => \N__27314\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__27359\,
            I => \N__27311\
        );

    \I__5833\ : InMux
    port map (
            O => \N__27358\,
            I => \N__27308\
        );

    \I__5832\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27301\
        );

    \I__5831\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27301\
        );

    \I__5830\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27301\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__27350\,
            I => \N__27298\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__27347\,
            I => \N__27295\
        );

    \I__5827\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27290\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__27343\,
            I => \N__27287\
        );

    \I__5825\ : Span4Mux_h
    port map (
            O => \N__27340\,
            I => \N__27284\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__27337\,
            I => \N__27277\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__27334\,
            I => \N__27277\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__27331\,
            I => \N__27277\
        );

    \I__5821\ : Span4Mux_v
    port map (
            O => \N__27328\,
            I => \N__27272\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__27325\,
            I => \N__27272\
        );

    \I__5819\ : Span4Mux_h
    port map (
            O => \N__27320\,
            I => \N__27269\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__27317\,
            I => \N__27266\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__27314\,
            I => \N__27263\
        );

    \I__5816\ : Span4Mux_h
    port map (
            O => \N__27311\,
            I => \N__27255\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__27308\,
            I => \N__27255\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__27301\,
            I => \N__27255\
        );

    \I__5813\ : Span4Mux_v
    port map (
            O => \N__27298\,
            I => \N__27250\
        );

    \I__5812\ : Span4Mux_h
    port map (
            O => \N__27295\,
            I => \N__27250\
        );

    \I__5811\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27245\
        );

    \I__5810\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27245\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__27290\,
            I => \N__27242\
        );

    \I__5808\ : Span4Mux_v
    port map (
            O => \N__27287\,
            I => \N__27233\
        );

    \I__5807\ : Span4Mux_v
    port map (
            O => \N__27284\,
            I => \N__27233\
        );

    \I__5806\ : Span4Mux_v
    port map (
            O => \N__27277\,
            I => \N__27233\
        );

    \I__5805\ : Span4Mux_h
    port map (
            O => \N__27272\,
            I => \N__27233\
        );

    \I__5804\ : Span4Mux_v
    port map (
            O => \N__27269\,
            I => \N__27226\
        );

    \I__5803\ : Span4Mux_h
    port map (
            O => \N__27266\,
            I => \N__27226\
        );

    \I__5802\ : Span4Mux_v
    port map (
            O => \N__27263\,
            I => \N__27226\
        );

    \I__5801\ : InMux
    port map (
            O => \N__27262\,
            I => \N__27223\
        );

    \I__5800\ : Span4Mux_h
    port map (
            O => \N__27255\,
            I => \N__27218\
        );

    \I__5799\ : Span4Mux_h
    port map (
            O => \N__27250\,
            I => \N__27218\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__27245\,
            I => \tok.A_low_4\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__27242\,
            I => \tok.A_low_4\
        );

    \I__5796\ : Odrv4
    port map (
            O => \N__27233\,
            I => \tok.A_low_4\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__27226\,
            I => \tok.A_low_4\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__27223\,
            I => \tok.A_low_4\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__27218\,
            I => \tok.A_low_4\
        );

    \I__5792\ : InMux
    port map (
            O => \N__27205\,
            I => \N__27202\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__27202\,
            I => \N__27199\
        );

    \I__5790\ : Span4Mux_v
    port map (
            O => \N__27199\,
            I => \N__27196\
        );

    \I__5789\ : Span4Mux_h
    port map (
            O => \N__27196\,
            I => \N__27193\
        );

    \I__5788\ : Odrv4
    port map (
            O => \N__27193\,
            I => \tok.uart.sender_6\
        );

    \I__5787\ : InMux
    port map (
            O => \N__27190\,
            I => \N__27187\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__27187\,
            I => \tok.uart.sender_7\
        );

    \I__5785\ : InMux
    port map (
            O => \N__27184\,
            I => \N__27181\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__27181\,
            I => \tok.uart.sender_8\
        );

    \I__5783\ : CEMux
    port map (
            O => \N__27178\,
            I => \N__27175\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__27175\,
            I => \N__27172\
        );

    \I__5781\ : Span4Mux_s3_h
    port map (
            O => \N__27172\,
            I => \N__27167\
        );

    \I__5780\ : CEMux
    port map (
            O => \N__27171\,
            I => \N__27164\
        );

    \I__5779\ : CEMux
    port map (
            O => \N__27170\,
            I => \N__27160\
        );

    \I__5778\ : Span4Mux_h
    port map (
            O => \N__27167\,
            I => \N__27155\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__27164\,
            I => \N__27155\
        );

    \I__5776\ : CEMux
    port map (
            O => \N__27163\,
            I => \N__27152\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__27160\,
            I => \N__27149\
        );

    \I__5774\ : Span4Mux_h
    port map (
            O => \N__27155\,
            I => \N__27144\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__27152\,
            I => \N__27144\
        );

    \I__5772\ : Span4Mux_h
    port map (
            O => \N__27149\,
            I => \N__27141\
        );

    \I__5771\ : Span4Mux_s1_v
    port map (
            O => \N__27144\,
            I => \N__27138\
        );

    \I__5770\ : Odrv4
    port map (
            O => \N__27141\,
            I => \tok.uart.n950\
        );

    \I__5769\ : Odrv4
    port map (
            O => \N__27138\,
            I => \tok.uart.n950\
        );

    \I__5768\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27130\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__27130\,
            I => \N__27126\
        );

    \I__5766\ : InMux
    port map (
            O => \N__27129\,
            I => \N__27123\
        );

    \I__5765\ : Span4Mux_v
    port map (
            O => \N__27126\,
            I => \N__27119\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__27123\,
            I => \N__27116\
        );

    \I__5763\ : InMux
    port map (
            O => \N__27122\,
            I => \N__27113\
        );

    \I__5762\ : Span4Mux_v
    port map (
            O => \N__27119\,
            I => \N__27110\
        );

    \I__5761\ : Span4Mux_h
    port map (
            O => \N__27116\,
            I => \N__27107\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__27113\,
            I => \N__27104\
        );

    \I__5759\ : Span4Mux_h
    port map (
            O => \N__27110\,
            I => \N__27099\
        );

    \I__5758\ : Span4Mux_v
    port map (
            O => \N__27107\,
            I => \N__27099\
        );

    \I__5757\ : Span4Mux_v
    port map (
            O => \N__27104\,
            I => \N__27096\
        );

    \I__5756\ : Odrv4
    port map (
            O => \N__27099\,
            I => \tok.n274\
        );

    \I__5755\ : Odrv4
    port map (
            O => \N__27096\,
            I => \tok.n274\
        );

    \I__5754\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27087\
        );

    \I__5753\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27084\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__27087\,
            I => \N__27080\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__27084\,
            I => \N__27077\
        );

    \I__5750\ : InMux
    port map (
            O => \N__27083\,
            I => \N__27074\
        );

    \I__5749\ : Span4Mux_s2_h
    port map (
            O => \N__27080\,
            I => \N__27069\
        );

    \I__5748\ : Span4Mux_h
    port map (
            O => \N__27077\,
            I => \N__27069\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__27074\,
            I => \N__27066\
        );

    \I__5746\ : Span4Mux_v
    port map (
            O => \N__27069\,
            I => \N__27063\
        );

    \I__5745\ : Odrv4
    port map (
            O => \N__27066\,
            I => \tok.n185\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__27063\,
            I => \tok.n185\
        );

    \I__5743\ : InMux
    port map (
            O => \N__27058\,
            I => \N__27055\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__27055\,
            I => \N__27052\
        );

    \I__5741\ : Span4Mux_h
    port map (
            O => \N__27052\,
            I => \N__27049\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__27049\,
            I => \tok.n7410\
        );

    \I__5739\ : CascadeMux
    port map (
            O => \N__27046\,
            I => \tok.n2598_cascade_\
        );

    \I__5738\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27040\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__27040\,
            I => \N__27033\
        );

    \I__5736\ : InMux
    port map (
            O => \N__27039\,
            I => \N__27030\
        );

    \I__5735\ : InMux
    port map (
            O => \N__27038\,
            I => \N__27027\
        );

    \I__5734\ : InMux
    port map (
            O => \N__27037\,
            I => \N__27024\
        );

    \I__5733\ : InMux
    port map (
            O => \N__27036\,
            I => \N__27019\
        );

    \I__5732\ : Span4Mux_v
    port map (
            O => \N__27033\,
            I => \N__27013\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__27030\,
            I => \N__27013\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__27027\,
            I => \N__27008\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__27005\
        );

    \I__5728\ : InMux
    port map (
            O => \N__27023\,
            I => \N__27000\
        );

    \I__5727\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27000\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__27019\,
            I => \N__26997\
        );

    \I__5725\ : InMux
    port map (
            O => \N__27018\,
            I => \N__26994\
        );

    \I__5724\ : Span4Mux_s3_h
    port map (
            O => \N__27013\,
            I => \N__26991\
        );

    \I__5723\ : CascadeMux
    port map (
            O => \N__27012\,
            I => \N__26988\
        );

    \I__5722\ : InMux
    port map (
            O => \N__27011\,
            I => \N__26984\
        );

    \I__5721\ : Span12Mux_s8_v
    port map (
            O => \N__27008\,
            I => \N__26981\
        );

    \I__5720\ : Span4Mux_h
    port map (
            O => \N__27005\,
            I => \N__26976\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__27000\,
            I => \N__26976\
        );

    \I__5718\ : Span4Mux_h
    port map (
            O => \N__26997\,
            I => \N__26973\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__26994\,
            I => \N__26970\
        );

    \I__5716\ : Span4Mux_h
    port map (
            O => \N__26991\,
            I => \N__26967\
        );

    \I__5715\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26962\
        );

    \I__5714\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26962\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__26984\,
            I => \tok.n45\
        );

    \I__5712\ : Odrv12
    port map (
            O => \N__26981\,
            I => \tok.n45\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__26976\,
            I => \tok.n45\
        );

    \I__5710\ : Odrv4
    port map (
            O => \N__26973\,
            I => \tok.n45\
        );

    \I__5709\ : Odrv12
    port map (
            O => \N__26970\,
            I => \tok.n45\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__26967\,
            I => \tok.n45\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__26962\,
            I => \tok.n45\
        );

    \I__5706\ : InMux
    port map (
            O => \N__26947\,
            I => \N__26944\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__26944\,
            I => \N__26941\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__26941\,
            I => \tok.n6390\
        );

    \I__5703\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26934\
        );

    \I__5702\ : CascadeMux
    port map (
            O => \N__26937\,
            I => \N__26928\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__26934\,
            I => \N__26923\
        );

    \I__5700\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26920\
        );

    \I__5699\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26917\
        );

    \I__5698\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26912\
        );

    \I__5697\ : InMux
    port map (
            O => \N__26928\,
            I => \N__26912\
        );

    \I__5696\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26907\
        );

    \I__5695\ : InMux
    port map (
            O => \N__26926\,
            I => \N__26907\
        );

    \I__5694\ : Span4Mux_h
    port map (
            O => \N__26923\,
            I => \N__26899\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__26920\,
            I => \N__26899\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__26917\,
            I => \N__26899\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__26912\,
            I => \N__26894\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26894\
        );

    \I__5689\ : InMux
    port map (
            O => \N__26906\,
            I => \N__26891\
        );

    \I__5688\ : Span4Mux_h
    port map (
            O => \N__26899\,
            I => \N__26888\
        );

    \I__5687\ : Span4Mux_h
    port map (
            O => \N__26894\,
            I => \N__26883\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__26891\,
            I => \N__26883\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__26888\,
            I => \tok.n821\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__26883\,
            I => \tok.n821\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__26878\,
            I => \tok.n215_cascade_\
        );

    \I__5682\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26872\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__26872\,
            I => \N__26869\
        );

    \I__5680\ : Span4Mux_v
    port map (
            O => \N__26869\,
            I => \N__26866\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__26866\,
            I => \tok.n6547\
        );

    \I__5678\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26860\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__26860\,
            I => \N__26857\
        );

    \I__5676\ : Span4Mux_s2_h
    port map (
            O => \N__26857\,
            I => \N__26853\
        );

    \I__5675\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26850\
        );

    \I__5674\ : Span4Mux_v
    port map (
            O => \N__26853\,
            I => \N__26845\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__26850\,
            I => \N__26845\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__26845\,
            I => \tok.n4_adj_712\
        );

    \I__5671\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26839\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__26839\,
            I => \N__26835\
        );

    \I__5669\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26832\
        );

    \I__5668\ : Span4Mux_s3_h
    port map (
            O => \N__26835\,
            I => \N__26828\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__26832\,
            I => \N__26825\
        );

    \I__5666\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26822\
        );

    \I__5665\ : Span4Mux_v
    port map (
            O => \N__26828\,
            I => \N__26815\
        );

    \I__5664\ : Span4Mux_s3_h
    port map (
            O => \N__26825\,
            I => \N__26815\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__26822\,
            I => \N__26815\
        );

    \I__5662\ : Span4Mux_h
    port map (
            O => \N__26815\,
            I => \N__26812\
        );

    \I__5661\ : Span4Mux_h
    port map (
            O => \N__26812\,
            I => \N__26809\
        );

    \I__5660\ : Odrv4
    port map (
            O => \N__26809\,
            I => \tok.n238\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__26806\,
            I => \tok.n6650_cascade_\
        );

    \I__5658\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26799\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__26802\,
            I => \N__26794\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__26799\,
            I => \N__26789\
        );

    \I__5655\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26786\
        );

    \I__5654\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26781\
        );

    \I__5653\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26781\
        );

    \I__5652\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26776\
        );

    \I__5651\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26769\
        );

    \I__5650\ : Span4Mux_v
    port map (
            O => \N__26789\,
            I => \N__26762\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__26786\,
            I => \N__26762\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__26781\,
            I => \N__26759\
        );

    \I__5647\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26755\
        );

    \I__5646\ : InMux
    port map (
            O => \N__26779\,
            I => \N__26752\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__26776\,
            I => \N__26749\
        );

    \I__5644\ : InMux
    port map (
            O => \N__26775\,
            I => \N__26746\
        );

    \I__5643\ : InMux
    port map (
            O => \N__26774\,
            I => \N__26739\
        );

    \I__5642\ : InMux
    port map (
            O => \N__26773\,
            I => \N__26739\
        );

    \I__5641\ : InMux
    port map (
            O => \N__26772\,
            I => \N__26739\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__26769\,
            I => \N__26733\
        );

    \I__5639\ : InMux
    port map (
            O => \N__26768\,
            I => \N__26728\
        );

    \I__5638\ : InMux
    port map (
            O => \N__26767\,
            I => \N__26728\
        );

    \I__5637\ : Span4Mux_h
    port map (
            O => \N__26762\,
            I => \N__26723\
        );

    \I__5636\ : Span4Mux_h
    port map (
            O => \N__26759\,
            I => \N__26723\
        );

    \I__5635\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26720\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__26755\,
            I => \N__26717\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__26752\,
            I => \N__26714\
        );

    \I__5632\ : Span4Mux_v
    port map (
            O => \N__26749\,
            I => \N__26709\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26709\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__26739\,
            I => \N__26706\
        );

    \I__5629\ : InMux
    port map (
            O => \N__26738\,
            I => \N__26703\
        );

    \I__5628\ : InMux
    port map (
            O => \N__26737\,
            I => \N__26698\
        );

    \I__5627\ : InMux
    port map (
            O => \N__26736\,
            I => \N__26698\
        );

    \I__5626\ : Span4Mux_s1_v
    port map (
            O => \N__26733\,
            I => \N__26689\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__26728\,
            I => \N__26689\
        );

    \I__5624\ : Span4Mux_h
    port map (
            O => \N__26723\,
            I => \N__26689\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__26720\,
            I => \N__26689\
        );

    \I__5622\ : Span4Mux_v
    port map (
            O => \N__26717\,
            I => \N__26680\
        );

    \I__5621\ : Span4Mux_v
    port map (
            O => \N__26714\,
            I => \N__26680\
        );

    \I__5620\ : Span4Mux_h
    port map (
            O => \N__26709\,
            I => \N__26680\
        );

    \I__5619\ : Span4Mux_v
    port map (
            O => \N__26706\,
            I => \N__26680\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__26703\,
            I => \tok.n48\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__26698\,
            I => \tok.n48\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__26689\,
            I => \tok.n48\
        );

    \I__5615\ : Odrv4
    port map (
            O => \N__26680\,
            I => \tok.n48\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__26671\,
            I => \tok.n211_cascade_\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__26668\,
            I => \N__26665\
        );

    \I__5612\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26662\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__26662\,
            I => \N__26659\
        );

    \I__5610\ : Span4Mux_s3_v
    port map (
            O => \N__26659\,
            I => \N__26656\
        );

    \I__5609\ : Span4Mux_h
    port map (
            O => \N__26656\,
            I => \N__26653\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__26653\,
            I => \N__26650\
        );

    \I__5607\ : Span4Mux_v
    port map (
            O => \N__26650\,
            I => \N__26647\
        );

    \I__5606\ : Odrv4
    port map (
            O => \N__26647\,
            I => \tok.n6644\
        );

    \I__5605\ : CascadeMux
    port map (
            O => \N__26644\,
            I => \tok.n260_cascade_\
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__26641\,
            I => \N__26638\
        );

    \I__5603\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26635\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__26635\,
            I => \N__26632\
        );

    \I__5601\ : Odrv4
    port map (
            O => \N__26632\,
            I => \tok.n6501\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__26629\,
            I => \tok.n186_adj_798_cascade_\
        );

    \I__5599\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26623\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__26623\,
            I => \N__26620\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__26620\,
            I => \tok.n6496\
        );

    \I__5596\ : CascadeMux
    port map (
            O => \N__26617\,
            I => \N__26612\
        );

    \I__5595\ : CascadeMux
    port map (
            O => \N__26616\,
            I => \N__26605\
        );

    \I__5594\ : CascadeMux
    port map (
            O => \N__26615\,
            I => \N__26602\
        );

    \I__5593\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26597\
        );

    \I__5592\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26597\
        );

    \I__5591\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26594\
        );

    \I__5590\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26591\
        );

    \I__5589\ : InMux
    port map (
            O => \N__26608\,
            I => \N__26588\
        );

    \I__5588\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26578\
        );

    \I__5587\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26578\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__26597\,
            I => \N__26575\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__26594\,
            I => \N__26570\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26570\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__26588\,
            I => \N__26567\
        );

    \I__5582\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26564\
        );

    \I__5581\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26561\
        );

    \I__5580\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26556\
        );

    \I__5579\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26556\
        );

    \I__5578\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26553\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__26578\,
            I => \N__26548\
        );

    \I__5576\ : Span4Mux_h
    port map (
            O => \N__26575\,
            I => \N__26548\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__26570\,
            I => \N__26543\
        );

    \I__5574\ : Span4Mux_h
    port map (
            O => \N__26567\,
            I => \N__26543\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__26564\,
            I => \tok.n194\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__26561\,
            I => \tok.n194\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__26556\,
            I => \tok.n194\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__26553\,
            I => \tok.n194\
        );

    \I__5569\ : Odrv4
    port map (
            O => \N__26548\,
            I => \tok.n194\
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__26543\,
            I => \tok.n194\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__26530\,
            I => \tok.n338_adj_805_cascade_\
        );

    \I__5566\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26524\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__26524\,
            I => \N__26521\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__26521\,
            I => \N__26518\
        );

    \I__5563\ : Span4Mux_v
    port map (
            O => \N__26518\,
            I => \N__26515\
        );

    \I__5562\ : Odrv4
    port map (
            O => \N__26515\,
            I => \tok.n6608\
        );

    \I__5561\ : InMux
    port map (
            O => \N__26512\,
            I => \N__26508\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__26511\,
            I => \N__26505\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__26508\,
            I => \N__26501\
        );

    \I__5558\ : InMux
    port map (
            O => \N__26505\,
            I => \N__26497\
        );

    \I__5557\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26493\
        );

    \I__5556\ : Span4Mux_h
    port map (
            O => \N__26501\,
            I => \N__26490\
        );

    \I__5555\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26487\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__26497\,
            I => \N__26484\
        );

    \I__5553\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26480\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__26493\,
            I => \N__26477\
        );

    \I__5551\ : Span4Mux_v
    port map (
            O => \N__26490\,
            I => \N__26474\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__26487\,
            I => \N__26469\
        );

    \I__5549\ : Span4Mux_h
    port map (
            O => \N__26484\,
            I => \N__26469\
        );

    \I__5548\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26466\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__26480\,
            I => \N__26463\
        );

    \I__5546\ : Span4Mux_h
    port map (
            O => \N__26477\,
            I => \N__26458\
        );

    \I__5545\ : Span4Mux_h
    port map (
            O => \N__26474\,
            I => \N__26458\
        );

    \I__5544\ : Span4Mux_v
    port map (
            O => \N__26469\,
            I => \N__26453\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__26466\,
            I => \N__26453\
        );

    \I__5542\ : Odrv4
    port map (
            O => \N__26463\,
            I => \tok.n219\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__26458\,
            I => \tok.n219\
        );

    \I__5540\ : Odrv4
    port map (
            O => \N__26453\,
            I => \tok.n219\
        );

    \I__5539\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26440\
        );

    \I__5538\ : InMux
    port map (
            O => \N__26445\,
            I => \N__26440\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__26440\,
            I => \N__26437\
        );

    \I__5536\ : Odrv4
    port map (
            O => \N__26437\,
            I => \tok.n190_adj_792\
        );

    \I__5535\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26431\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__26431\,
            I => \N__26428\
        );

    \I__5533\ : Odrv12
    port map (
            O => \N__26428\,
            I => \tok.n4_adj_804\
        );

    \I__5532\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26422\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__26422\,
            I => \N__26419\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__26419\,
            I => \tok.n174_adj_803\
        );

    \I__5529\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26413\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__26413\,
            I => \tok.n205_adj_806\
        );

    \I__5527\ : InMux
    port map (
            O => \N__26410\,
            I => \N__26407\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__26407\,
            I => \N__26404\
        );

    \I__5525\ : Span4Mux_v
    port map (
            O => \N__26404\,
            I => \N__26401\
        );

    \I__5524\ : Span4Mux_h
    port map (
            O => \N__26401\,
            I => \N__26398\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__26398\,
            I => \tok.n177_adj_813\
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__26395\,
            I => \tok.n252_adj_801_cascade_\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__26392\,
            I => \N__26388\
        );

    \I__5520\ : CascadeMux
    port map (
            O => \N__26391\,
            I => \N__26385\
        );

    \I__5519\ : InMux
    port map (
            O => \N__26388\,
            I => \N__26380\
        );

    \I__5518\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26377\
        );

    \I__5517\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26374\
        );

    \I__5516\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26371\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__26380\,
            I => \N__26368\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__26377\,
            I => \N__26365\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__26374\,
            I => \N__26360\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__26371\,
            I => \N__26360\
        );

    \I__5511\ : Span4Mux_h
    port map (
            O => \N__26368\,
            I => \N__26355\
        );

    \I__5510\ : Span4Mux_s3_h
    port map (
            O => \N__26365\,
            I => \N__26355\
        );

    \I__5509\ : Odrv12
    port map (
            O => \N__26360\,
            I => \tok.n867\
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__26355\,
            I => \tok.n867\
        );

    \I__5507\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26346\
        );

    \I__5506\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26343\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26340\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__26343\,
            I => \N__26337\
        );

    \I__5503\ : Span4Mux_s2_h
    port map (
            O => \N__26340\,
            I => \N__26334\
        );

    \I__5502\ : Span4Mux_h
    port map (
            O => \N__26337\,
            I => \N__26331\
        );

    \I__5501\ : Span4Mux_h
    port map (
            O => \N__26334\,
            I => \N__26328\
        );

    \I__5500\ : Span4Mux_h
    port map (
            O => \N__26331\,
            I => \N__26325\
        );

    \I__5499\ : Span4Mux_h
    port map (
            O => \N__26328\,
            I => \N__26322\
        );

    \I__5498\ : Odrv4
    port map (
            O => \N__26325\,
            I => \tok.n233\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__26322\,
            I => \tok.n233\
        );

    \I__5496\ : InMux
    port map (
            O => \N__26317\,
            I => \N__26312\
        );

    \I__5495\ : InMux
    port map (
            O => \N__26316\,
            I => \N__26309\
        );

    \I__5494\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26306\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__26312\,
            I => \N__26302\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__26309\,
            I => \N__26299\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__26306\,
            I => \N__26296\
        );

    \I__5490\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26293\
        );

    \I__5489\ : Span4Mux_v
    port map (
            O => \N__26302\,
            I => \N__26288\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__26299\,
            I => \N__26288\
        );

    \I__5487\ : Span4Mux_v
    port map (
            O => \N__26296\,
            I => \N__26282\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__26293\,
            I => \N__26282\
        );

    \I__5485\ : Span4Mux_h
    port map (
            O => \N__26288\,
            I => \N__26279\
        );

    \I__5484\ : InMux
    port map (
            O => \N__26287\,
            I => \N__26276\
        );

    \I__5483\ : Odrv4
    port map (
            O => \N__26282\,
            I => \tok.n5_adj_745\
        );

    \I__5482\ : Odrv4
    port map (
            O => \N__26279\,
            I => \tok.n5_adj_745\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__26276\,
            I => \tok.n5_adj_745\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__26269\,
            I => \tok.n255_adj_793_cascade_\
        );

    \I__5479\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26263\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__26263\,
            I => \tok.n258_adj_800\
        );

    \I__5477\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26256\
        );

    \I__5476\ : InMux
    port map (
            O => \N__26259\,
            I => \N__26253\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__26256\,
            I => \N__26250\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__26253\,
            I => \N__26247\
        );

    \I__5473\ : Sp12to4
    port map (
            O => \N__26250\,
            I => \N__26244\
        );

    \I__5472\ : Span12Mux_s11_v
    port map (
            O => \N__26247\,
            I => \N__26241\
        );

    \I__5471\ : Odrv12
    port map (
            O => \N__26244\,
            I => \tok.n6183\
        );

    \I__5470\ : Odrv12
    port map (
            O => \N__26241\,
            I => \tok.n6183\
        );

    \I__5469\ : CascadeMux
    port map (
            O => \N__26236\,
            I => \tok.n6162_cascade_\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__26233\,
            I => \tok.n865_cascade_\
        );

    \I__5467\ : CascadeMux
    port map (
            O => \N__26230\,
            I => \tok.n222_cascade_\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__26227\,
            I => \N__26223\
        );

    \I__5465\ : CascadeMux
    port map (
            O => \N__26226\,
            I => \N__26218\
        );

    \I__5464\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26214\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__26222\,
            I => \N__26211\
        );

    \I__5462\ : CascadeMux
    port map (
            O => \N__26221\,
            I => \N__26208\
        );

    \I__5461\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26204\
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__26217\,
            I => \N__26201\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__26214\,
            I => \N__26198\
        );

    \I__5458\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26195\
        );

    \I__5457\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26192\
        );

    \I__5456\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26189\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__26204\,
            I => \N__26186\
        );

    \I__5454\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26183\
        );

    \I__5453\ : Span4Mux_h
    port map (
            O => \N__26198\,
            I => \N__26176\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__26195\,
            I => \N__26176\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__26192\,
            I => \N__26173\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__26189\,
            I => \N__26166\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__26186\,
            I => \N__26166\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26166\
        );

    \I__5447\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26163\
        );

    \I__5446\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26160\
        );

    \I__5445\ : Span4Mux_v
    port map (
            O => \N__26176\,
            I => \N__26157\
        );

    \I__5444\ : Span4Mux_v
    port map (
            O => \N__26173\,
            I => \N__26152\
        );

    \I__5443\ : Span4Mux_v
    port map (
            O => \N__26166\,
            I => \N__26152\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__26163\,
            I => \N__26147\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__26160\,
            I => \N__26147\
        );

    \I__5440\ : Span4Mux_h
    port map (
            O => \N__26157\,
            I => \N__26144\
        );

    \I__5439\ : Span4Mux_h
    port map (
            O => \N__26152\,
            I => \N__26141\
        );

    \I__5438\ : Span12Mux_s4_h
    port map (
            O => \N__26147\,
            I => \N__26138\
        );

    \I__5437\ : Odrv4
    port map (
            O => \N__26144\,
            I => \tok.n245\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__26141\,
            I => \tok.n245\
        );

    \I__5435\ : Odrv12
    port map (
            O => \N__26138\,
            I => \tok.n245\
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__26131\,
            I => \N__26126\
        );

    \I__5433\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26123\
        );

    \I__5432\ : InMux
    port map (
            O => \N__26129\,
            I => \N__26120\
        );

    \I__5431\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26117\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__26123\,
            I => \N__26114\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__26120\,
            I => \N__26111\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__26117\,
            I => \N__26106\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__26114\,
            I => \N__26106\
        );

    \I__5426\ : Span4Mux_h
    port map (
            O => \N__26111\,
            I => \N__26103\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__26106\,
            I => \tok.n4_adj_648\
        );

    \I__5424\ : Odrv4
    port map (
            O => \N__26103\,
            I => \tok.n4_adj_648\
        );

    \I__5423\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26095\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__26095\,
            I => \N__26092\
        );

    \I__5421\ : Span4Mux_v
    port map (
            O => \N__26092\,
            I => \N__26089\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__26089\,
            I => \N__26086\
        );

    \I__5419\ : Span4Mux_h
    port map (
            O => \N__26086\,
            I => \N__26083\
        );

    \I__5418\ : Odrv4
    port map (
            O => \N__26083\,
            I => \tok.n2635\
        );

    \I__5417\ : CascadeMux
    port map (
            O => \N__26080\,
            I => \tok.n6653_cascade_\
        );

    \I__5416\ : CascadeMux
    port map (
            O => \N__26077\,
            I => \tok.n6646_cascade_\
        );

    \I__5415\ : CascadeMux
    port map (
            O => \N__26074\,
            I => \N__26071\
        );

    \I__5414\ : InMux
    port map (
            O => \N__26071\,
            I => \N__26068\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__26068\,
            I => \tok.n6167\
        );

    \I__5412\ : InMux
    port map (
            O => \N__26065\,
            I => \N__26062\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__26062\,
            I => \N__26059\
        );

    \I__5410\ : Span4Mux_v
    port map (
            O => \N__26059\,
            I => \N__26056\
        );

    \I__5409\ : Odrv4
    port map (
            O => \N__26056\,
            I => \tok.n6645\
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__26053\,
            I => \N__26050\
        );

    \I__5407\ : InMux
    port map (
            O => \N__26050\,
            I => \N__26047\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__26047\,
            I => \N__26044\
        );

    \I__5405\ : Span4Mux_h
    port map (
            O => \N__26044\,
            I => \N__26041\
        );

    \I__5404\ : Odrv4
    port map (
            O => \N__26041\,
            I => \tok.n247\
        );

    \I__5403\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26035\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__26035\,
            I => \tok.n6639\
        );

    \I__5401\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__26029\,
            I => \tok.n280\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__26026\,
            I => \tok.n6638_cascade_\
        );

    \I__5398\ : InMux
    port map (
            O => \N__26023\,
            I => \N__26020\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__26020\,
            I => \N__26017\
        );

    \I__5396\ : Odrv4
    port map (
            O => \N__26017\,
            I => \tok.n6636\
        );

    \I__5395\ : InMux
    port map (
            O => \N__26014\,
            I => \N__26010\
        );

    \I__5394\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26007\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__26010\,
            I => \N__26004\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__26007\,
            I => \N__25999\
        );

    \I__5391\ : Span4Mux_v
    port map (
            O => \N__26004\,
            I => \N__25999\
        );

    \I__5390\ : Span4Mux_h
    port map (
            O => \N__25999\,
            I => \N__25996\
        );

    \I__5389\ : Odrv4
    port map (
            O => \N__25996\,
            I => \tok.n260_adj_717\
        );

    \I__5388\ : InMux
    port map (
            O => \N__25993\,
            I => \N__25989\
        );

    \I__5387\ : CascadeMux
    port map (
            O => \N__25992\,
            I => \N__25985\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__25989\,
            I => \N__25981\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__25988\,
            I => \N__25978\
        );

    \I__5384\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25975\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__25984\,
            I => \N__25972\
        );

    \I__5382\ : Span4Mux_v
    port map (
            O => \N__25981\,
            I => \N__25968\
        );

    \I__5381\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25965\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__25975\,
            I => \N__25961\
        );

    \I__5379\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25958\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__25971\,
            I => \N__25955\
        );

    \I__5377\ : Span4Mux_h
    port map (
            O => \N__25968\,
            I => \N__25950\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__25965\,
            I => \N__25950\
        );

    \I__5375\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25947\
        );

    \I__5374\ : Span4Mux_v
    port map (
            O => \N__25961\,
            I => \N__25944\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__25958\,
            I => \N__25941\
        );

    \I__5372\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25938\
        );

    \I__5371\ : Span4Mux_v
    port map (
            O => \N__25950\,
            I => \N__25933\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__25947\,
            I => \N__25930\
        );

    \I__5369\ : Span4Mux_h
    port map (
            O => \N__25944\,
            I => \N__25927\
        );

    \I__5368\ : Span4Mux_v
    port map (
            O => \N__25941\,
            I => \N__25924\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__25938\,
            I => \N__25921\
        );

    \I__5366\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25918\
        );

    \I__5365\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25915\
        );

    \I__5364\ : Span4Mux_h
    port map (
            O => \N__25933\,
            I => \N__25912\
        );

    \I__5363\ : Span4Mux_h
    port map (
            O => \N__25930\,
            I => \N__25903\
        );

    \I__5362\ : Span4Mux_h
    port map (
            O => \N__25927\,
            I => \N__25903\
        );

    \I__5361\ : Span4Mux_v
    port map (
            O => \N__25924\,
            I => \N__25903\
        );

    \I__5360\ : Span4Mux_v
    port map (
            O => \N__25921\,
            I => \N__25903\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__25918\,
            I => \tok.S_6\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__25915\,
            I => \tok.S_6\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__25912\,
            I => \tok.S_6\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__25903\,
            I => \tok.S_6\
        );

    \I__5355\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25889\
        );

    \I__5354\ : InMux
    port map (
            O => \N__25893\,
            I => \N__25886\
        );

    \I__5353\ : InMux
    port map (
            O => \N__25892\,
            I => \N__25883\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__25889\,
            I => \N__25879\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__25886\,
            I => \N__25876\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__25883\,
            I => \N__25872\
        );

    \I__5349\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25869\
        );

    \I__5348\ : Span4Mux_h
    port map (
            O => \N__25879\,
            I => \N__25864\
        );

    \I__5347\ : Span4Mux_v
    port map (
            O => \N__25876\,
            I => \N__25864\
        );

    \I__5346\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25861\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__25872\,
            I => \N__25858\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__25869\,
            I => \N__25855\
        );

    \I__5343\ : Span4Mux_v
    port map (
            O => \N__25864\,
            I => \N__25852\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__25861\,
            I => \N__25845\
        );

    \I__5341\ : Span4Mux_h
    port map (
            O => \N__25858\,
            I => \N__25845\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__25855\,
            I => \N__25845\
        );

    \I__5339\ : Odrv4
    port map (
            O => \N__25852\,
            I => \tok.n815\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__25845\,
            I => \tok.n815\
        );

    \I__5337\ : InMux
    port map (
            O => \N__25840\,
            I => \N__25837\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__25837\,
            I => \N__25834\
        );

    \I__5335\ : Odrv4
    port map (
            O => \N__25834\,
            I => \tok.n6510\
        );

    \I__5334\ : CascadeMux
    port map (
            O => \N__25831\,
            I => \tok.n177_adj_799_cascade_\
        );

    \I__5333\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25825\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__25825\,
            I => \N__25822\
        );

    \I__5331\ : Odrv12
    port map (
            O => \N__25822\,
            I => \tok.n127_adj_772\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__25819\,
            I => \tok.n10_adj_773_cascade_\
        );

    \I__5329\ : CascadeMux
    port map (
            O => \N__25816\,
            I => \tok.n6146_cascade_\
        );

    \I__5328\ : InMux
    port map (
            O => \N__25813\,
            I => \N__25810\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__25810\,
            I => \N__25801\
        );

    \I__5326\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25798\
        );

    \I__5325\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25794\
        );

    \I__5324\ : InMux
    port map (
            O => \N__25807\,
            I => \N__25791\
        );

    \I__5323\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25788\
        );

    \I__5322\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25785\
        );

    \I__5321\ : InMux
    port map (
            O => \N__25804\,
            I => \N__25782\
        );

    \I__5320\ : Span4Mux_h
    port map (
            O => \N__25801\,
            I => \N__25779\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__25798\,
            I => \N__25776\
        );

    \I__5318\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25773\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__25794\,
            I => \N__25768\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__25791\,
            I => \N__25768\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__25788\,
            I => \N__25763\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__25785\,
            I => \N__25763\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__25782\,
            I => \N__25756\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__25779\,
            I => \N__25756\
        );

    \I__5311\ : Span4Mux_h
    port map (
            O => \N__25776\,
            I => \N__25756\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__25773\,
            I => \N__25749\
        );

    \I__5309\ : Span4Mux_s3_v
    port map (
            O => \N__25768\,
            I => \N__25749\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__25763\,
            I => \N__25749\
        );

    \I__5307\ : Span4Mux_h
    port map (
            O => \N__25756\,
            I => \N__25746\
        );

    \I__5306\ : Span4Mux_h
    port map (
            O => \N__25749\,
            I => \N__25743\
        );

    \I__5305\ : Odrv4
    port map (
            O => \N__25746\,
            I => \tok.n86\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__25743\,
            I => \tok.n86\
        );

    \I__5303\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25734\
        );

    \I__5302\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25731\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__25734\,
            I => \N__25728\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__25731\,
            I => \N__25724\
        );

    \I__5299\ : Span4Mux_s2_h
    port map (
            O => \N__25728\,
            I => \N__25721\
        );

    \I__5298\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25718\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__25724\,
            I => \N__25715\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__25721\,
            I => \N__25712\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__25718\,
            I => \tok.n5_adj_715\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__25715\,
            I => \tok.n5_adj_715\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__25712\,
            I => \tok.n5_adj_715\
        );

    \I__5292\ : CascadeMux
    port map (
            O => \N__25705\,
            I => \tok.n369_cascade_\
        );

    \I__5291\ : InMux
    port map (
            O => \N__25702\,
            I => \N__25699\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__25699\,
            I => \N__25696\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__25696\,
            I => \N__25693\
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__25693\,
            I => \tok.n278\
        );

    \I__5287\ : CascadeMux
    port map (
            O => \N__25690\,
            I => \tok.n233_adj_716_cascade_\
        );

    \I__5286\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25684\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__25684\,
            I => \N__25681\
        );

    \I__5284\ : Span4Mux_s2_h
    port map (
            O => \N__25681\,
            I => \N__25678\
        );

    \I__5283\ : Span4Mux_v
    port map (
            O => \N__25678\,
            I => \N__25675\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__25675\,
            I => \tok.n229\
        );

    \I__5281\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25669\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__25669\,
            I => \N__25666\
        );

    \I__5279\ : Span4Mux_h
    port map (
            O => \N__25666\,
            I => \N__25663\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__25663\,
            I => \tok.n6156\
        );

    \I__5277\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25657\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__25657\,
            I => \tok.n7\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__25654\,
            I => \tok.n53_cascade_\
        );

    \I__5274\ : CEMux
    port map (
            O => \N__25651\,
            I => \N__25646\
        );

    \I__5273\ : CEMux
    port map (
            O => \N__25650\,
            I => \N__25636\
        );

    \I__5272\ : CEMux
    port map (
            O => \N__25649\,
            I => \N__25632\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__25646\,
            I => \N__25629\
        );

    \I__5270\ : CEMux
    port map (
            O => \N__25645\,
            I => \N__25626\
        );

    \I__5269\ : CEMux
    port map (
            O => \N__25644\,
            I => \N__25623\
        );

    \I__5268\ : CEMux
    port map (
            O => \N__25643\,
            I => \N__25620\
        );

    \I__5267\ : CEMux
    port map (
            O => \N__25642\,
            I => \N__25617\
        );

    \I__5266\ : CEMux
    port map (
            O => \N__25641\,
            I => \N__25614\
        );

    \I__5265\ : CEMux
    port map (
            O => \N__25640\,
            I => \N__25611\
        );

    \I__5264\ : CEMux
    port map (
            O => \N__25639\,
            I => \N__25608\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__25636\,
            I => \N__25604\
        );

    \I__5262\ : CEMux
    port map (
            O => \N__25635\,
            I => \N__25601\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__25632\,
            I => \N__25598\
        );

    \I__5260\ : Span4Mux_v
    port map (
            O => \N__25629\,
            I => \N__25593\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__25626\,
            I => \N__25593\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__25623\,
            I => \N__25590\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__25620\,
            I => \N__25587\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__25617\,
            I => \N__25584\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__25614\,
            I => \N__25577\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__25611\,
            I => \N__25577\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__25608\,
            I => \N__25577\
        );

    \I__5252\ : CEMux
    port map (
            O => \N__25607\,
            I => \N__25574\
        );

    \I__5251\ : Span4Mux_v
    port map (
            O => \N__25604\,
            I => \N__25571\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__25601\,
            I => \N__25568\
        );

    \I__5249\ : Span4Mux_h
    port map (
            O => \N__25598\,
            I => \N__25563\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__25593\,
            I => \N__25563\
        );

    \I__5247\ : Span4Mux_v
    port map (
            O => \N__25590\,
            I => \N__25560\
        );

    \I__5246\ : Span4Mux_h
    port map (
            O => \N__25587\,
            I => \N__25555\
        );

    \I__5245\ : Span4Mux_h
    port map (
            O => \N__25584\,
            I => \N__25555\
        );

    \I__5244\ : Span4Mux_v
    port map (
            O => \N__25577\,
            I => \N__25552\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__25574\,
            I => \N__25547\
        );

    \I__5242\ : Span4Mux_h
    port map (
            O => \N__25571\,
            I => \N__25547\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__25568\,
            I => \N__25544\
        );

    \I__5240\ : Span4Mux_s2_h
    port map (
            O => \N__25563\,
            I => \N__25537\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__25560\,
            I => \N__25537\
        );

    \I__5238\ : Span4Mux_h
    port map (
            O => \N__25555\,
            I => \N__25537\
        );

    \I__5237\ : Span4Mux_h
    port map (
            O => \N__25552\,
            I => \N__25532\
        );

    \I__5236\ : Span4Mux_v
    port map (
            O => \N__25547\,
            I => \N__25532\
        );

    \I__5235\ : Sp12to4
    port map (
            O => \N__25544\,
            I => \N__25527\
        );

    \I__5234\ : Sp12to4
    port map (
            O => \N__25537\,
            I => \N__25527\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__25532\,
            I => \tok.n992\
        );

    \I__5232\ : Odrv12
    port map (
            O => \N__25527\,
            I => \tok.n992\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__25522\,
            I => \tok.n2_cascade_\
        );

    \I__5230\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25512\
        );

    \I__5229\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25507\
        );

    \I__5228\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25507\
        );

    \I__5227\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25504\
        );

    \I__5226\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25501\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__25512\,
            I => \N__25494\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__25507\,
            I => \N__25494\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__25504\,
            I => \N__25489\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__25501\,
            I => \N__25489\
        );

    \I__5221\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25486\
        );

    \I__5220\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25483\
        );

    \I__5219\ : Span4Mux_v
    port map (
            O => \N__25494\,
            I => \N__25468\
        );

    \I__5218\ : Span4Mux_v
    port map (
            O => \N__25489\,
            I => \N__25468\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__25486\,
            I => \N__25468\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__25483\,
            I => \N__25468\
        );

    \I__5215\ : InMux
    port map (
            O => \N__25482\,
            I => \N__25463\
        );

    \I__5214\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25460\
        );

    \I__5213\ : InMux
    port map (
            O => \N__25480\,
            I => \N__25455\
        );

    \I__5212\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25455\
        );

    \I__5211\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25450\
        );

    \I__5210\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25450\
        );

    \I__5209\ : Span4Mux_v
    port map (
            O => \N__25468\,
            I => \N__25446\
        );

    \I__5208\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25441\
        );

    \I__5207\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25441\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__25463\,
            I => \N__25438\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__25460\,
            I => \N__25435\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__25455\,
            I => \N__25430\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__25450\,
            I => \N__25430\
        );

    \I__5202\ : InMux
    port map (
            O => \N__25449\,
            I => \N__25427\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__25446\,
            I => \N__25424\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__25441\,
            I => \N__25419\
        );

    \I__5199\ : Span4Mux_v
    port map (
            O => \N__25438\,
            I => \N__25419\
        );

    \I__5198\ : Span4Mux_h
    port map (
            O => \N__25435\,
            I => \N__25416\
        );

    \I__5197\ : Span4Mux_h
    port map (
            O => \N__25430\,
            I => \N__25413\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__25427\,
            I => \N__25410\
        );

    \I__5195\ : Sp12to4
    port map (
            O => \N__25424\,
            I => \N__25406\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__25419\,
            I => \N__25403\
        );

    \I__5193\ : Span4Mux_s1_h
    port map (
            O => \N__25416\,
            I => \N__25400\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__25413\,
            I => \N__25395\
        );

    \I__5191\ : Span4Mux_h
    port map (
            O => \N__25410\,
            I => \N__25395\
        );

    \I__5190\ : InMux
    port map (
            O => \N__25409\,
            I => \N__25392\
        );

    \I__5189\ : Odrv12
    port map (
            O => \N__25406\,
            I => \tok.n23\
        );

    \I__5188\ : Odrv4
    port map (
            O => \N__25403\,
            I => \tok.n23\
        );

    \I__5187\ : Odrv4
    port map (
            O => \N__25400\,
            I => \tok.n23\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__25395\,
            I => \tok.n23\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__25392\,
            I => \tok.n23\
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__25381\,
            I => \tok.n174_cascade_\
        );

    \I__5183\ : InMux
    port map (
            O => \N__25378\,
            I => \N__25369\
        );

    \I__5182\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25369\
        );

    \I__5181\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25364\
        );

    \I__5180\ : CascadeMux
    port map (
            O => \N__25375\,
            I => \N__25361\
        );

    \I__5179\ : CascadeMux
    port map (
            O => \N__25374\,
            I => \N__25355\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__25369\,
            I => \N__25350\
        );

    \I__5177\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25347\
        );

    \I__5176\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25344\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__25364\,
            I => \N__25340\
        );

    \I__5174\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25333\
        );

    \I__5173\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25333\
        );

    \I__5172\ : CascadeMux
    port map (
            O => \N__25359\,
            I => \N__25330\
        );

    \I__5171\ : CascadeMux
    port map (
            O => \N__25358\,
            I => \N__25326\
        );

    \I__5170\ : InMux
    port map (
            O => \N__25355\,
            I => \N__25320\
        );

    \I__5169\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25320\
        );

    \I__5168\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25317\
        );

    \I__5167\ : Span4Mux_s3_h
    port map (
            O => \N__25350\,
            I => \N__25312\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25312\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__25344\,
            I => \N__25309\
        );

    \I__5164\ : InMux
    port map (
            O => \N__25343\,
            I => \N__25306\
        );

    \I__5163\ : Span4Mux_h
    port map (
            O => \N__25340\,
            I => \N__25303\
        );

    \I__5162\ : InMux
    port map (
            O => \N__25339\,
            I => \N__25298\
        );

    \I__5161\ : InMux
    port map (
            O => \N__25338\,
            I => \N__25298\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__25333\,
            I => \N__25295\
        );

    \I__5159\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25290\
        );

    \I__5158\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25290\
        );

    \I__5157\ : InMux
    port map (
            O => \N__25326\,
            I => \N__25285\
        );

    \I__5156\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25285\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__25320\,
            I => \N__25282\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__25317\,
            I => \N__25275\
        );

    \I__5153\ : Span4Mux_h
    port map (
            O => \N__25312\,
            I => \N__25275\
        );

    \I__5152\ : Span4Mux_v
    port map (
            O => \N__25309\,
            I => \N__25275\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__25306\,
            I => \N__25270\
        );

    \I__5150\ : Span4Mux_v
    port map (
            O => \N__25303\,
            I => \N__25270\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__25298\,
            I => \tok.stall\
        );

    \I__5148\ : Odrv12
    port map (
            O => \N__25295\,
            I => \tok.stall\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__25290\,
            I => \tok.stall\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__25285\,
            I => \tok.stall\
        );

    \I__5145\ : Odrv4
    port map (
            O => \N__25282\,
            I => \tok.stall\
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__25275\,
            I => \tok.stall\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__25270\,
            I => \tok.stall\
        );

    \I__5142\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25249\
        );

    \I__5141\ : InMux
    port map (
            O => \N__25254\,
            I => \N__25249\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__25249\,
            I => \N__25244\
        );

    \I__5139\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25239\
        );

    \I__5138\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25239\
        );

    \I__5137\ : Span4Mux_v
    port map (
            O => \N__25244\,
            I => \N__25235\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__25239\,
            I => \N__25232\
        );

    \I__5135\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25229\
        );

    \I__5134\ : Sp12to4
    port map (
            O => \N__25235\,
            I => \N__25226\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__25232\,
            I => \N__25221\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__25229\,
            I => \N__25221\
        );

    \I__5131\ : Odrv12
    port map (
            O => \N__25226\,
            I => \tok.n6189\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__25221\,
            I => \tok.n6189\
        );

    \I__5129\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25213\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__25213\,
            I => \tok.n6_adj_722\
        );

    \I__5127\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25206\
        );

    \I__5126\ : InMux
    port map (
            O => \N__25209\,
            I => \N__25203\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__25206\,
            I => \N__25200\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__25203\,
            I => tail_49_adj_899
        );

    \I__5123\ : Odrv12
    port map (
            O => \N__25200\,
            I => tail_49_adj_899
        );

    \I__5122\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25189\
        );

    \I__5121\ : InMux
    port map (
            O => \N__25194\,
            I => \N__25189\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__25189\,
            I => \tok.C_stk.tail_33\
        );

    \I__5119\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25182\
        );

    \I__5118\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25179\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__25182\,
            I => \N__25176\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__25179\,
            I => tail_41
        );

    \I__5115\ : Odrv4
    port map (
            O => \N__25176\,
            I => tail_41
        );

    \I__5114\ : InMux
    port map (
            O => \N__25171\,
            I => \N__25168\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__25168\,
            I => \tok.n156\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__25165\,
            I => \tok.n211_adj_741_cascade_\
        );

    \I__5111\ : CascadeMux
    port map (
            O => \N__25162\,
            I => \tok.n277_cascade_\
        );

    \I__5110\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25156\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__25156\,
            I => \tok.n265\
        );

    \I__5108\ : InMux
    port map (
            O => \N__25153\,
            I => \N__25150\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__25150\,
            I => \N__25147\
        );

    \I__5106\ : Span4Mux_h
    port map (
            O => \N__25147\,
            I => \N__25144\
        );

    \I__5105\ : Span4Mux_h
    port map (
            O => \N__25144\,
            I => \N__25141\
        );

    \I__5104\ : Odrv4
    port map (
            O => \N__25141\,
            I => \tok.n6_adj_748\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__25138\,
            I => \N__25135\
        );

    \I__5102\ : InMux
    port map (
            O => \N__25135\,
            I => \N__25132\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__25132\,
            I => \N__25129\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__25129\,
            I => \N__25126\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__25126\,
            I => \tok.n6331\
        );

    \I__5098\ : CascadeMux
    port map (
            O => \N__25123\,
            I => \tok.n238_adj_855_cascade_\
        );

    \I__5097\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25117\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__25117\,
            I => \N__25114\
        );

    \I__5095\ : Odrv12
    port map (
            O => \N__25114\,
            I => \tok.n4_adj_859\
        );

    \I__5094\ : CascadeMux
    port map (
            O => \N__25111\,
            I => \N__25107\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__25110\,
            I => \N__25103\
        );

    \I__5092\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25100\
        );

    \I__5091\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25097\
        );

    \I__5090\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25094\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__25100\,
            I => \N__25091\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__25097\,
            I => \N__25088\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__25094\,
            I => \N__25083\
        );

    \I__5086\ : Span4Mux_s3_h
    port map (
            O => \N__25091\,
            I => \N__25083\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__25088\,
            I => \N__25080\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__25083\,
            I => \tok.n6_adj_676\
        );

    \I__5083\ : Odrv4
    port map (
            O => \N__25080\,
            I => \tok.n6_adj_676\
        );

    \I__5082\ : InMux
    port map (
            O => \N__25075\,
            I => \N__25072\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__25072\,
            I => \tok.n298_adj_856\
        );

    \I__5080\ : InMux
    port map (
            O => \N__25069\,
            I => \N__25063\
        );

    \I__5079\ : InMux
    port map (
            O => \N__25068\,
            I => \N__25063\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__25063\,
            I => \N__25060\
        );

    \I__5077\ : Span4Mux_h
    port map (
            O => \N__25060\,
            I => \N__25057\
        );

    \I__5076\ : Sp12to4
    port map (
            O => \N__25057\,
            I => \N__25054\
        );

    \I__5075\ : Odrv12
    port map (
            O => \N__25054\,
            I => \tok.n37\
        );

    \I__5074\ : InMux
    port map (
            O => \N__25051\,
            I => \N__25045\
        );

    \I__5073\ : InMux
    port map (
            O => \N__25050\,
            I => \N__25045\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__25045\,
            I => \N__25042\
        );

    \I__5071\ : Span4Mux_v
    port map (
            O => \N__25042\,
            I => \N__25039\
        );

    \I__5070\ : Sp12to4
    port map (
            O => \N__25039\,
            I => \N__25036\
        );

    \I__5069\ : Odrv12
    port map (
            O => \N__25036\,
            I => \tok.n2559\
        );

    \I__5068\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25030\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__25026\
        );

    \I__5066\ : InMux
    port map (
            O => \N__25029\,
            I => \N__25023\
        );

    \I__5065\ : Span4Mux_h
    port map (
            O => \N__25026\,
            I => \N__25018\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__25023\,
            I => \N__25018\
        );

    \I__5063\ : Odrv4
    port map (
            O => \N__25018\,
            I => \tok.tail_53\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__25015\,
            I => \rd_7__N_373_cascade_\
        );

    \I__5061\ : InMux
    port map (
            O => \N__25012\,
            I => \N__25008\
        );

    \I__5060\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25005\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__25008\,
            I => \tok.tail_61\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__25005\,
            I => \tok.tail_61\
        );

    \I__5057\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24997\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__24997\,
            I => \N__24992\
        );

    \I__5055\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24987\
        );

    \I__5054\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24987\
        );

    \I__5053\ : Span4Mux_s3_h
    port map (
            O => \N__24992\,
            I => \N__24981\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__24987\,
            I => \N__24981\
        );

    \I__5051\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24978\
        );

    \I__5050\ : Span4Mux_h
    port map (
            O => \N__24981\,
            I => \N__24975\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__24978\,
            I => tc_plus_1_1
        );

    \I__5048\ : Odrv4
    port map (
            O => \N__24975\,
            I => tc_plus_1_1
        );

    \I__5047\ : CascadeMux
    port map (
            O => \N__24970\,
            I => \tok.C_stk.n6248_cascade_\
        );

    \I__5046\ : InMux
    port map (
            O => \N__24967\,
            I => \N__24964\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__24964\,
            I => \N__24960\
        );

    \I__5044\ : InMux
    port map (
            O => \N__24963\,
            I => \N__24956\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__24960\,
            I => \N__24952\
        );

    \I__5042\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24949\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__24956\,
            I => \N__24946\
        );

    \I__5040\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24943\
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__24952\,
            I => tc_1
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__24949\,
            I => tc_1
        );

    \I__5037\ : Odrv12
    port map (
            O => \N__24946\,
            I => tc_1
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__24943\,
            I => tc_1
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__24934\,
            I => \N__24930\
        );

    \I__5034\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24921\
        );

    \I__5033\ : InMux
    port map (
            O => \N__24930\,
            I => \N__24921\
        );

    \I__5032\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24921\
        );

    \I__5031\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24918\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__24921\,
            I => \N__24915\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__24918\,
            I => c_stk_r_1
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__24915\,
            I => c_stk_r_1
        );

    \I__5027\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24904\
        );

    \I__5026\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24904\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__24904\,
            I => \tok.C_stk.tail_1\
        );

    \I__5024\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24895\
        );

    \I__5023\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24895\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__24895\,
            I => tail_9
        );

    \I__5021\ : CascadeMux
    port map (
            O => \N__24892\,
            I => \N__24889\
        );

    \I__5020\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24883\
        );

    \I__5019\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24883\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__24883\,
            I => \tok.C_stk.tail_17\
        );

    \I__5017\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24874\
        );

    \I__5016\ : InMux
    port map (
            O => \N__24879\,
            I => \N__24874\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__24874\,
            I => tail_25
        );

    \I__5014\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24867\
        );

    \I__5013\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24864\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__24867\,
            I => \N__24861\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__24864\,
            I => \tok.tail_44\
        );

    \I__5010\ : Odrv12
    port map (
            O => \N__24861\,
            I => \tok.tail_44\
        );

    \I__5009\ : InMux
    port map (
            O => \N__24856\,
            I => \N__24852\
        );

    \I__5008\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24849\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__24852\,
            I => \N__24844\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24844\
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__24844\,
            I => \tok.tail_42\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__24841\,
            I => \N__24837\
        );

    \I__5003\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24834\
        );

    \I__5002\ : InMux
    port map (
            O => \N__24837\,
            I => \N__24831\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__24834\,
            I => \N__24828\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__24831\,
            I => \N__24825\
        );

    \I__4999\ : Span4Mux_v
    port map (
            O => \N__24828\,
            I => \N__24822\
        );

    \I__4998\ : Odrv4
    port map (
            O => \N__24825\,
            I => tail_51
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__24822\,
            I => tail_51
        );

    \I__4996\ : InMux
    port map (
            O => \N__24817\,
            I => \N__24813\
        );

    \I__4995\ : InMux
    port map (
            O => \N__24816\,
            I => \N__24810\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__24813\,
            I => tail_59
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__24810\,
            I => tail_59
        );

    \I__4992\ : CascadeMux
    port map (
            O => \N__24805\,
            I => \N__24802\
        );

    \I__4991\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24798\
        );

    \I__4990\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24795\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__24798\,
            I => \N__24792\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__24795\,
            I => \N__24789\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__24792\,
            I => tail_48_adj_900
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__24789\,
            I => tail_48_adj_900
        );

    \I__4985\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24781\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__24781\,
            I => \N__24777\
        );

    \I__4983\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24774\
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__24777\,
            I => tail_56
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__24774\,
            I => tail_56
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__24769\,
            I => \C_stk_delta_1_cascade_\
        );

    \I__4979\ : InMux
    port map (
            O => \N__24766\,
            I => \N__24763\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__24763\,
            I => \N__24759\
        );

    \I__4977\ : InMux
    port map (
            O => \N__24762\,
            I => \N__24756\
        );

    \I__4976\ : Odrv12
    port map (
            O => \N__24759\,
            I => tail_57
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__24756\,
            I => tail_57
        );

    \I__4974\ : InMux
    port map (
            O => \N__24751\,
            I => \N__24747\
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__24750\,
            I => \N__24744\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__24747\,
            I => \N__24741\
        );

    \I__4971\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24738\
        );

    \I__4970\ : Odrv12
    port map (
            O => \N__24741\,
            I => \tok.tail_52\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__24738\,
            I => \tok.tail_52\
        );

    \I__4968\ : InMux
    port map (
            O => \N__24733\,
            I => \N__24729\
        );

    \I__4967\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24726\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__24729\,
            I => \tok.tail_60\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__24726\,
            I => \tok.tail_60\
        );

    \I__4964\ : InMux
    port map (
            O => \N__24721\,
            I => \N__24718\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__24718\,
            I => \N__24714\
        );

    \I__4962\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24711\
        );

    \I__4961\ : Odrv12
    port map (
            O => \N__24714\,
            I => \tok.tail_62\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__24711\,
            I => \tok.tail_62\
        );

    \I__4959\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24700\
        );

    \I__4958\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24700\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__24700\,
            I => tail_40
        );

    \I__4956\ : InMux
    port map (
            O => \N__24697\,
            I => \N__24693\
        );

    \I__4955\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24690\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__24693\,
            I => \N__24687\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__24690\,
            I => tail_8
        );

    \I__4952\ : Odrv4
    port map (
            O => \N__24687\,
            I => tail_8
        );

    \I__4951\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24678\
        );

    \I__4950\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24675\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__24678\,
            I => \tok.C_stk.tail_32\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__24675\,
            I => \tok.C_stk.tail_32\
        );

    \I__4947\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24667\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__24667\,
            I => \N__24664\
        );

    \I__4945\ : Span4Mux_h
    port map (
            O => \N__24664\,
            I => \N__24660\
        );

    \I__4944\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24657\
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__24660\,
            I => \tok.C_stk.tail_16\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__24657\,
            I => \tok.C_stk.tail_16\
        );

    \I__4941\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24648\
        );

    \I__4940\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24645\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__24648\,
            I => tail_24
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__24645\,
            I => tail_24
        );

    \I__4937\ : InMux
    port map (
            O => \N__24640\,
            I => \N__24637\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__24637\,
            I => \N__24633\
        );

    \I__4935\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24630\
        );

    \I__4934\ : Span4Mux_s3_h
    port map (
            O => \N__24633\,
            I => \N__24627\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__24630\,
            I => \tok.C_stk.tail_43\
        );

    \I__4932\ : Odrv4
    port map (
            O => \N__24627\,
            I => \tok.C_stk.tail_43\
        );

    \I__4931\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24619\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__24619\,
            I => \N__24615\
        );

    \I__4929\ : InMux
    port map (
            O => \N__24618\,
            I => \N__24612\
        );

    \I__4928\ : Span4Mux_s3_h
    port map (
            O => \N__24615\,
            I => \N__24609\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__24612\,
            I => \tok.tail_45\
        );

    \I__4926\ : Odrv4
    port map (
            O => \N__24609\,
            I => \tok.tail_45\
        );

    \I__4925\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24601\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__24601\,
            I => \tok.n6442\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__24598\,
            I => \tok.n6433_cascade_\
        );

    \I__4922\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24592\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__24592\,
            I => \N__24589\
        );

    \I__4920\ : Span4Mux_h
    port map (
            O => \N__24589\,
            I => \N__24586\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__24586\,
            I => \tok.n215_adj_841\
        );

    \I__4918\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24580\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__24580\,
            I => \tok.n179_adj_842\
        );

    \I__4916\ : CascadeMux
    port map (
            O => \N__24577\,
            I => \tok.n6602_cascade_\
        );

    \I__4915\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24571\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__24571\,
            I => \N__24568\
        );

    \I__4913\ : Odrv4
    port map (
            O => \N__24568\,
            I => \tok.n6601\
        );

    \I__4912\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24562\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__24562\,
            I => \N__24559\
        );

    \I__4910\ : Odrv4
    port map (
            O => \N__24559\,
            I => \tok.n6375\
        );

    \I__4909\ : InMux
    port map (
            O => \N__24556\,
            I => \N__24548\
        );

    \I__4908\ : CascadeMux
    port map (
            O => \N__24555\,
            I => \N__24545\
        );

    \I__4907\ : CascadeMux
    port map (
            O => \N__24554\,
            I => \N__24542\
        );

    \I__4906\ : CascadeMux
    port map (
            O => \N__24553\,
            I => \N__24537\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__24552\,
            I => \N__24534\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__24551\,
            I => \N__24531\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__24548\,
            I => \N__24528\
        );

    \I__4902\ : InMux
    port map (
            O => \N__24545\,
            I => \N__24525\
        );

    \I__4901\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24518\
        );

    \I__4900\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24518\
        );

    \I__4899\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24518\
        );

    \I__4898\ : InMux
    port map (
            O => \N__24537\,
            I => \N__24515\
        );

    \I__4897\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24512\
        );

    \I__4896\ : InMux
    port map (
            O => \N__24531\,
            I => \N__24509\
        );

    \I__4895\ : Span4Mux_v
    port map (
            O => \N__24528\,
            I => \N__24502\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__24525\,
            I => \N__24502\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24502\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__24515\,
            I => \tok.n847\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__24512\,
            I => \tok.n847\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__24509\,
            I => \tok.n847\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__24502\,
            I => \tok.n847\
        );

    \I__4888\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24490\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__24490\,
            I => \tok.n6544\
        );

    \I__4886\ : CascadeMux
    port map (
            O => \N__24487\,
            I => \tok.n179_adj_657_cascade_\
        );

    \I__4885\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24481\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__24481\,
            I => \N__24478\
        );

    \I__4883\ : Span4Mux_h
    port map (
            O => \N__24478\,
            I => \N__24475\
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__24475\,
            I => \tok.n6543\
        );

    \I__4881\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24469\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__24469\,
            I => \N__24466\
        );

    \I__4879\ : Odrv12
    port map (
            O => \N__24466\,
            I => \tok.n464\
        );

    \I__4878\ : CascadeMux
    port map (
            O => \N__24463\,
            I => \N__24455\
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__24462\,
            I => \N__24449\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__24461\,
            I => \N__24445\
        );

    \I__4875\ : CascadeMux
    port map (
            O => \N__24460\,
            I => \N__24442\
        );

    \I__4874\ : CascadeMux
    port map (
            O => \N__24459\,
            I => \N__24438\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__24458\,
            I => \N__24434\
        );

    \I__4872\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24430\
        );

    \I__4871\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24427\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__24453\,
            I => \N__24422\
        );

    \I__4869\ : InMux
    port map (
            O => \N__24452\,
            I => \N__24413\
        );

    \I__4868\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24413\
        );

    \I__4867\ : InMux
    port map (
            O => \N__24448\,
            I => \N__24413\
        );

    \I__4866\ : InMux
    port map (
            O => \N__24445\,
            I => \N__24413\
        );

    \I__4865\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24410\
        );

    \I__4864\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24405\
        );

    \I__4863\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24405\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__24437\,
            I => \N__24402\
        );

    \I__4861\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24399\
        );

    \I__4860\ : CascadeMux
    port map (
            O => \N__24433\,
            I => \N__24396\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__24430\,
            I => \N__24391\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__24427\,
            I => \N__24391\
        );

    \I__4857\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24384\
        );

    \I__4856\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24384\
        );

    \I__4855\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24384\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__24413\,
            I => \N__24379\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__24410\,
            I => \N__24379\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__24405\,
            I => \N__24376\
        );

    \I__4851\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24373\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__24399\,
            I => \N__24370\
        );

    \I__4849\ : InMux
    port map (
            O => \N__24396\,
            I => \N__24367\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__24391\,
            I => \N__24362\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__24384\,
            I => \N__24362\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__24379\,
            I => \N__24359\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__24376\,
            I => \N__24356\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__24373\,
            I => \tok.n8\
        );

    \I__4843\ : Odrv4
    port map (
            O => \N__24370\,
            I => \tok.n8\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__24367\,
            I => \tok.n8\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__24362\,
            I => \tok.n8\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__24359\,
            I => \tok.n8\
        );

    \I__4839\ : Odrv4
    port map (
            O => \N__24356\,
            I => \tok.n8\
        );

    \I__4838\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24340\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__24340\,
            I => \tok.n6382\
        );

    \I__4836\ : CascadeMux
    port map (
            O => \N__24337\,
            I => \N__24334\
        );

    \I__4835\ : InMux
    port map (
            O => \N__24334\,
            I => \N__24330\
        );

    \I__4834\ : InMux
    port map (
            O => \N__24333\,
            I => \N__24325\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__24330\,
            I => \N__24319\
        );

    \I__4832\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24314\
        );

    \I__4831\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24311\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__24325\,
            I => \N__24308\
        );

    \I__4829\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24305\
        );

    \I__4828\ : InMux
    port map (
            O => \N__24323\,
            I => \N__24300\
        );

    \I__4827\ : InMux
    port map (
            O => \N__24322\,
            I => \N__24300\
        );

    \I__4826\ : Span4Mux_v
    port map (
            O => \N__24319\,
            I => \N__24297\
        );

    \I__4825\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24294\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__24317\,
            I => \N__24291\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24284\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__24311\,
            I => \N__24279\
        );

    \I__4821\ : Span4Mux_v
    port map (
            O => \N__24308\,
            I => \N__24279\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24274\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__24300\,
            I => \N__24274\
        );

    \I__4818\ : Sp12to4
    port map (
            O => \N__24297\,
            I => \N__24269\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__24294\,
            I => \N__24269\
        );

    \I__4816\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24266\
        );

    \I__4815\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24259\
        );

    \I__4814\ : InMux
    port map (
            O => \N__24289\,
            I => \N__24259\
        );

    \I__4813\ : InMux
    port map (
            O => \N__24288\,
            I => \N__24259\
        );

    \I__4812\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24256\
        );

    \I__4811\ : Span4Mux_s2_v
    port map (
            O => \N__24284\,
            I => \N__24249\
        );

    \I__4810\ : Span4Mux_s2_v
    port map (
            O => \N__24279\,
            I => \N__24249\
        );

    \I__4809\ : Span4Mux_v
    port map (
            O => \N__24274\,
            I => \N__24249\
        );

    \I__4808\ : Span12Mux_h
    port map (
            O => \N__24269\,
            I => \N__24246\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__24266\,
            I => \N__24237\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__24259\,
            I => \N__24237\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__24256\,
            I => \N__24237\
        );

    \I__4804\ : Sp12to4
    port map (
            O => \N__24249\,
            I => \N__24237\
        );

    \I__4803\ : Odrv12
    port map (
            O => \N__24246\,
            I => \tok.n4_adj_636\
        );

    \I__4802\ : Odrv12
    port map (
            O => \N__24237\,
            I => \tok.n4_adj_636\
        );

    \I__4801\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24229\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__24229\,
            I => \tok.n213_adj_795\
        );

    \I__4799\ : CascadeMux
    port map (
            O => \N__24226\,
            I => \tok.n207_adj_796_cascade_\
        );

    \I__4798\ : InMux
    port map (
            O => \N__24223\,
            I => \N__24220\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__24220\,
            I => \N__24215\
        );

    \I__4796\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24210\
        );

    \I__4795\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24210\
        );

    \I__4794\ : Span4Mux_s3_v
    port map (
            O => \N__24215\,
            I => \N__24205\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__24210\,
            I => \N__24205\
        );

    \I__4792\ : Odrv4
    port map (
            O => \N__24205\,
            I => \tok.n872\
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__24202\,
            I => \tok.n6505_cascade_\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__24199\,
            I => \N__24193\
        );

    \I__4789\ : InMux
    port map (
            O => \N__24198\,
            I => \N__24190\
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__24197\,
            I => \N__24187\
        );

    \I__4787\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24181\
        );

    \I__4786\ : InMux
    port map (
            O => \N__24193\,
            I => \N__24176\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__24190\,
            I => \N__24173\
        );

    \I__4784\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24170\
        );

    \I__4783\ : InMux
    port map (
            O => \N__24186\,
            I => \N__24166\
        );

    \I__4782\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24161\
        );

    \I__4781\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24161\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__24181\,
            I => \N__24158\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__24180\,
            I => \N__24155\
        );

    \I__4778\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24152\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24149\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__24173\,
            I => \N__24144\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__24170\,
            I => \N__24144\
        );

    \I__4774\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24140\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__24166\,
            I => \N__24137\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__24161\,
            I => \N__24134\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__24158\,
            I => \N__24130\
        );

    \I__4770\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24127\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__24152\,
            I => \N__24124\
        );

    \I__4768\ : Span4Mux_v
    port map (
            O => \N__24149\,
            I => \N__24119\
        );

    \I__4767\ : Span4Mux_s1_h
    port map (
            O => \N__24144\,
            I => \N__24119\
        );

    \I__4766\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24116\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__24140\,
            I => \N__24113\
        );

    \I__4764\ : Span4Mux_h
    port map (
            O => \N__24137\,
            I => \N__24108\
        );

    \I__4763\ : Span4Mux_h
    port map (
            O => \N__24134\,
            I => \N__24108\
        );

    \I__4762\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24105\
        );

    \I__4761\ : Span4Mux_v
    port map (
            O => \N__24130\,
            I => \N__24102\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N__24099\
        );

    \I__4759\ : Span4Mux_h
    port map (
            O => \N__24124\,
            I => \N__24094\
        );

    \I__4758\ : Span4Mux_h
    port map (
            O => \N__24119\,
            I => \N__24094\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__24116\,
            I => \N__24091\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__24113\,
            I => \N__24086\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__24108\,
            I => \N__24086\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__24105\,
            I => \tok.n42\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__24102\,
            I => \tok.n42\
        );

    \I__4752\ : Odrv12
    port map (
            O => \N__24099\,
            I => \tok.n42\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__24094\,
            I => \tok.n42\
        );

    \I__4750\ : Odrv12
    port map (
            O => \N__24091\,
            I => \tok.n42\
        );

    \I__4749\ : Odrv4
    port map (
            O => \N__24086\,
            I => \tok.n42\
        );

    \I__4748\ : InMux
    port map (
            O => \N__24073\,
            I => \N__24070\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__24070\,
            I => \N__24067\
        );

    \I__4746\ : Span4Mux_s2_v
    port map (
            O => \N__24067\,
            I => \N__24064\
        );

    \I__4745\ : Odrv4
    port map (
            O => \N__24064\,
            I => \tok.n6360\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__24061\,
            I => \N__24057\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__24060\,
            I => \N__24054\
        );

    \I__4742\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24051\
        );

    \I__4741\ : InMux
    port map (
            O => \N__24054\,
            I => \N__24048\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__24051\,
            I => \N__24045\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24042\
        );

    \I__4738\ : Span4Mux_v
    port map (
            O => \N__24045\,
            I => \N__24039\
        );

    \I__4737\ : Span4Mux_v
    port map (
            O => \N__24042\,
            I => \N__24036\
        );

    \I__4736\ : Span4Mux_h
    port map (
            O => \N__24039\,
            I => \N__24031\
        );

    \I__4735\ : Span4Mux_v
    port map (
            O => \N__24036\,
            I => \N__24031\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__24031\,
            I => \tok.table_rd_6\
        );

    \I__4733\ : InMux
    port map (
            O => \N__24028\,
            I => \N__24025\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__24025\,
            I => \N__24022\
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__24022\,
            I => \tok.n210_adj_802\
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__24019\,
            I => \N__24016\
        );

    \I__4729\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24013\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__24013\,
            I => \N__24010\
        );

    \I__4727\ : Span4Mux_h
    port map (
            O => \N__24010\,
            I => \N__24007\
        );

    \I__4726\ : Odrv4
    port map (
            O => \N__24007\,
            I => \tok.n316\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__24004\,
            I => \tok.n6409_cascade_\
        );

    \I__4724\ : InMux
    port map (
            O => \N__24001\,
            I => \N__23996\
        );

    \I__4723\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23989\
        );

    \I__4722\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23984\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__23996\,
            I => \N__23981\
        );

    \I__4720\ : InMux
    port map (
            O => \N__23995\,
            I => \N__23978\
        );

    \I__4719\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23975\
        );

    \I__4718\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23972\
        );

    \I__4717\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23969\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__23989\,
            I => \N__23962\
        );

    \I__4715\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23957\
        );

    \I__4714\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23957\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__23984\,
            I => \N__23954\
        );

    \I__4712\ : Span4Mux_v
    port map (
            O => \N__23981\,
            I => \N__23945\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__23978\,
            I => \N__23945\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__23975\,
            I => \N__23945\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__23972\,
            I => \N__23942\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__23969\,
            I => \N__23939\
        );

    \I__4707\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23936\
        );

    \I__4706\ : InMux
    port map (
            O => \N__23967\,
            I => \N__23929\
        );

    \I__4705\ : InMux
    port map (
            O => \N__23966\,
            I => \N__23929\
        );

    \I__4704\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23929\
        );

    \I__4703\ : Span12Mux_v
    port map (
            O => \N__23962\,
            I => \N__23926\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__23957\,
            I => \N__23921\
        );

    \I__4701\ : Span4Mux_v
    port map (
            O => \N__23954\,
            I => \N__23921\
        );

    \I__4700\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23916\
        );

    \I__4699\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23916\
        );

    \I__4698\ : Span4Mux_v
    port map (
            O => \N__23945\,
            I => \N__23913\
        );

    \I__4697\ : Span4Mux_v
    port map (
            O => \N__23942\,
            I => \N__23906\
        );

    \I__4696\ : Span4Mux_h
    port map (
            O => \N__23939\,
            I => \N__23906\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__23936\,
            I => \N__23906\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__23929\,
            I => \N__23903\
        );

    \I__4693\ : Odrv12
    port map (
            O => \N__23926\,
            I => \tok.n46\
        );

    \I__4692\ : Odrv4
    port map (
            O => \N__23921\,
            I => \tok.n46\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__23916\,
            I => \tok.n46\
        );

    \I__4690\ : Odrv4
    port map (
            O => \N__23913\,
            I => \tok.n46\
        );

    \I__4689\ : Odrv4
    port map (
            O => \N__23906\,
            I => \tok.n46\
        );

    \I__4688\ : Odrv12
    port map (
            O => \N__23903\,
            I => \tok.n46\
        );

    \I__4687\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23887\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__23887\,
            I => \N__23884\
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__23884\,
            I => \tok.n215_adj_887\
        );

    \I__4684\ : CascadeMux
    port map (
            O => \N__23881\,
            I => \tok.n207_adj_811_cascade_\
        );

    \I__4683\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23875\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__23875\,
            I => \tok.n6481\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__23872\,
            I => \N__23869\
        );

    \I__4680\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23866\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__23866\,
            I => \tok.n6484\
        );

    \I__4678\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23860\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__23860\,
            I => \tok.n213_adj_810\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__23857\,
            I => \N__23853\
        );

    \I__4675\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23848\
        );

    \I__4674\ : InMux
    port map (
            O => \N__23853\,
            I => \N__23845\
        );

    \I__4673\ : CascadeMux
    port map (
            O => \N__23852\,
            I => \N__23840\
        );

    \I__4672\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23836\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__23848\,
            I => \N__23831\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__23845\,
            I => \N__23831\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__23844\,
            I => \N__23828\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__23843\,
            I => \N__23825\
        );

    \I__4667\ : InMux
    port map (
            O => \N__23840\,
            I => \N__23822\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__23839\,
            I => \N__23819\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__23836\,
            I => \N__23816\
        );

    \I__4664\ : Span4Mux_v
    port map (
            O => \N__23831\,
            I => \N__23813\
        );

    \I__4663\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23810\
        );

    \I__4662\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23807\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__23822\,
            I => \N__23804\
        );

    \I__4660\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23801\
        );

    \I__4659\ : Span4Mux_s3_v
    port map (
            O => \N__23816\,
            I => \N__23797\
        );

    \I__4658\ : Span4Mux_h
    port map (
            O => \N__23813\,
            I => \N__23790\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__23810\,
            I => \N__23790\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__23807\,
            I => \N__23790\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__23804\,
            I => \N__23785\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__23801\,
            I => \N__23785\
        );

    \I__4653\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23782\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__23797\,
            I => \N__23777\
        );

    \I__4651\ : Span4Mux_h
    port map (
            O => \N__23790\,
            I => \N__23777\
        );

    \I__4650\ : Span4Mux_h
    port map (
            O => \N__23785\,
            I => \N__23774\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__23782\,
            I => \tok.S_4\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__23777\,
            I => \tok.S_4\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__23774\,
            I => \tok.S_4\
        );

    \I__4646\ : CascadeMux
    port map (
            O => \N__23767\,
            I => \tok.n207_cascade_\
        );

    \I__4645\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23761\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__23761\,
            I => \N__23758\
        );

    \I__4643\ : Odrv4
    port map (
            O => \N__23758\,
            I => \tok.n210\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__23755\,
            I => \tok.n6572_cascade_\
        );

    \I__4641\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23749\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__23749\,
            I => \tok.n174_adj_768\
        );

    \I__4639\ : CascadeMux
    port map (
            O => \N__23746\,
            I => \N__23743\
        );

    \I__4638\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23738\
        );

    \I__4637\ : InMux
    port map (
            O => \N__23742\,
            I => \N__23733\
        );

    \I__4636\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23733\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__23738\,
            I => \N__23721\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__23733\,
            I => \N__23721\
        );

    \I__4633\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23716\
        );

    \I__4632\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23711\
        );

    \I__4631\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23711\
        );

    \I__4630\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23706\
        );

    \I__4629\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23706\
        );

    \I__4628\ : InMux
    port map (
            O => \N__23727\,
            I => \N__23701\
        );

    \I__4627\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23701\
        );

    \I__4626\ : Span4Mux_h
    port map (
            O => \N__23721\,
            I => \N__23698\
        );

    \I__4625\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23693\
        );

    \I__4624\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23693\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__23716\,
            I => \N__23690\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__23711\,
            I => \tok.n31\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__23706\,
            I => \tok.n31\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__23701\,
            I => \tok.n31\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__23698\,
            I => \tok.n31\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__23693\,
            I => \tok.n31\
        );

    \I__4617\ : Odrv12
    port map (
            O => \N__23690\,
            I => \tok.n31\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__23677\,
            I => \N__23672\
        );

    \I__4615\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23669\
        );

    \I__4614\ : InMux
    port map (
            O => \N__23675\,
            I => \N__23666\
        );

    \I__4613\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23663\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__23669\,
            I => \tok.n26_adj_763\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__23666\,
            I => \tok.n26_adj_763\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__23663\,
            I => \tok.n26_adj_763\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__23656\,
            I => \tok.n26_adj_763_cascade_\
        );

    \I__4608\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23650\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23647\
        );

    \I__4606\ : Span4Mux_v
    port map (
            O => \N__23647\,
            I => \N__23644\
        );

    \I__4605\ : Sp12to4
    port map (
            O => \N__23644\,
            I => \N__23641\
        );

    \I__4604\ : Odrv12
    port map (
            O => \N__23641\,
            I => \tok.n6466\
        );

    \I__4603\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23635\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__23635\,
            I => \N__23632\
        );

    \I__4601\ : Odrv12
    port map (
            O => \N__23632\,
            I => \tok.n6467\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__23629\,
            I => \N__23626\
        );

    \I__4599\ : InMux
    port map (
            O => \N__23626\,
            I => \N__23623\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__23623\,
            I => \N__23620\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__23620\,
            I => \tok.n6486\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__23617\,
            I => \N__23613\
        );

    \I__4595\ : InMux
    port map (
            O => \N__23616\,
            I => \N__23609\
        );

    \I__4594\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23606\
        );

    \I__4593\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23603\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__23609\,
            I => \N__23600\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__23606\,
            I => \N__23597\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23594\
        );

    \I__4589\ : Span4Mux_h
    port map (
            O => \N__23600\,
            I => \N__23591\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__23597\,
            I => \N__23586\
        );

    \I__4587\ : Span4Mux_v
    port map (
            O => \N__23594\,
            I => \N__23586\
        );

    \I__4586\ : Odrv4
    port map (
            O => \N__23591\,
            I => \tok.n833\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__23586\,
            I => \tok.n833\
        );

    \I__4584\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23578\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__23578\,
            I => \N__23575\
        );

    \I__4582\ : Span4Mux_h
    port map (
            O => \N__23575\,
            I => \N__23572\
        );

    \I__4581\ : Odrv4
    port map (
            O => \N__23572\,
            I => \tok.n6490\
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__23569\,
            I => \N__23566\
        );

    \I__4579\ : InMux
    port map (
            O => \N__23566\,
            I => \N__23563\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__23563\,
            I => \N__23560\
        );

    \I__4577\ : Span4Mux_h
    port map (
            O => \N__23560\,
            I => \N__23557\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__23557\,
            I => \tok.n6491\
        );

    \I__4575\ : CascadeMux
    port map (
            O => \N__23554\,
            I => \N__23550\
        );

    \I__4574\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23543\
        );

    \I__4573\ : InMux
    port map (
            O => \N__23550\,
            I => \N__23540\
        );

    \I__4572\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23537\
        );

    \I__4571\ : InMux
    port map (
            O => \N__23548\,
            I => \N__23534\
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__23547\,
            I => \N__23531\
        );

    \I__4569\ : CascadeMux
    port map (
            O => \N__23546\,
            I => \N__23528\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__23543\,
            I => \N__23525\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__23540\,
            I => \N__23520\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__23537\,
            I => \N__23520\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23517\
        );

    \I__4564\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23514\
        );

    \I__4563\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23511\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__23525\,
            I => \N__23506\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__23520\,
            I => \N__23506\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__23517\,
            I => \N__23503\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23500\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__23511\,
            I => \N__23497\
        );

    \I__4557\ : Span4Mux_h
    port map (
            O => \N__23506\,
            I => \N__23486\
        );

    \I__4556\ : Span4Mux_h
    port map (
            O => \N__23503\,
            I => \N__23486\
        );

    \I__4555\ : Span4Mux_v
    port map (
            O => \N__23500\,
            I => \N__23486\
        );

    \I__4554\ : Span4Mux_v
    port map (
            O => \N__23497\,
            I => \N__23486\
        );

    \I__4553\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23483\
        );

    \I__4552\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23480\
        );

    \I__4551\ : Span4Mux_v
    port map (
            O => \N__23486\,
            I => \N__23477\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__23483\,
            I => \S_1\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__23480\,
            I => \S_1\
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__23477\,
            I => \S_1\
        );

    \I__4547\ : InMux
    port map (
            O => \N__23470\,
            I => \N__23467\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__23467\,
            I => \N__23464\
        );

    \I__4545\ : Span4Mux_h
    port map (
            O => \N__23464\,
            I => \N__23461\
        );

    \I__4544\ : Odrv4
    port map (
            O => \N__23461\,
            I => \tok.n208\
        );

    \I__4543\ : CascadeMux
    port map (
            O => \N__23458\,
            I => \N__23455\
        );

    \I__4542\ : InMux
    port map (
            O => \N__23455\,
            I => \N__23452\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__23452\,
            I => \N__23449\
        );

    \I__4540\ : Span4Mux_h
    port map (
            O => \N__23449\,
            I => \N__23446\
        );

    \I__4539\ : Span4Mux_s3_h
    port map (
            O => \N__23446\,
            I => \N__23443\
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__23443\,
            I => \tok.n6589\
        );

    \I__4537\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23437\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__23437\,
            I => \N__23434\
        );

    \I__4535\ : Span12Mux_s6_h
    port map (
            O => \N__23434\,
            I => \N__23431\
        );

    \I__4534\ : Odrv12
    port map (
            O => \N__23431\,
            I => \tok.n239_adj_727\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__23428\,
            I => \tok.n6_adj_728_cascade_\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__23425\,
            I => \tok.n200_adj_732_cascade_\
        );

    \I__4531\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23419\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23416\
        );

    \I__4529\ : Odrv12
    port map (
            O => \N__23416\,
            I => \tok.n203_adj_731\
        );

    \I__4528\ : InMux
    port map (
            O => \N__23413\,
            I => \N__23410\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__23410\,
            I => \N__23407\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__23407\,
            I => \N__23404\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__23404\,
            I => \tok.n6_adj_733\
        );

    \I__4524\ : InMux
    port map (
            O => \N__23401\,
            I => \N__23397\
        );

    \I__4523\ : InMux
    port map (
            O => \N__23400\,
            I => \N__23394\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__23397\,
            I => \N__23389\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23389\
        );

    \I__4520\ : Span4Mux_v
    port map (
            O => \N__23389\,
            I => \N__23386\
        );

    \I__4519\ : Span4Mux_v
    port map (
            O => \N__23386\,
            I => \N__23383\
        );

    \I__4518\ : Odrv4
    port map (
            O => \N__23383\,
            I => \tok.n206_adj_794\
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__23380\,
            I => \tok.n244_cascade_\
        );

    \I__4516\ : CascadeMux
    port map (
            O => \N__23377\,
            I => \tok.n4_adj_720_cascade_\
        );

    \I__4515\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23371\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__23371\,
            I => \N__23368\
        );

    \I__4513\ : Odrv12
    port map (
            O => \N__23368\,
            I => \tok.n145\
        );

    \I__4512\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23362\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__23362\,
            I => \tok.n251\
        );

    \I__4510\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23356\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__23356\,
            I => \N__23352\
        );

    \I__4508\ : InMux
    port map (
            O => \N__23355\,
            I => \N__23349\
        );

    \I__4507\ : Span4Mux_h
    port map (
            O => \N__23352\,
            I => \N__23346\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__23349\,
            I => \N__23343\
        );

    \I__4505\ : Span4Mux_v
    port map (
            O => \N__23346\,
            I => \N__23340\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__23343\,
            I => \N__23337\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__23340\,
            I => \tok.n2557\
        );

    \I__4502\ : Odrv4
    port map (
            O => \N__23337\,
            I => \tok.n2557\
        );

    \I__4501\ : CascadeMux
    port map (
            O => \N__23332\,
            I => \tok.n4_adj_714_cascade_\
        );

    \I__4500\ : InMux
    port map (
            O => \N__23329\,
            I => \N__23326\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__23326\,
            I => \tok.n218\
        );

    \I__4498\ : InMux
    port map (
            O => \N__23323\,
            I => \N__23320\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__23320\,
            I => \tok.n39\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__23317\,
            I => \tok.n6269_cascade_\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__23314\,
            I => \tok.n197_adj_729_cascade_\
        );

    \I__4494\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23308\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__23308\,
            I => \N__23305\
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__23305\,
            I => \tok.n7458\
        );

    \I__4491\ : InMux
    port map (
            O => \N__23302\,
            I => \N__23299\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__23299\,
            I => \tok.n2544\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__23296\,
            I => \N__23292\
        );

    \I__4488\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23289\
        );

    \I__4487\ : InMux
    port map (
            O => \N__23292\,
            I => \N__23286\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__23289\,
            I => \N__23283\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__23286\,
            I => \N__23280\
        );

    \I__4484\ : Span4Mux_v
    port map (
            O => \N__23283\,
            I => \N__23277\
        );

    \I__4483\ : Sp12to4
    port map (
            O => \N__23280\,
            I => \N__23274\
        );

    \I__4482\ : Span4Mux_h
    port map (
            O => \N__23277\,
            I => \N__23271\
        );

    \I__4481\ : Span12Mux_s10_h
    port map (
            O => \N__23274\,
            I => \N__23268\
        );

    \I__4480\ : Odrv4
    port map (
            O => \N__23271\,
            I => \tok.table_rd_1\
        );

    \I__4479\ : Odrv12
    port map (
            O => \N__23268\,
            I => \tok.table_rd_1\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__23263\,
            I => \tok.n7475_cascade_\
        );

    \I__4477\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23256\
        );

    \I__4476\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23253\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__23256\,
            I => \N__23248\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__23253\,
            I => \N__23248\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__23248\,
            I => \N__23245\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__23245\,
            I => \N__23242\
        );

    \I__4471\ : Odrv4
    port map (
            O => \N__23242\,
            I => \tok.n237\
        );

    \I__4470\ : CascadeMux
    port map (
            O => \N__23239\,
            I => \N__23236\
        );

    \I__4469\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23233\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__23233\,
            I => \N__23230\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__23230\,
            I => \tok.n180\
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__23227\,
            I => \N__23224\
        );

    \I__4465\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23221\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__23221\,
            I => \tok.n6628\
        );

    \I__4463\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23212\
        );

    \I__4462\ : InMux
    port map (
            O => \N__23217\,
            I => \N__23206\
        );

    \I__4461\ : InMux
    port map (
            O => \N__23216\,
            I => \N__23203\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__23215\,
            I => \N__23200\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__23212\,
            I => \N__23197\
        );

    \I__4458\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23194\
        );

    \I__4457\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23191\
        );

    \I__4456\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23188\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__23206\,
            I => \N__23185\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__23203\,
            I => \N__23182\
        );

    \I__4453\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23179\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__23197\,
            I => \N__23173\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__23194\,
            I => \N__23173\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__23191\,
            I => \N__23170\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__23188\,
            I => \N__23161\
        );

    \I__4448\ : Span4Mux_h
    port map (
            O => \N__23185\,
            I => \N__23161\
        );

    \I__4447\ : Span4Mux_v
    port map (
            O => \N__23182\,
            I => \N__23161\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__23179\,
            I => \N__23161\
        );

    \I__4445\ : InMux
    port map (
            O => \N__23178\,
            I => \N__23158\
        );

    \I__4444\ : Span4Mux_v
    port map (
            O => \N__23173\,
            I => \N__23155\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__23170\,
            I => \N__23150\
        );

    \I__4442\ : Span4Mux_h
    port map (
            O => \N__23161\,
            I => \N__23150\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__23158\,
            I => \tok.S_3\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__23155\,
            I => \tok.S_3\
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__23150\,
            I => \tok.S_3\
        );

    \I__4438\ : CascadeMux
    port map (
            O => \N__23143\,
            I => \N__23140\
        );

    \I__4437\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23137\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__23137\,
            I => \N__23134\
        );

    \I__4435\ : Odrv4
    port map (
            O => \N__23134\,
            I => \tok.n241\
        );

    \I__4434\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23128\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__23128\,
            I => \N__23125\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__23125\,
            I => \tok.n6637\
        );

    \I__4431\ : CascadeMux
    port map (
            O => \N__23122\,
            I => \tok.n284_cascade_\
        );

    \I__4430\ : InMux
    port map (
            O => \N__23119\,
            I => \N__23116\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__23116\,
            I => \tok.n17\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__23113\,
            I => \N__23110\
        );

    \I__4427\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23107\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__23107\,
            I => \N__23103\
        );

    \I__4425\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23100\
        );

    \I__4424\ : Span12Mux_s9_h
    port map (
            O => \N__23103\,
            I => \N__23097\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__23100\,
            I => \tok.n5_adj_821\
        );

    \I__4422\ : Odrv12
    port map (
            O => \N__23097\,
            I => \tok.n5_adj_821\
        );

    \I__4421\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23089\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__23089\,
            I => \tok.n2679\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__23086\,
            I => \tok.n17_cascade_\
        );

    \I__4418\ : CascadeMux
    port map (
            O => \N__23083\,
            I => \N__23080\
        );

    \I__4417\ : InMux
    port map (
            O => \N__23080\,
            I => \N__23077\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__23077\,
            I => \tok.n864\
        );

    \I__4415\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__23071\,
            I => \N__23068\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__23068\,
            I => \tok.n186\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__23065\,
            I => \tok.n6562_cascade_\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__23062\,
            I => \N__23059\
        );

    \I__4410\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23056\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__23056\,
            I => \N__23053\
        );

    \I__4408\ : Span4Mux_v
    port map (
            O => \N__23053\,
            I => \N__23050\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__23050\,
            I => \tok.n338\
        );

    \I__4406\ : InMux
    port map (
            O => \N__23047\,
            I => \N__23044\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__23044\,
            I => \tok.n162\
        );

    \I__4404\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23038\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__23038\,
            I => \tok.n179_adj_730\
        );

    \I__4402\ : InMux
    port map (
            O => \N__23035\,
            I => \N__23032\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__23032\,
            I => \N__23029\
        );

    \I__4400\ : Span4Mux_v
    port map (
            O => \N__23029\,
            I => \N__23026\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__23026\,
            I => \tok.n4926\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__23023\,
            I => \tok.n2692_cascade_\
        );

    \I__4397\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23017\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__23014\
        );

    \I__4395\ : Span4Mux_h
    port map (
            O => \N__23014\,
            I => \N__23011\
        );

    \I__4394\ : Odrv4
    port map (
            O => \N__23011\,
            I => \tok.n217\
        );

    \I__4393\ : InMux
    port map (
            O => \N__23008\,
            I => \N__23005\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__23005\,
            I => \tok.n7154\
        );

    \I__4391\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22999\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__22999\,
            I => \tok.n6_adj_701\
        );

    \I__4389\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22993\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__22993\,
            I => \tok.n2700\
        );

    \I__4387\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__22987\,
            I => \tok.n236_adj_737\
        );

    \I__4385\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22981\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__22981\,
            I => \N__22978\
        );

    \I__4383\ : Span4Mux_h
    port map (
            O => \N__22978\,
            I => \N__22975\
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__22975\,
            I => \tok.n239_adj_738\
        );

    \I__4381\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22966\
        );

    \I__4380\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22966\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__22966\,
            I => \tok.C_stk.tail_19\
        );

    \I__4378\ : InMux
    port map (
            O => \N__22963\,
            I => \N__22957\
        );

    \I__4377\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22957\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__22957\,
            I => \tok.C_stk.tail_27\
        );

    \I__4375\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22948\
        );

    \I__4374\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22948\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__22948\,
            I => \tok.C_stk.tail_35\
        );

    \I__4372\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22940\
        );

    \I__4371\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22936\
        );

    \I__4370\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22933\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__22940\,
            I => \N__22928\
        );

    \I__4368\ : InMux
    port map (
            O => \N__22939\,
            I => \N__22925\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__22936\,
            I => \N__22922\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__22933\,
            I => \N__22919\
        );

    \I__4365\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22916\
        );

    \I__4364\ : InMux
    port map (
            O => \N__22931\,
            I => \N__22911\
        );

    \I__4363\ : Span4Mux_v
    port map (
            O => \N__22928\,
            I => \N__22906\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__22925\,
            I => \N__22906\
        );

    \I__4361\ : Span4Mux_v
    port map (
            O => \N__22922\,
            I => \N__22903\
        );

    \I__4360\ : Span4Mux_v
    port map (
            O => \N__22919\,
            I => \N__22898\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22898\
        );

    \I__4358\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22895\
        );

    \I__4357\ : InMux
    port map (
            O => \N__22914\,
            I => \N__22892\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__22911\,
            I => \N__22885\
        );

    \I__4355\ : Span4Mux_h
    port map (
            O => \N__22906\,
            I => \N__22885\
        );

    \I__4354\ : Span4Mux_s2_v
    port map (
            O => \N__22903\,
            I => \N__22885\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__22898\,
            I => \tok.n4_adj_726\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__22895\,
            I => \tok.n4_adj_726\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__22892\,
            I => \tok.n4_adj_726\
        );

    \I__4350\ : Odrv4
    port map (
            O => \N__22885\,
            I => \tok.n4_adj_726\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__22876\,
            I => \N__22871\
        );

    \I__4348\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22865\
        );

    \I__4347\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22860\
        );

    \I__4346\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22857\
        );

    \I__4345\ : InMux
    port map (
            O => \N__22870\,
            I => \N__22854\
        );

    \I__4344\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22851\
        );

    \I__4343\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22848\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__22865\,
            I => \N__22845\
        );

    \I__4341\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22842\
        );

    \I__4340\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22839\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__22860\,
            I => \N__22832\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__22857\,
            I => \N__22832\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__22854\,
            I => \N__22832\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__22851\,
            I => \N__22827\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__22848\,
            I => \N__22827\
        );

    \I__4334\ : Span4Mux_h
    port map (
            O => \N__22845\,
            I => \N__22818\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__22842\,
            I => \N__22818\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__22839\,
            I => \N__22818\
        );

    \I__4331\ : Span4Mux_h
    port map (
            O => \N__22832\,
            I => \N__22818\
        );

    \I__4330\ : Span4Mux_h
    port map (
            O => \N__22827\,
            I => \N__22815\
        );

    \I__4329\ : Span4Mux_v
    port map (
            O => \N__22818\,
            I => \N__22812\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__22815\,
            I => \tok.tc__7__N_133\
        );

    \I__4327\ : Odrv4
    port map (
            O => \N__22812\,
            I => \tok.tc__7__N_133\
        );

    \I__4326\ : InMux
    port map (
            O => \N__22807\,
            I => \N__22803\
        );

    \I__4325\ : InMux
    port map (
            O => \N__22806\,
            I => \N__22798\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__22803\,
            I => \N__22795\
        );

    \I__4323\ : InMux
    port map (
            O => \N__22802\,
            I => \N__22792\
        );

    \I__4322\ : InMux
    port map (
            O => \N__22801\,
            I => \N__22787\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__22798\,
            I => \N__22780\
        );

    \I__4320\ : Span4Mux_s3_v
    port map (
            O => \N__22795\,
            I => \N__22780\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__22792\,
            I => \N__22780\
        );

    \I__4318\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22776\
        );

    \I__4317\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22772\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__22787\,
            I => \N__22769\
        );

    \I__4315\ : Span4Mux_h
    port map (
            O => \N__22780\,
            I => \N__22766\
        );

    \I__4314\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22763\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__22776\,
            I => \N__22760\
        );

    \I__4312\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22757\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__22772\,
            I => \tok.n2573\
        );

    \I__4310\ : Odrv12
    port map (
            O => \N__22769\,
            I => \tok.n2573\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__22766\,
            I => \tok.n2573\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__22763\,
            I => \tok.n2573\
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__22760\,
            I => \tok.n2573\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__22757\,
            I => \tok.n2573\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__22744\,
            I => \tok.n6291_cascade_\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__22741\,
            I => \tok.n80_adj_735_cascade_\
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__22738\,
            I => \tok.n83_adj_725_cascade_\
        );

    \I__4302\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22732\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__22732\,
            I => \tok.n6287\
        );

    \I__4300\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22726\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__22726\,
            I => \tok.n89_adj_736\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__22723\,
            I => \N__22720\
        );

    \I__4297\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22716\
        );

    \I__4296\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22713\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22710\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__22713\,
            I => \N__22707\
        );

    \I__4293\ : Span4Mux_h
    port map (
            O => \N__22710\,
            I => \N__22702\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__22707\,
            I => \N__22702\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__22702\,
            I => n92
        );

    \I__4290\ : InMux
    port map (
            O => \N__22699\,
            I => \N__22693\
        );

    \I__4289\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22693\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__22693\,
            I => \tok.tail_10\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__22690\,
            I => \N__22687\
        );

    \I__4286\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22681\
        );

    \I__4285\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22681\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__22681\,
            I => \tok.C_stk.tail_18\
        );

    \I__4283\ : InMux
    port map (
            O => \N__22678\,
            I => \N__22672\
        );

    \I__4282\ : InMux
    port map (
            O => \N__22677\,
            I => \N__22672\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__22672\,
            I => \tok.tail_26\
        );

    \I__4280\ : InMux
    port map (
            O => \N__22669\,
            I => \N__22663\
        );

    \I__4279\ : InMux
    port map (
            O => \N__22668\,
            I => \N__22663\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__22663\,
            I => \tok.C_stk.tail_34\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__22660\,
            I => \N__22656\
        );

    \I__4276\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22650\
        );

    \I__4275\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22650\
        );

    \I__4274\ : InMux
    port map (
            O => \N__22655\,
            I => \N__22647\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__22650\,
            I => \N__22643\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__22647\,
            I => \N__22640\
        );

    \I__4271\ : InMux
    port map (
            O => \N__22646\,
            I => \N__22637\
        );

    \I__4270\ : Span4Mux_v
    port map (
            O => \N__22643\,
            I => \N__22634\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__22640\,
            I => \N__22627\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__22637\,
            I => \N__22627\
        );

    \I__4267\ : Span4Mux_s1_v
    port map (
            O => \N__22634\,
            I => \N__22627\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__22627\,
            I => \tok.tc_plus_1_3\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__22624\,
            I => \tok.C_stk.n6242_cascade_\
        );

    \I__4264\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22617\
        );

    \I__4263\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22614\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__22617\,
            I => \N__22611\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__22614\,
            I => \N__22607\
        );

    \I__4260\ : Span4Mux_h
    port map (
            O => \N__22611\,
            I => \N__22603\
        );

    \I__4259\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22600\
        );

    \I__4258\ : Span4Mux_v
    port map (
            O => \N__22607\,
            I => \N__22597\
        );

    \I__4257\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22594\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__22603\,
            I => tc_3
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__22600\,
            I => tc_3
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__22597\,
            I => tc_3
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__22594\,
            I => tc_3
        );

    \I__4252\ : InMux
    port map (
            O => \N__22585\,
            I => \N__22579\
        );

    \I__4251\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22572\
        );

    \I__4250\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22572\
        );

    \I__4249\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22572\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__22579\,
            I => \tok.c_stk_r_3\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__22572\,
            I => \tok.c_stk_r_3\
        );

    \I__4246\ : InMux
    port map (
            O => \N__22567\,
            I => \N__22561\
        );

    \I__4245\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22561\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__22561\,
            I => \tok.C_stk.tail_3\
        );

    \I__4243\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22552\
        );

    \I__4242\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22552\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__22552\,
            I => \tok.C_stk.tail_11\
        );

    \I__4240\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22543\
        );

    \I__4239\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22543\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__22543\,
            I => \tok.C_stk.tail_5\
        );

    \I__4237\ : InMux
    port map (
            O => \N__22540\,
            I => \N__22534\
        );

    \I__4236\ : InMux
    port map (
            O => \N__22539\,
            I => \N__22534\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__22534\,
            I => \tok.tail_13\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__22531\,
            I => \N__22528\
        );

    \I__4233\ : InMux
    port map (
            O => \N__22528\,
            I => \N__22522\
        );

    \I__4232\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22522\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__22522\,
            I => \tok.C_stk.tail_21\
        );

    \I__4230\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22513\
        );

    \I__4229\ : InMux
    port map (
            O => \N__22518\,
            I => \N__22513\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__22513\,
            I => \tok.tail_29\
        );

    \I__4227\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22504\
        );

    \I__4226\ : InMux
    port map (
            O => \N__22509\,
            I => \N__22504\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__22504\,
            I => \tok.C_stk.tail_37\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__22501\,
            I => \N__22498\
        );

    \I__4223\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22491\
        );

    \I__4222\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22491\
        );

    \I__4221\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22488\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__22491\,
            I => \N__22484\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__22488\,
            I => \N__22481\
        );

    \I__4218\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22478\
        );

    \I__4217\ : Span4Mux_h
    port map (
            O => \N__22484\,
            I => \N__22475\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__22481\,
            I => \tok.tc_plus_1_2\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__22478\,
            I => \tok.tc_plus_1_2\
        );

    \I__4214\ : Odrv4
    port map (
            O => \N__22475\,
            I => \tok.tc_plus_1_2\
        );

    \I__4213\ : CascadeMux
    port map (
            O => \N__22468\,
            I => \tok.C_stk.n6245_cascade_\
        );

    \I__4212\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22461\
        );

    \I__4211\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22457\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__22461\,
            I => \N__22453\
        );

    \I__4209\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22450\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__22457\,
            I => \N__22447\
        );

    \I__4207\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22444\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__22453\,
            I => tc_2
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__22450\,
            I => tc_2
        );

    \I__4204\ : Odrv12
    port map (
            O => \N__22447\,
            I => tc_2
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__22444\,
            I => tc_2
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__22435\,
            I => \N__22429\
        );

    \I__4201\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22426\
        );

    \I__4200\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22421\
        );

    \I__4199\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22421\
        );

    \I__4198\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22418\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__22426\,
            I => \tok.c_stk_r_2\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__22421\,
            I => \tok.c_stk_r_2\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__22418\,
            I => \tok.c_stk_r_2\
        );

    \I__4194\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22405\
        );

    \I__4193\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22405\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__22405\,
            I => \tok.C_stk.tail_2\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__22402\,
            I => \tok.n6404_cascade_\
        );

    \I__4190\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22396\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__22396\,
            I => \tok.n179_adj_888\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__22393\,
            I => \tok.n6550_cascade_\
        );

    \I__4187\ : InMux
    port map (
            O => \N__22390\,
            I => \N__22387\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__22387\,
            I => \N__22384\
        );

    \I__4185\ : Odrv4
    port map (
            O => \N__22384\,
            I => \tok.n6549\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__22381\,
            I => \N__22378\
        );

    \I__4183\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22375\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__22375\,
            I => \tok.n6419\
        );

    \I__4181\ : InMux
    port map (
            O => \N__22372\,
            I => \N__22369\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__22369\,
            I => \N__22366\
        );

    \I__4179\ : Span4Mux_s1_v
    port map (
            O => \N__22366\,
            I => \N__22363\
        );

    \I__4178\ : Odrv4
    port map (
            O => \N__22363\,
            I => \tok.n215_adj_697\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__22360\,
            I => \tok.n6337_cascade_\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__22357\,
            I => \N__22354\
        );

    \I__4175\ : InMux
    port map (
            O => \N__22354\,
            I => \N__22351\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__22351\,
            I => \tok.n6538\
        );

    \I__4173\ : InMux
    port map (
            O => \N__22348\,
            I => \N__22344\
        );

    \I__4172\ : InMux
    port map (
            O => \N__22347\,
            I => \N__22341\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__22344\,
            I => \N__22338\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__22341\,
            I => \N__22335\
        );

    \I__4169\ : Span4Mux_h
    port map (
            O => \N__22338\,
            I => \N__22328\
        );

    \I__4168\ : Span4Mux_v
    port map (
            O => \N__22335\,
            I => \N__22328\
        );

    \I__4167\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22323\
        );

    \I__4166\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22323\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__22328\,
            I => \tok.tc_plus_1_5\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__22323\,
            I => \tok.tc_plus_1_5\
        );

    \I__4163\ : CascadeMux
    port map (
            O => \N__22318\,
            I => \tok.C_stk.n6236_cascade_\
        );

    \I__4162\ : InMux
    port map (
            O => \N__22315\,
            I => \N__22312\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__22312\,
            I => \N__22309\
        );

    \I__4160\ : Span4Mux_s2_v
    port map (
            O => \N__22309\,
            I => \N__22303\
        );

    \I__4159\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22298\
        );

    \I__4158\ : InMux
    port map (
            O => \N__22307\,
            I => \N__22298\
        );

    \I__4157\ : InMux
    port map (
            O => \N__22306\,
            I => \N__22295\
        );

    \I__4156\ : Odrv4
    port map (
            O => \N__22303\,
            I => tc_5
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__22298\,
            I => tc_5
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__22295\,
            I => tc_5
        );

    \I__4153\ : InMux
    port map (
            O => \N__22288\,
            I => \N__22279\
        );

    \I__4152\ : InMux
    port map (
            O => \N__22287\,
            I => \N__22279\
        );

    \I__4151\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22279\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__22279\,
            I => \N__22275\
        );

    \I__4149\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22272\
        );

    \I__4148\ : Span4Mux_v
    port map (
            O => \N__22275\,
            I => \N__22269\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__22272\,
            I => \tok.c_stk_r_5\
        );

    \I__4146\ : Odrv4
    port map (
            O => \N__22269\,
            I => \tok.c_stk_r_5\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__22264\,
            I => \N__22261\
        );

    \I__4144\ : InMux
    port map (
            O => \N__22261\,
            I => \N__22258\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__22258\,
            I => \tok.n6320\
        );

    \I__4142\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22252\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__22252\,
            I => \N__22246\
        );

    \I__4140\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22237\
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__22250\,
            I => \N__22234\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__22249\,
            I => \N__22229\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__22246\,
            I => \N__22225\
        );

    \I__4136\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22218\
        );

    \I__4135\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22218\
        );

    \I__4134\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22218\
        );

    \I__4133\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22215\
        );

    \I__4132\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22212\
        );

    \I__4131\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22209\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22206\
        );

    \I__4129\ : InMux
    port map (
            O => \N__22234\,
            I => \N__22203\
        );

    \I__4128\ : InMux
    port map (
            O => \N__22233\,
            I => \N__22200\
        );

    \I__4127\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22195\
        );

    \I__4126\ : InMux
    port map (
            O => \N__22229\,
            I => \N__22195\
        );

    \I__4125\ : InMux
    port map (
            O => \N__22228\,
            I => \N__22192\
        );

    \I__4124\ : Span4Mux_v
    port map (
            O => \N__22225\,
            I => \N__22185\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__22218\,
            I => \N__22182\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__22215\,
            I => \N__22179\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__22212\,
            I => \N__22176\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__22209\,
            I => \N__22173\
        );

    \I__4119\ : Span4Mux_v
    port map (
            O => \N__22206\,
            I => \N__22168\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__22203\,
            I => \N__22168\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__22200\,
            I => \N__22162\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__22195\,
            I => \N__22162\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__22192\,
            I => \N__22159\
        );

    \I__4114\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22154\
        );

    \I__4113\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22154\
        );

    \I__4112\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22149\
        );

    \I__4111\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22149\
        );

    \I__4110\ : Span4Mux_s3_h
    port map (
            O => \N__22185\,
            I => \N__22144\
        );

    \I__4109\ : Span4Mux_s2_v
    port map (
            O => \N__22182\,
            I => \N__22144\
        );

    \I__4108\ : Span4Mux_h
    port map (
            O => \N__22179\,
            I => \N__22139\
        );

    \I__4107\ : Span4Mux_h
    port map (
            O => \N__22176\,
            I => \N__22139\
        );

    \I__4106\ : Span4Mux_h
    port map (
            O => \N__22173\,
            I => \N__22134\
        );

    \I__4105\ : Span4Mux_h
    port map (
            O => \N__22168\,
            I => \N__22134\
        );

    \I__4104\ : InMux
    port map (
            O => \N__22167\,
            I => \N__22131\
        );

    \I__4103\ : Span4Mux_v
    port map (
            O => \N__22162\,
            I => \N__22128\
        );

    \I__4102\ : Span4Mux_s2_v
    port map (
            O => \N__22159\,
            I => \N__22123\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__22154\,
            I => \N__22123\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__22149\,
            I => \tok.n49\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__22144\,
            I => \tok.n49\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__22139\,
            I => \tok.n49\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__22134\,
            I => \tok.n49\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__22131\,
            I => \tok.n49\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__22128\,
            I => \tok.n49\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__22123\,
            I => \tok.n49\
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__22108\,
            I => \tok.n6380_cascade_\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__22105\,
            I => \tok.n215_adj_656_cascade_\
        );

    \I__4091\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22099\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__22099\,
            I => \N__22096\
        );

    \I__4089\ : Odrv4
    port map (
            O => \N__22096\,
            I => \tok.n2665\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__22093\,
            I => \N__22090\
        );

    \I__4087\ : InMux
    port map (
            O => \N__22090\,
            I => \N__22087\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__22087\,
            I => \tok.n4_adj_719\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__22084\,
            I => \tok.n4_adj_719_cascade_\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__22081\,
            I => \N__22078\
        );

    \I__4083\ : InMux
    port map (
            O => \N__22078\,
            I => \N__22075\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__22075\,
            I => \N__22072\
        );

    \I__4081\ : Span12Mux_s7_v
    port map (
            O => \N__22072\,
            I => \N__22069\
        );

    \I__4080\ : Odrv12
    port map (
            O => \N__22069\,
            I => \tok.n10_adj_809\
        );

    \I__4079\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22063\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__22063\,
            I => \N__22060\
        );

    \I__4077\ : Odrv12
    port map (
            O => \N__22060\,
            I => \tok.n6411\
        );

    \I__4076\ : InMux
    port map (
            O => \N__22057\,
            I => \N__22054\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__22054\,
            I => \N__22051\
        );

    \I__4074\ : Span4Mux_h
    port map (
            O => \N__22051\,
            I => \N__22048\
        );

    \I__4073\ : Span4Mux_v
    port map (
            O => \N__22048\,
            I => \N__22045\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__22045\,
            I => \tok.n6532\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__22042\,
            I => \tok.n207_adj_771_cascade_\
        );

    \I__4070\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22036\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__22036\,
            I => \N__22033\
        );

    \I__4068\ : Odrv12
    port map (
            O => \N__22033\,
            I => \tok.n6583\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__22030\,
            I => \N__22024\
        );

    \I__4066\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22021\
        );

    \I__4065\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22018\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__22027\,
            I => \N__22015\
        );

    \I__4063\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22011\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__22021\,
            I => \N__22006\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__22018\,
            I => \N__22006\
        );

    \I__4060\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22003\
        );

    \I__4059\ : InMux
    port map (
            O => \N__22014\,
            I => \N__22000\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__22011\,
            I => \N__21997\
        );

    \I__4057\ : Span4Mux_v
    port map (
            O => \N__22006\,
            I => \N__21992\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__22003\,
            I => \N__21992\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__22000\,
            I => \N__21988\
        );

    \I__4054\ : Span4Mux_h
    port map (
            O => \N__21997\,
            I => \N__21983\
        );

    \I__4053\ : Span4Mux_h
    port map (
            O => \N__21992\,
            I => \N__21980\
        );

    \I__4052\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21977\
        );

    \I__4051\ : Span4Mux_v
    port map (
            O => \N__21988\,
            I => \N__21974\
        );

    \I__4050\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21971\
        );

    \I__4049\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21968\
        );

    \I__4048\ : Span4Mux_h
    port map (
            O => \N__21983\,
            I => \N__21965\
        );

    \I__4047\ : Span4Mux_h
    port map (
            O => \N__21980\,
            I => \N__21962\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__21977\,
            I => \N__21955\
        );

    \I__4045\ : Sp12to4
    port map (
            O => \N__21974\,
            I => \N__21955\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__21971\,
            I => \N__21955\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__21968\,
            I => \tok.S_5\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__21965\,
            I => \tok.S_5\
        );

    \I__4041\ : Odrv4
    port map (
            O => \N__21962\,
            I => \tok.S_5\
        );

    \I__4040\ : Odrv12
    port map (
            O => \N__21955\,
            I => \tok.S_5\
        );

    \I__4039\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21943\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__21943\,
            I => \tok.n213\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__21940\,
            I => \tok.n207_adj_776_cascade_\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__21937\,
            I => \tok.n6529_cascade_\
        );

    \I__4035\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21931\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__21931\,
            I => \N__21928\
        );

    \I__4033\ : Span4Mux_v
    port map (
            O => \N__21928\,
            I => \N__21925\
        );

    \I__4032\ : Odrv4
    port map (
            O => \N__21925\,
            I => \tok.n210_adj_784\
        );

    \I__4031\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21919\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__21919\,
            I => \tok.n174_adj_785\
        );

    \I__4029\ : InMux
    port map (
            O => \N__21916\,
            I => \N__21913\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__21913\,
            I => \N__21910\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__21910\,
            I => \N__21907\
        );

    \I__4026\ : Span4Mux_v
    port map (
            O => \N__21907\,
            I => \N__21904\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__21904\,
            I => \tok.n229_adj_861\
        );

    \I__4024\ : CascadeMux
    port map (
            O => \N__21901\,
            I => \N__21898\
        );

    \I__4023\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21895\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__21895\,
            I => \tok.n6365\
        );

    \I__4021\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21889\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__21889\,
            I => \N__21886\
        );

    \I__4019\ : Sp12to4
    port map (
            O => \N__21886\,
            I => \N__21883\
        );

    \I__4018\ : Odrv12
    port map (
            O => \N__21883\,
            I => \tok.n215_adj_672\
        );

    \I__4017\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21877\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__21877\,
            I => \N__21874\
        );

    \I__4015\ : Span4Mux_h
    port map (
            O => \N__21874\,
            I => \N__21871\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__21871\,
            I => \tok.n252\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__21868\,
            I => \tok.n4_adj_769_cascade_\
        );

    \I__4012\ : InMux
    port map (
            O => \N__21865\,
            I => \N__21862\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__21862\,
            I => \tok.n205_adj_770\
        );

    \I__4010\ : InMux
    port map (
            O => \N__21859\,
            I => \N__21855\
        );

    \I__4009\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21852\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__21855\,
            I => \N__21849\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__21852\,
            I => \N__21846\
        );

    \I__4006\ : Span4Mux_v
    port map (
            O => \N__21849\,
            I => \N__21841\
        );

    \I__4005\ : Span4Mux_v
    port map (
            O => \N__21846\,
            I => \N__21841\
        );

    \I__4004\ : Sp12to4
    port map (
            O => \N__21841\,
            I => \N__21838\
        );

    \I__4003\ : Odrv12
    port map (
            O => \N__21838\,
            I => \tok.n235\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__21835\,
            I => \tok.n190_cascade_\
        );

    \I__4001\ : InMux
    port map (
            O => \N__21832\,
            I => \N__21829\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__21829\,
            I => \tok.n190\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__21826\,
            I => \tok.n255_cascade_\
        );

    \I__3998\ : InMux
    port map (
            O => \N__21823\,
            I => \N__21820\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__21820\,
            I => \tok.n258\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__21817\,
            I => \tok.n6508_cascade_\
        );

    \I__3995\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21811\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__21811\,
            I => \tok.n210_adj_816\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__21808\,
            I => \tok.n872_cascade_\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__21805\,
            I => \tok.n174_adj_817_cascade_\
        );

    \I__3991\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21799\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__21799\,
            I => \tok.n4_adj_818\
        );

    \I__3989\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21793\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__21793\,
            I => \tok.n205_adj_820\
        );

    \I__3987\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__21787\,
            I => \N__21784\
        );

    \I__3985\ : Odrv12
    port map (
            O => \N__21784\,
            I => \tok.n200_adj_840\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__21781\,
            I => \tok.n6_adj_843_cascade_\
        );

    \I__3983\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21774\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__21777\,
            I => \N__21769\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__21774\,
            I => \N__21765\
        );

    \I__3980\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21762\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__21772\,
            I => \N__21758\
        );

    \I__3978\ : InMux
    port map (
            O => \N__21769\,
            I => \N__21755\
        );

    \I__3977\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21752\
        );

    \I__3976\ : Span4Mux_v
    port map (
            O => \N__21765\,
            I => \N__21747\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__21762\,
            I => \N__21747\
        );

    \I__3974\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21744\
        );

    \I__3973\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21741\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__21755\,
            I => \N__21738\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__21752\,
            I => \N__21734\
        );

    \I__3970\ : Span4Mux_h
    port map (
            O => \N__21747\,
            I => \N__21731\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__21744\,
            I => \N__21726\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__21741\,
            I => \N__21726\
        );

    \I__3967\ : Span4Mux_v
    port map (
            O => \N__21738\,
            I => \N__21723\
        );

    \I__3966\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21720\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__21734\,
            I => \N__21717\
        );

    \I__3964\ : Span4Mux_h
    port map (
            O => \N__21731\,
            I => \N__21714\
        );

    \I__3963\ : Span4Mux_v
    port map (
            O => \N__21726\,
            I => \N__21711\
        );

    \I__3962\ : Span4Mux_h
    port map (
            O => \N__21723\,
            I => \N__21708\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__21720\,
            I => \tok.S_9\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__21717\,
            I => \tok.S_9\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__21714\,
            I => \tok.S_9\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__21711\,
            I => \tok.S_9\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__21708\,
            I => \tok.S_9\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__21697\,
            I => \tok.n6440_cascade_\
        );

    \I__3955\ : CascadeMux
    port map (
            O => \N__21694\,
            I => \tok.n6612_cascade_\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__21691\,
            I => \tok.n179_cascade_\
        );

    \I__3953\ : InMux
    port map (
            O => \N__21688\,
            I => \N__21685\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__21685\,
            I => \tok.n6546\
        );

    \I__3951\ : CascadeMux
    port map (
            O => \N__21682\,
            I => \N__21678\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__21681\,
            I => \N__21675\
        );

    \I__3949\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21672\
        );

    \I__3948\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21669\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__21672\,
            I => \N__21666\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__21669\,
            I => \N__21663\
        );

    \I__3945\ : Span4Mux_v
    port map (
            O => \N__21666\,
            I => \N__21660\
        );

    \I__3944\ : Span4Mux_v
    port map (
            O => \N__21663\,
            I => \N__21657\
        );

    \I__3943\ : Span4Mux_h
    port map (
            O => \N__21660\,
            I => \N__21654\
        );

    \I__3942\ : Span4Mux_v
    port map (
            O => \N__21657\,
            I => \N__21651\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__21654\,
            I => \tok.table_rd_7\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__21651\,
            I => \tok.table_rd_7\
        );

    \I__3939\ : CascadeMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__3938\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21639\
        );

    \I__3937\ : InMux
    port map (
            O => \N__21642\,
            I => \N__21636\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__21639\,
            I => \N__21633\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__21636\,
            I => \N__21630\
        );

    \I__3934\ : Span4Mux_v
    port map (
            O => \N__21633\,
            I => \N__21627\
        );

    \I__3933\ : Span12Mux_s9_v
    port map (
            O => \N__21630\,
            I => \N__21624\
        );

    \I__3932\ : Span4Mux_h
    port map (
            O => \N__21627\,
            I => \N__21621\
        );

    \I__3931\ : Odrv12
    port map (
            O => \N__21624\,
            I => \tok.table_rd_4\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__21621\,
            I => \tok.table_rd_4\
        );

    \I__3929\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21613\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__21613\,
            I => \tok.n258_adj_814\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__21610\,
            I => \tok.n252_adj_815_cascade_\
        );

    \I__3926\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21603\
        );

    \I__3925\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21600\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__21603\,
            I => \N__21595\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__21600\,
            I => \N__21595\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__21595\,
            I => \N__21592\
        );

    \I__3921\ : Span4Mux_h
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__21589\,
            I => \tok.n232\
        );

    \I__3919\ : InMux
    port map (
            O => \N__21586\,
            I => \N__21583\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__21583\,
            I => \tok.n255_adj_808\
        );

    \I__3917\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21577\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__21577\,
            I => \tok.n311_adj_721\
        );

    \I__3915\ : CascadeMux
    port map (
            O => \N__21574\,
            I => \tok.n167_cascade_\
        );

    \I__3914\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21568\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__21568\,
            I => \N__21565\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__21565\,
            I => \tok.n6567\
        );

    \I__3911\ : InMux
    port map (
            O => \N__21562\,
            I => \N__21558\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__21561\,
            I => \N__21555\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__21558\,
            I => \N__21552\
        );

    \I__3908\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21549\
        );

    \I__3907\ : Span4Mux_v
    port map (
            O => \N__21552\,
            I => \N__21544\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__21549\,
            I => \N__21544\
        );

    \I__3905\ : Span4Mux_v
    port map (
            O => \N__21544\,
            I => \N__21541\
        );

    \I__3904\ : Span4Mux_h
    port map (
            O => \N__21541\,
            I => \N__21538\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__21538\,
            I => \tok.table_rd_2\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__21535\,
            I => \tok.n209_cascade_\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__21532\,
            I => \tok.n6625_cascade_\
        );

    \I__3900\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21526\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__21526\,
            I => \tok.n6624\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__21523\,
            I => \tok.n168_adj_700_cascade_\
        );

    \I__3897\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21517\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__21517\,
            I => \tok.n6569\
        );

    \I__3895\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21511\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__21511\,
            I => \N__21508\
        );

    \I__3893\ : Span4Mux_h
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__21505\,
            I => \tok.n2548\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__21502\,
            I => \N__21499\
        );

    \I__3890\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21496\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__3888\ : Span4Mux_v
    port map (
            O => \N__21493\,
            I => \N__21490\
        );

    \I__3887\ : Odrv4
    port map (
            O => \N__21490\,
            I => \tok.n6396\
        );

    \I__3886\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21481\
        );

    \I__3885\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21481\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__21481\,
            I => \N__21477\
        );

    \I__3883\ : InMux
    port map (
            O => \N__21480\,
            I => \N__21474\
        );

    \I__3882\ : Span4Mux_v
    port map (
            O => \N__21477\,
            I => \N__21471\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__21474\,
            I => \N__21468\
        );

    \I__3880\ : Span4Mux_v
    port map (
            O => \N__21471\,
            I => \N__21465\
        );

    \I__3879\ : Span4Mux_h
    port map (
            O => \N__21468\,
            I => \N__21462\
        );

    \I__3878\ : Span4Mux_h
    port map (
            O => \N__21465\,
            I => \N__21459\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__21462\,
            I => \N__21456\
        );

    \I__3876\ : Odrv4
    port map (
            O => \N__21459\,
            I => \tok.n236\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__21456\,
            I => \tok.n236\
        );

    \I__3874\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21448\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__21448\,
            I => \tok.n4925\
        );

    \I__3872\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21442\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__21442\,
            I => \N__21439\
        );

    \I__3870\ : Span4Mux_h
    port map (
            O => \N__21439\,
            I => \N__21436\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__21436\,
            I => \tok.n288\
        );

    \I__3868\ : InMux
    port map (
            O => \N__21433\,
            I => \N__21430\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__21430\,
            I => \N__21427\
        );

    \I__3866\ : Span4Mux_v
    port map (
            O => \N__21427\,
            I => \N__21424\
        );

    \I__3865\ : Span4Mux_h
    port map (
            O => \N__21424\,
            I => \N__21421\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__21421\,
            I => \tok.n2613\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__21418\,
            I => \tok.n6578_cascade_\
        );

    \I__3862\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21412\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__21412\,
            I => \N__21409\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__21409\,
            I => \tok.n6581\
        );

    \I__3859\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21403\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__21403\,
            I => \tok.n4_adj_739\
        );

    \I__3857\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21397\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__21397\,
            I => \tok.n2611\
        );

    \I__3855\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21391\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__21391\,
            I => \N__21388\
        );

    \I__3853\ : Span4Mux_h
    port map (
            O => \N__21388\,
            I => \N__21385\
        );

    \I__3852\ : Odrv4
    port map (
            O => \N__21385\,
            I => \tok.n6580\
        );

    \I__3851\ : InMux
    port map (
            O => \N__21382\,
            I => \N__21376\
        );

    \I__3850\ : InMux
    port map (
            O => \N__21381\,
            I => \N__21376\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__21376\,
            I => \tok.n4_adj_684\
        );

    \I__3848\ : CascadeMux
    port map (
            O => \N__21373\,
            I => \tok.n6620_cascade_\
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__21370\,
            I => \tok.n14_adj_683_cascade_\
        );

    \I__3846\ : InMux
    port map (
            O => \N__21367\,
            I => \N__21364\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__21364\,
            I => \N__21360\
        );

    \I__3844\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21357\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__21360\,
            I => \tok.n9_adj_651\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__21357\,
            I => \tok.n9_adj_651\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__21352\,
            I => \tok.n15_adj_807_cascade_\
        );

    \I__3840\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21343\
        );

    \I__3839\ : InMux
    port map (
            O => \N__21348\,
            I => \N__21343\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__21343\,
            I => \N__21340\
        );

    \I__3837\ : Odrv12
    port map (
            O => \N__21340\,
            I => \tok.n903\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__21337\,
            I => \N__21334\
        );

    \I__3835\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21331\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__21331\,
            I => \N__21328\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__21328\,
            I => \tok.n14_adj_683\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__21325\,
            I => \N__21322\
        );

    \I__3831\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21319\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__21319\,
            I => \tok.n6621\
        );

    \I__3829\ : InMux
    port map (
            O => \N__21316\,
            I => \N__21313\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__21313\,
            I => \tok.n241_adj_747\
        );

    \I__3827\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21307\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21304\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__21304\,
            I => \tok.n6593\
        );

    \I__3824\ : InMux
    port map (
            O => \N__21301\,
            I => \N__21298\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__21298\,
            I => \tok.n6664\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__21295\,
            I => \tok.n1600_cascade_\
        );

    \I__3821\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21289\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__21289\,
            I => \tok.n13_adj_742\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__21286\,
            I => \tok.n6301_cascade_\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__21283\,
            I => \tok.n80_adj_751_cascade_\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__21280\,
            I => \tok.n83_adj_746_cascade_\
        );

    \I__3816\ : InMux
    port map (
            O => \N__21277\,
            I => \N__21274\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__21274\,
            I => \tok.n6297\
        );

    \I__3814\ : InMux
    port map (
            O => \N__21271\,
            I => \N__21268\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__21268\,
            I => \tok.n89_adj_754\
        );

    \I__3812\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21261\
        );

    \I__3811\ : InMux
    port map (
            O => \N__21264\,
            I => \N__21258\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__21261\,
            I => \N__21255\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__21258\,
            I => \N__21252\
        );

    \I__3808\ : Span4Mux_h
    port map (
            O => \N__21255\,
            I => \N__21249\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__21252\,
            I => n92_adj_898
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__21249\,
            I => n92_adj_898
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__21244\,
            I => \N__21240\
        );

    \I__3804\ : InMux
    port map (
            O => \N__21243\,
            I => \N__21235\
        );

    \I__3803\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21235\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__21235\,
            I => \N__21232\
        );

    \I__3801\ : Span4Mux_h
    port map (
            O => \N__21232\,
            I => \N__21229\
        );

    \I__3800\ : Span4Mux_h
    port map (
            O => \N__21229\,
            I => \N__21226\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__21226\,
            I => \N__21223\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__21223\,
            I => \tok.table_rd_3\
        );

    \I__3797\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21214\
        );

    \I__3796\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21214\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__21214\,
            I => \tok.tail_28\
        );

    \I__3794\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21205\
        );

    \I__3793\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21205\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__21205\,
            I => \tok.C_stk.tail_36\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__21202\,
            I => \tok.n83_adj_723_cascade_\
        );

    \I__3790\ : InMux
    port map (
            O => \N__21199\,
            I => \N__21195\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__21198\,
            I => \N__21192\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__21195\,
            I => \N__21189\
        );

    \I__3787\ : InMux
    port map (
            O => \N__21192\,
            I => \N__21186\
        );

    \I__3786\ : Span4Mux_s1_v
    port map (
            O => \N__21189\,
            I => \N__21181\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21181\
        );

    \I__3784\ : Odrv4
    port map (
            O => \N__21181\,
            I => n10_adj_908
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__21178\,
            I => \tok.n4_adj_726_cascade_\
        );

    \I__3782\ : CascadeMux
    port map (
            O => \N__21175\,
            I => \tok.ram.n6257_cascade_\
        );

    \I__3781\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21168\
        );

    \I__3780\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21164\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__21168\,
            I => \N__21161\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__21167\,
            I => \N__21157\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__21164\,
            I => \N__21154\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__21161\,
            I => \N__21151\
        );

    \I__3775\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21146\
        );

    \I__3774\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21146\
        );

    \I__3773\ : Span4Mux_s1_v
    port map (
            O => \N__21154\,
            I => \N__21143\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__21151\,
            I => \N__21138\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__21146\,
            I => \N__21138\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__21143\,
            I => tc_plus_1_0
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__21138\,
            I => tc_plus_1_0
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__21133\,
            I => \tok.C_stk.n6230_cascade_\
        );

    \I__3767\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21125\
        );

    \I__3766\ : InMux
    port map (
            O => \N__21129\,
            I => \N__21121\
        );

    \I__3765\ : InMux
    port map (
            O => \N__21128\,
            I => \N__21118\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__21125\,
            I => \N__21115\
        );

    \I__3763\ : InMux
    port map (
            O => \N__21124\,
            I => \N__21112\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__21121\,
            I => tc_0
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__21118\,
            I => tc_0
        );

    \I__3760\ : Odrv12
    port map (
            O => \N__21115\,
            I => tc_0
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__21112\,
            I => tc_0
        );

    \I__3758\ : CascadeMux
    port map (
            O => \N__21103\,
            I => \N__21098\
        );

    \I__3757\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21095\
        );

    \I__3756\ : InMux
    port map (
            O => \N__21101\,
            I => \N__21090\
        );

    \I__3755\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21090\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__21095\,
            I => \N__21084\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__21090\,
            I => \N__21084\
        );

    \I__3752\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21081\
        );

    \I__3751\ : Span4Mux_h
    port map (
            O => \N__21084\,
            I => \N__21078\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__21081\,
            I => c_stk_r_0
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__21078\,
            I => c_stk_r_0
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__21073\,
            I => \N__21070\
        );

    \I__3747\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21064\
        );

    \I__3746\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21064\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__21064\,
            I => \tok.C_stk.tail_0\
        );

    \I__3744\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21058\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21052\
        );

    \I__3742\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21049\
        );

    \I__3741\ : InMux
    port map (
            O => \N__21056\,
            I => \N__21044\
        );

    \I__3740\ : InMux
    port map (
            O => \N__21055\,
            I => \N__21044\
        );

    \I__3739\ : Odrv4
    port map (
            O => \N__21052\,
            I => \tok.tc_plus_1_4\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__21049\,
            I => \tok.tc_plus_1_4\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__21044\,
            I => \tok.tc_plus_1_4\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__21037\,
            I => \tok.C_stk.n6239_cascade_\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__21034\,
            I => \N__21030\
        );

    \I__3734\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21025\
        );

    \I__3733\ : InMux
    port map (
            O => \N__21030\,
            I => \N__21020\
        );

    \I__3732\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21020\
        );

    \I__3731\ : InMux
    port map (
            O => \N__21028\,
            I => \N__21017\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__21025\,
            I => tc_4
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__21020\,
            I => tc_4
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__21017\,
            I => tc_4
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__21010\,
            I => \N__21005\
        );

    \I__3726\ : InMux
    port map (
            O => \N__21009\,
            I => \N__21001\
        );

    \I__3725\ : InMux
    port map (
            O => \N__21008\,
            I => \N__20998\
        );

    \I__3724\ : InMux
    port map (
            O => \N__21005\,
            I => \N__20993\
        );

    \I__3723\ : InMux
    port map (
            O => \N__21004\,
            I => \N__20993\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__21001\,
            I => \tok.c_stk_r_4\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__20998\,
            I => \tok.c_stk_r_4\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__20993\,
            I => \tok.c_stk_r_4\
        );

    \I__3719\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20980\
        );

    \I__3718\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20980\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__20980\,
            I => \tok.C_stk.tail_4\
        );

    \I__3716\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20971\
        );

    \I__3715\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20971\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__20971\,
            I => \tok.tail_12\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__20968\,
            I => \N__20965\
        );

    \I__3712\ : InMux
    port map (
            O => \N__20965\,
            I => \N__20959\
        );

    \I__3711\ : InMux
    port map (
            O => \N__20964\,
            I => \N__20959\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__20959\,
            I => \tok.C_stk.tail_20\
        );

    \I__3709\ : InMux
    port map (
            O => \N__20956\,
            I => \N__20953\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__20953\,
            I => \tok.n6425\
        );

    \I__3707\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20947\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__20947\,
            I => \tok.n6346\
        );

    \I__3705\ : InMux
    port map (
            O => \N__20944\,
            I => \N__20941\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__20941\,
            I => \N__20938\
        );

    \I__3703\ : Odrv12
    port map (
            O => \N__20938\,
            I => \tok.n215_adj_876\
        );

    \I__3702\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20932\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__20932\,
            I => \tok.n179_adj_877\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__20929\,
            I => \tok.n6553_cascade_\
        );

    \I__3699\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20923\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__20923\,
            I => \N__20920\
        );

    \I__3697\ : Span4Mux_v
    port map (
            O => \N__20920\,
            I => \N__20917\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__20917\,
            I => \tok.n6552\
        );

    \I__3695\ : InMux
    port map (
            O => \N__20914\,
            I => \N__20911\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__20911\,
            I => \tok.n179_adj_698\
        );

    \I__3693\ : InMux
    port map (
            O => \N__20908\,
            I => \N__20905\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__20905\,
            I => \N__20902\
        );

    \I__3691\ : Odrv12
    port map (
            O => \N__20902\,
            I => \tok.n6537\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__20899\,
            I => \tok.n6541_cascade_\
        );

    \I__3689\ : InMux
    port map (
            O => \N__20896\,
            I => \N__20893\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__20893\,
            I => \N__20890\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__20890\,
            I => \N__20887\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__20887\,
            I => \tok.n6540\
        );

    \I__3685\ : InMux
    port map (
            O => \N__20884\,
            I => \N__20881\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__20881\,
            I => \N__20878\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__20878\,
            I => \tok.n6367\
        );

    \I__3682\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20872\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__20872\,
            I => \tok.n179_adj_673\
        );

    \I__3680\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20866\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__20866\,
            I => \tok.uart.sender_4\
        );

    \I__3678\ : InMux
    port map (
            O => \N__20863\,
            I => \N__20860\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__20860\,
            I => \N__20857\
        );

    \I__3676\ : Span4Mux_s2_v
    port map (
            O => \N__20857\,
            I => \N__20854\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__20854\,
            I => \tok.uart.sender_3\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__20851\,
            I => \N__20848\
        );

    \I__3673\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20845\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__20845\,
            I => \N__20842\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__20842\,
            I => \N__20839\
        );

    \I__3670\ : Odrv4
    port map (
            O => \N__20839\,
            I => \tok.n2602\
        );

    \I__3669\ : InMux
    port map (
            O => \N__20836\,
            I => \N__20833\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__20833\,
            I => \tok.n6450\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__20830\,
            I => \tok.n215_adj_830_cascade_\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__20827\,
            I => \tok.n6605_cascade_\
        );

    \I__3665\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__20821\,
            I => \N__20818\
        );

    \I__3663\ : Span4Mux_h
    port map (
            O => \N__20818\,
            I => \N__20815\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__20815\,
            I => \tok.n6604\
        );

    \I__3661\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20809\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__20809\,
            I => \N__20806\
        );

    \I__3659\ : Span4Mux_h
    port map (
            O => \N__20806\,
            I => \N__20803\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__20803\,
            I => \tok.n6456\
        );

    \I__3657\ : InMux
    port map (
            O => \N__20800\,
            I => \N__20797\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__20797\,
            I => \tok.n179_adj_831\
        );

    \I__3655\ : InMux
    port map (
            O => \N__20794\,
            I => \N__20789\
        );

    \I__3654\ : InMux
    port map (
            O => \N__20793\,
            I => \N__20786\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__20792\,
            I => \N__20782\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__20789\,
            I => \N__20778\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__20786\,
            I => \N__20775\
        );

    \I__3650\ : InMux
    port map (
            O => \N__20785\,
            I => \N__20770\
        );

    \I__3649\ : InMux
    port map (
            O => \N__20782\,
            I => \N__20770\
        );

    \I__3648\ : CascadeMux
    port map (
            O => \N__20781\,
            I => \N__20762\
        );

    \I__3647\ : Span4Mux_h
    port map (
            O => \N__20778\,
            I => \N__20751\
        );

    \I__3646\ : Span4Mux_h
    port map (
            O => \N__20775\,
            I => \N__20751\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__20770\,
            I => \N__20751\
        );

    \I__3644\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20748\
        );

    \I__3643\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20741\
        );

    \I__3642\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20741\
        );

    \I__3641\ : InMux
    port map (
            O => \N__20766\,
            I => \N__20741\
        );

    \I__3640\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20737\
        );

    \I__3639\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20734\
        );

    \I__3638\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20731\
        );

    \I__3637\ : InMux
    port map (
            O => \N__20760\,
            I => \N__20724\
        );

    \I__3636\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20724\
        );

    \I__3635\ : InMux
    port map (
            O => \N__20758\,
            I => \N__20724\
        );

    \I__3634\ : Span4Mux_h
    port map (
            O => \N__20751\,
            I => \N__20721\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__20748\,
            I => \N__20716\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__20741\,
            I => \N__20716\
        );

    \I__3631\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20713\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__20737\,
            I => \tok.n214\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__20734\,
            I => \tok.n214\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__20731\,
            I => \tok.n214\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__20724\,
            I => \tok.n214\
        );

    \I__3626\ : Odrv4
    port map (
            O => \N__20721\,
            I => \tok.n214\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__20716\,
            I => \tok.n214\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__20713\,
            I => \tok.n214\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__20698\,
            I => \tok.n6462_cascade_\
        );

    \I__3622\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20692\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__20692\,
            I => \N__20686\
        );

    \I__3620\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20683\
        );

    \I__3619\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20680\
        );

    \I__3618\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20674\
        );

    \I__3617\ : Span4Mux_v
    port map (
            O => \N__20686\,
            I => \N__20671\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__20683\,
            I => \N__20665\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__20680\,
            I => \N__20665\
        );

    \I__3614\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20660\
        );

    \I__3613\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20660\
        );

    \I__3612\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20657\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__20674\,
            I => \N__20653\
        );

    \I__3610\ : Span4Mux_v
    port map (
            O => \N__20671\,
            I => \N__20650\
        );

    \I__3609\ : InMux
    port map (
            O => \N__20670\,
            I => \N__20647\
        );

    \I__3608\ : Span12Mux_s11_h
    port map (
            O => \N__20665\,
            I => \N__20644\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__20660\,
            I => \N__20639\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__20657\,
            I => \N__20639\
        );

    \I__3605\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20636\
        );

    \I__3604\ : Span4Mux_s2_h
    port map (
            O => \N__20653\,
            I => \N__20633\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__20650\,
            I => \tok.n786\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__20647\,
            I => \tok.n786\
        );

    \I__3601\ : Odrv12
    port map (
            O => \N__20644\,
            I => \tok.n786\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__20639\,
            I => \tok.n786\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__20636\,
            I => \tok.n786\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__20633\,
            I => \tok.n786\
        );

    \I__3597\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20617\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__20617\,
            I => \tok.n206_adj_823\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__20614\,
            I => \N__20611\
        );

    \I__3594\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20607\
        );

    \I__3593\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20604\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__20607\,
            I => \N__20601\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__20604\,
            I => \N__20598\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__20601\,
            I => \N__20595\
        );

    \I__3589\ : Span4Mux_h
    port map (
            O => \N__20598\,
            I => \N__20590\
        );

    \I__3588\ : Span4Mux_v
    port map (
            O => \N__20595\,
            I => \N__20590\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__20590\,
            I => \tok.n314\
        );

    \I__3586\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20584\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__20584\,
            I => \N__20581\
        );

    \I__3584\ : Span4Mux_v
    port map (
            O => \N__20581\,
            I => \N__20578\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__20578\,
            I => \tok.n321\
        );

    \I__3582\ : InMux
    port map (
            O => \N__20575\,
            I => \N__20566\
        );

    \I__3581\ : InMux
    port map (
            O => \N__20574\,
            I => \N__20566\
        );

    \I__3580\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20566\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20563\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__20563\,
            I => \tok.n4_adj_640\
        );

    \I__3577\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20553\
        );

    \I__3576\ : InMux
    port map (
            O => \N__20559\,
            I => \N__20553\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__20558\,
            I => \N__20550\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__20553\,
            I => \N__20547\
        );

    \I__3573\ : InMux
    port map (
            O => \N__20550\,
            I => \N__20544\
        );

    \I__3572\ : Span4Mux_h
    port map (
            O => \N__20547\,
            I => \N__20541\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__20544\,
            I => \N__20538\
        );

    \I__3570\ : Span4Mux_v
    port map (
            O => \N__20541\,
            I => \N__20535\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__20538\,
            I => \tok.n4_adj_680\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__20535\,
            I => \tok.n4_adj_680\
        );

    \I__3567\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20527\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__20527\,
            I => \N__20524\
        );

    \I__3565\ : Span4Mux_v
    port map (
            O => \N__20524\,
            I => \N__20521\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__20521\,
            I => \tok.n239_adj_679\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__20518\,
            I => \tok.n238_adj_681_cascade_\
        );

    \I__3562\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20511\
        );

    \I__3561\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20508\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__20511\,
            I => \N__20505\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__20508\,
            I => \tok.n900\
        );

    \I__3558\ : Odrv12
    port map (
            O => \N__20505\,
            I => \tok.n900\
        );

    \I__3557\ : InMux
    port map (
            O => \N__20500\,
            I => \N__20497\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__20497\,
            I => \N__20494\
        );

    \I__3555\ : Span4Mux_v
    port map (
            O => \N__20494\,
            I => \N__20491\
        );

    \I__3554\ : Odrv4
    port map (
            O => \N__20491\,
            I => \tok.n317_adj_659\
        );

    \I__3553\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20485\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__20485\,
            I => \N__20482\
        );

    \I__3551\ : Odrv12
    port map (
            O => \N__20482\,
            I => \tok.n2663\
        );

    \I__3550\ : InMux
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__20476\,
            I => \tok.uart.sender_5\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__20473\,
            I => \tok.n2600_cascade_\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__20470\,
            I => \tok.n6610_cascade_\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__20467\,
            I => \N__20464\
        );

    \I__3545\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20461\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__20461\,
            I => \tok.n6344\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__20458\,
            I => \tok.n269_cascade_\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__20455\,
            I => \N__20452\
        );

    \I__3541\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20449\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__20449\,
            I => \tok.n4_adj_786\
        );

    \I__3539\ : InMux
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__20443\,
            I => \N__20440\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__20440\,
            I => \tok.n205_adj_789\
        );

    \I__3536\ : InMux
    port map (
            O => \N__20437\,
            I => \N__20434\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__20434\,
            I => \N__20430\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__20433\,
            I => \N__20427\
        );

    \I__3533\ : Span4Mux_v
    port map (
            O => \N__20430\,
            I => \N__20422\
        );

    \I__3532\ : InMux
    port map (
            O => \N__20427\,
            I => \N__20417\
        );

    \I__3531\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20417\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__20425\,
            I => \N__20413\
        );

    \I__3529\ : Span4Mux_h
    port map (
            O => \N__20422\,
            I => \N__20407\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__20417\,
            I => \N__20407\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__20416\,
            I => \N__20401\
        );

    \I__3526\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20397\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__20412\,
            I => \N__20393\
        );

    \I__3524\ : Span4Mux_h
    port map (
            O => \N__20407\,
            I => \N__20390\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__20406\,
            I => \N__20387\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__20405\,
            I => \N__20384\
        );

    \I__3521\ : InMux
    port map (
            O => \N__20404\,
            I => \N__20377\
        );

    \I__3520\ : InMux
    port map (
            O => \N__20401\,
            I => \N__20377\
        );

    \I__3519\ : InMux
    port map (
            O => \N__20400\,
            I => \N__20377\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__20397\,
            I => \N__20374\
        );

    \I__3517\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20369\
        );

    \I__3516\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20369\
        );

    \I__3515\ : Span4Mux_h
    port map (
            O => \N__20390\,
            I => \N__20366\
        );

    \I__3514\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20361\
        );

    \I__3513\ : InMux
    port map (
            O => \N__20384\,
            I => \N__20361\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__20377\,
            I => \N__20356\
        );

    \I__3511\ : Span4Mux_h
    port map (
            O => \N__20374\,
            I => \N__20356\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__20369\,
            I => \tok.n4_adj_635\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__20366\,
            I => \tok.n4_adj_635\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__20361\,
            I => \tok.n4_adj_635\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__20356\,
            I => \tok.n4_adj_635\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__20347\,
            I => \tok.n6341_cascade_\
        );

    \I__3505\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20336\
        );

    \I__3504\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20329\
        );

    \I__3503\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20329\
        );

    \I__3502\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20329\
        );

    \I__3501\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20326\
        );

    \I__3500\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20323\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__20336\,
            I => \N__20318\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__20329\,
            I => \N__20315\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__20326\,
            I => \N__20310\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__20323\,
            I => \N__20310\
        );

    \I__3495\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20307\
        );

    \I__3494\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20304\
        );

    \I__3493\ : Span4Mux_s3_v
    port map (
            O => \N__20318\,
            I => \N__20301\
        );

    \I__3492\ : Span4Mux_s3_v
    port map (
            O => \N__20315\,
            I => \N__20298\
        );

    \I__3491\ : Span4Mux_s3_v
    port map (
            O => \N__20310\,
            I => \N__20291\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__20307\,
            I => \N__20291\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__20304\,
            I => \N__20291\
        );

    \I__3488\ : Odrv4
    port map (
            O => \N__20301\,
            I => \tok.n170\
        );

    \I__3487\ : Odrv4
    port map (
            O => \N__20298\,
            I => \tok.n170\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__20291\,
            I => \tok.n170\
        );

    \I__3485\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20281\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__20281\,
            I => \tok.n197\
        );

    \I__3483\ : InMux
    port map (
            O => \N__20278\,
            I => \N__20275\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__20275\,
            I => \tok.n248\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__20272\,
            I => \tok.n6606_cascade_\
        );

    \I__3480\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20266\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__20266\,
            I => \tok.n200\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__20263\,
            I => \tok.n6_cascade_\
        );

    \I__3477\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20253\
        );

    \I__3476\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20253\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__20258\,
            I => \N__20250\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__20253\,
            I => \N__20245\
        );

    \I__3473\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20242\
        );

    \I__3472\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20239\
        );

    \I__3471\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20235\
        );

    \I__3470\ : Span4Mux_h
    port map (
            O => \N__20245\,
            I => \N__20230\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__20242\,
            I => \N__20230\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__20239\,
            I => \N__20227\
        );

    \I__3467\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20223\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__20235\,
            I => \N__20216\
        );

    \I__3465\ : Span4Mux_v
    port map (
            O => \N__20230\,
            I => \N__20216\
        );

    \I__3464\ : Span4Mux_h
    port map (
            O => \N__20227\,
            I => \N__20216\
        );

    \I__3463\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20213\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__20223\,
            I => \N__20208\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__20216\,
            I => \N__20208\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__20213\,
            I => \tok.S_12\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__20208\,
            I => \tok.S_12\
        );

    \I__3458\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20200\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__20200\,
            I => \N__20197\
        );

    \I__3456\ : Odrv12
    port map (
            O => \N__20197\,
            I => \tok.n200_adj_875\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__20194\,
            I => \tok.n6_adj_878_cascade_\
        );

    \I__3454\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20187\
        );

    \I__3453\ : InMux
    port map (
            O => \N__20190\,
            I => \N__20184\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__20187\,
            I => \N__20181\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__20184\,
            I => \N__20174\
        );

    \I__3450\ : Span4Mux_v
    port map (
            O => \N__20181\,
            I => \N__20170\
        );

    \I__3449\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20167\
        );

    \I__3448\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20164\
        );

    \I__3447\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20161\
        );

    \I__3446\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20158\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__20174\,
            I => \N__20155\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__20173\,
            I => \N__20152\
        );

    \I__3443\ : Span4Mux_h
    port map (
            O => \N__20170\,
            I => \N__20145\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__20167\,
            I => \N__20145\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__20164\,
            I => \N__20145\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__20161\,
            I => \N__20142\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__20158\,
            I => \N__20139\
        );

    \I__3438\ : Span4Mux_h
    port map (
            O => \N__20155\,
            I => \N__20136\
        );

    \I__3437\ : InMux
    port map (
            O => \N__20152\,
            I => \N__20133\
        );

    \I__3436\ : Span4Mux_h
    port map (
            O => \N__20145\,
            I => \N__20130\
        );

    \I__3435\ : Span4Mux_s2_v
    port map (
            O => \N__20142\,
            I => \N__20123\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__20139\,
            I => \N__20123\
        );

    \I__3433\ : Span4Mux_v
    port map (
            O => \N__20136\,
            I => \N__20123\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__20133\,
            I => \N__20120\
        );

    \I__3431\ : Span4Mux_v
    port map (
            O => \N__20130\,
            I => \N__20117\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__20123\,
            I => \tok.S_10\
        );

    \I__3429\ : Odrv12
    port map (
            O => \N__20120\,
            I => \tok.S_10\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__20117\,
            I => \tok.S_10\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__20110\,
            I => \tok.n4842_cascade_\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__20107\,
            I => \tok.n7451_cascade_\
        );

    \I__3425\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20101\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__20101\,
            I => \N__20098\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__20098\,
            I => \tok.n6616\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__20095\,
            I => \N__20091\
        );

    \I__3421\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20084\
        );

    \I__3420\ : InMux
    port map (
            O => \N__20091\,
            I => \N__20081\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__20090\,
            I => \N__20078\
        );

    \I__3418\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20071\
        );

    \I__3417\ : InMux
    port map (
            O => \N__20088\,
            I => \N__20071\
        );

    \I__3416\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20068\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__20084\,
            I => \N__20065\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20062\
        );

    \I__3413\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20059\
        );

    \I__3412\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20056\
        );

    \I__3411\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20053\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__20071\,
            I => \N__20050\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__20068\,
            I => \N__20047\
        );

    \I__3408\ : Span4Mux_v
    port map (
            O => \N__20065\,
            I => \N__20042\
        );

    \I__3407\ : Span4Mux_v
    port map (
            O => \N__20062\,
            I => \N__20042\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__20059\,
            I => \N__20037\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__20056\,
            I => \N__20037\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__20053\,
            I => \tok.S_2\
        );

    \I__3403\ : Odrv4
    port map (
            O => \N__20050\,
            I => \tok.S_2\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__20047\,
            I => \tok.S_2\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__20042\,
            I => \tok.S_2\
        );

    \I__3400\ : Odrv12
    port map (
            O => \N__20037\,
            I => \tok.S_2\
        );

    \I__3399\ : InMux
    port map (
            O => \N__20026\,
            I => \N__20023\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__20023\,
            I => \N__20020\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__20020\,
            I => \tok.n164\
        );

    \I__3396\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__20014\,
            I => \tok.n6597\
        );

    \I__3394\ : InMux
    port map (
            O => \N__20011\,
            I => \N__20008\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__20008\,
            I => \N__20005\
        );

    \I__3392\ : Span4Mux_v
    port map (
            O => \N__20005\,
            I => \N__20002\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__20002\,
            I => \tok.n4_adj_711\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__19999\,
            I => \N__19996\
        );

    \I__3389\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19993\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__19993\,
            I => \N__19990\
        );

    \I__3387\ : Odrv12
    port map (
            O => \N__19990\,
            I => \tok.n307\
        );

    \I__3386\ : InMux
    port map (
            O => \N__19987\,
            I => \N__19984\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__19984\,
            I => \N__19981\
        );

    \I__3384\ : Odrv12
    port map (
            O => \N__19981\,
            I => \tok.n6397\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__19978\,
            I => \tok.n242_cascade_\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__19975\,
            I => \N__19972\
        );

    \I__3381\ : InMux
    port map (
            O => \N__19972\,
            I => \N__19969\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__19969\,
            I => \tok.n6582\
        );

    \I__3379\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19963\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__19963\,
            I => \N__19960\
        );

    \I__3377\ : Span12Mux_s7_v
    port map (
            O => \N__19960\,
            I => \N__19957\
        );

    \I__3376\ : Odrv12
    port map (
            O => \N__19957\,
            I => \tok.table_wr_data_5\
        );

    \I__3375\ : CascadeMux
    port map (
            O => \N__19954\,
            I => \tok.n199_cascade_\
        );

    \I__3374\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19948\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__19948\,
            I => \tok.n262\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__19945\,
            I => \tok.n4_adj_648_cascade_\
        );

    \I__3371\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19939\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__19939\,
            I => \tok.n326\
        );

    \I__3369\ : InMux
    port map (
            O => \N__19936\,
            I => \N__19932\
        );

    \I__3368\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19929\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__19932\,
            I => \N__19926\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__19929\,
            I => \N__19923\
        );

    \I__3365\ : Span4Mux_v
    port map (
            O => \N__19926\,
            I => \N__19920\
        );

    \I__3364\ : Span4Mux_v
    port map (
            O => \N__19923\,
            I => \N__19917\
        );

    \I__3363\ : Span4Mux_h
    port map (
            O => \N__19920\,
            I => \N__19914\
        );

    \I__3362\ : Span4Mux_h
    port map (
            O => \N__19917\,
            I => \N__19911\
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__19914\,
            I => \tok.n234\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__19911\,
            I => \tok.n234\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__19906\,
            I => \N__19902\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__19905\,
            I => \N__19899\
        );

    \I__3357\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19896\
        );

    \I__3356\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19893\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__19896\,
            I => \N__19890\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__19893\,
            I => \N__19887\
        );

    \I__3353\ : Span4Mux_h
    port map (
            O => \N__19890\,
            I => \N__19884\
        );

    \I__3352\ : Span12Mux_s10_h
    port map (
            O => \N__19887\,
            I => \N__19881\
        );

    \I__3351\ : Span4Mux_v
    port map (
            O => \N__19884\,
            I => \N__19878\
        );

    \I__3350\ : Odrv12
    port map (
            O => \N__19881\,
            I => \tok.table_rd_5\
        );

    \I__3349\ : Odrv4
    port map (
            O => \N__19878\,
            I => \tok.table_rd_5\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__19873\,
            I => \tok.n286_cascade_\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__19870\,
            I => \N__19867\
        );

    \I__3346\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19864\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__19864\,
            I => \N__19861\
        );

    \I__3344\ : Span4Mux_h
    port map (
            O => \N__19861\,
            I => \N__19857\
        );

    \I__3343\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19854\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__19857\,
            I => \tok.n877\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__19854\,
            I => \tok.n877\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__19849\,
            I => \tok.n394_cascade_\
        );

    \I__3339\ : CascadeMux
    port map (
            O => \N__19846\,
            I => \N__19843\
        );

    \I__3338\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19840\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__19840\,
            I => \N__19837\
        );

    \I__3336\ : Span4Mux_h
    port map (
            O => \N__19837\,
            I => \N__19834\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__19834\,
            I => \tok.n6143\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__19831\,
            I => \N__19828\
        );

    \I__3333\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19825\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__19825\,
            I => \N__19822\
        );

    \I__3331\ : Span4Mux_h
    port map (
            O => \N__19822\,
            I => \N__19819\
        );

    \I__3330\ : Span4Mux_v
    port map (
            O => \N__19819\,
            I => \N__19816\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__19816\,
            I => \tok.tc_3\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__19813\,
            I => \N__19810\
        );

    \I__3327\ : InMux
    port map (
            O => \N__19810\,
            I => \N__19807\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__19807\,
            I => \N__19804\
        );

    \I__3325\ : Span4Mux_v
    port map (
            O => \N__19804\,
            I => \N__19801\
        );

    \I__3324\ : Span4Mux_h
    port map (
            O => \N__19801\,
            I => \N__19798\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__19798\,
            I => \tok.tc_1\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__19795\,
            I => \N__19791\
        );

    \I__3321\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19788\
        );

    \I__3320\ : InMux
    port map (
            O => \N__19791\,
            I => \N__19785\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__19788\,
            I => \N__19782\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19779\
        );

    \I__3317\ : Span4Mux_s3_v
    port map (
            O => \N__19782\,
            I => \N__19774\
        );

    \I__3316\ : Span4Mux_v
    port map (
            O => \N__19779\,
            I => \N__19774\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__19774\,
            I => n92_adj_897
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__19771\,
            I => \N__19768\
        );

    \I__3313\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19765\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__19765\,
            I => \N__19762\
        );

    \I__3311\ : Span4Mux_v
    port map (
            O => \N__19762\,
            I => \N__19759\
        );

    \I__3310\ : Span4Mux_h
    port map (
            O => \N__19759\,
            I => \N__19756\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__19756\,
            I => \tok.tc_0\
        );

    \I__3308\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19739\
        );

    \I__3307\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19739\
        );

    \I__3306\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19739\
        );

    \I__3305\ : InMux
    port map (
            O => \N__19750\,
            I => \N__19739\
        );

    \I__3304\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19732\
        );

    \I__3303\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19732\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__19739\,
            I => \N__19725\
        );

    \I__3301\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19720\
        );

    \I__3300\ : InMux
    port map (
            O => \N__19737\,
            I => \N__19720\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__19732\,
            I => \N__19713\
        );

    \I__3298\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19708\
        );

    \I__3297\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19708\
        );

    \I__3296\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19703\
        );

    \I__3295\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19703\
        );

    \I__3294\ : Span4Mux_h
    port map (
            O => \N__19725\,
            I => \N__19698\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__19720\,
            I => \N__19698\
        );

    \I__3292\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19689\
        );

    \I__3291\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19689\
        );

    \I__3290\ : InMux
    port map (
            O => \N__19717\,
            I => \N__19689\
        );

    \I__3289\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19689\
        );

    \I__3288\ : Span4Mux_v
    port map (
            O => \N__19713\,
            I => \N__19686\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__19708\,
            I => \N__19681\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19681\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__19698\,
            I => \N__19676\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__19689\,
            I => \N__19676\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__19686\,
            I => \stall_\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__19681\,
            I => \stall_\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__19676\,
            I => \stall_\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__19669\,
            I => \N__19666\
        );

    \I__3279\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19663\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__19663\,
            I => \N__19660\
        );

    \I__3277\ : Span4Mux_v
    port map (
            O => \N__19660\,
            I => \N__19657\
        );

    \I__3276\ : Span4Mux_v
    port map (
            O => \N__19657\,
            I => \N__19654\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__19654\,
            I => \tok.tc_2\
        );

    \I__3274\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19648\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__19648\,
            I => \tok.n6140\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__19645\,
            I => \tok.n225_adj_678_cascade_\
        );

    \I__3271\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19639\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__19639\,
            I => \tok.n6351\
        );

    \I__3269\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19633\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__19633\,
            I => \tok.n6632\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__19630\,
            I => \tok.n7456_cascade_\
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__19627\,
            I => \N__19624\
        );

    \I__3265\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19621\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19618\
        );

    \I__3263\ : Span4Mux_v
    port map (
            O => \N__19618\,
            I => \N__19615\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__19615\,
            I => \N__19612\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__19612\,
            I => \tok.n176\
        );

    \I__3260\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19606\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__19606\,
            I => \N__19603\
        );

    \I__3258\ : Odrv12
    port map (
            O => \N__19603\,
            I => \tok.n8_adj_686\
        );

    \I__3257\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19597\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__19597\,
            I => \tok.n6622\
        );

    \I__3255\ : CascadeMux
    port map (
            O => \N__19594\,
            I => \tok.n237_adj_724_cascade_\
        );

    \I__3254\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19588\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__19588\,
            I => \N__19585\
        );

    \I__3252\ : Span4Mux_v
    port map (
            O => \N__19585\,
            I => \N__19582\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__19582\,
            I => \tok.n4893\
        );

    \I__3250\ : InMux
    port map (
            O => \N__19579\,
            I => \N__19576\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__19576\,
            I => \tok.n286\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__19573\,
            I => \tok.ram.n6260_cascade_\
        );

    \I__3247\ : InMux
    port map (
            O => \N__19570\,
            I => \N__19567\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__19567\,
            I => \tok.n6295\
        );

    \I__3245\ : CascadeMux
    port map (
            O => \N__19564\,
            I => \tok.n1565_cascade_\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__19561\,
            I => \tok.n13_adj_757_cascade_\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__19558\,
            I => \n10_adj_906_cascade_\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__19555\,
            I => \N__19552\
        );

    \I__3241\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19549\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__19549\,
            I => \N__19546\
        );

    \I__3239\ : Span4Mux_v
    port map (
            O => \N__19546\,
            I => \N__19543\
        );

    \I__3238\ : Span4Mux_v
    port map (
            O => \N__19543\,
            I => \N__19540\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__19540\,
            I => \tok.tc_4\
        );

    \I__3236\ : InMux
    port map (
            O => \N__19537\,
            I => \N__19534\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__19534\,
            I => n10_adj_906
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__19531\,
            I => \tok.n324_cascade_\
        );

    \I__3233\ : InMux
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__19525\,
            I => \tok.n225_adj_678\
        );

    \I__3231\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19518\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__19521\,
            I => \N__19515\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__19518\,
            I => \N__19511\
        );

    \I__3228\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19508\
        );

    \I__3227\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19505\
        );

    \I__3226\ : Span4Mux_h
    port map (
            O => \N__19511\,
            I => \N__19500\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19497\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__19505\,
            I => \N__19494\
        );

    \I__3223\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19491\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__19503\,
            I => \N__19488\
        );

    \I__3221\ : Span4Mux_s0_v
    port map (
            O => \N__19500\,
            I => \N__19482\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__19497\,
            I => \N__19482\
        );

    \I__3219\ : Span4Mux_v
    port map (
            O => \N__19494\,
            I => \N__19477\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__19491\,
            I => \N__19477\
        );

    \I__3217\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19474\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__19487\,
            I => \N__19471\
        );

    \I__3215\ : Span4Mux_v
    port map (
            O => \N__19482\,
            I => \N__19463\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__19477\,
            I => \N__19463\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19463\
        );

    \I__3212\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19460\
        );

    \I__3211\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19457\
        );

    \I__3210\ : Span4Mux_h
    port map (
            O => \N__19463\,
            I => \N__19454\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__19460\,
            I => \N__19451\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__19457\,
            I => \N__19448\
        );

    \I__3207\ : Span4Mux_s1_h
    port map (
            O => \N__19454\,
            I => \N__19445\
        );

    \I__3206\ : Span4Mux_h
    port map (
            O => \N__19451\,
            I => \N__19442\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__19448\,
            I => \tok.S_11\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__19445\,
            I => \tok.S_11\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__19442\,
            I => \tok.S_11\
        );

    \I__3202\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19432\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__19432\,
            I => \N__19429\
        );

    \I__3200\ : Span4Mux_s1_v
    port map (
            O => \N__19429\,
            I => \N__19426\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__19426\,
            I => \tok.n197_adj_883\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__19423\,
            I => \N__19420\
        );

    \I__3197\ : InMux
    port map (
            O => \N__19420\,
            I => \N__19417\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__19417\,
            I => \tok.n248_adj_884\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__19414\,
            I => \tok.n83_adj_756_cascade_\
        );

    \I__3194\ : InMux
    port map (
            O => \N__19411\,
            I => \N__19408\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__19408\,
            I => \N__19405\
        );

    \I__3192\ : Span4Mux_s2_v
    port map (
            O => \N__19405\,
            I => \N__19402\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__19402\,
            I => \tok.n248_adj_827\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__19399\,
            I => \tok.n242_adj_828_cascade_\
        );

    \I__3189\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19393\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__19393\,
            I => \tok.n200_adj_829\
        );

    \I__3187\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19384\
        );

    \I__3186\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19384\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__19384\,
            I => \tok.n231\
        );

    \I__3184\ : InMux
    port map (
            O => \N__19381\,
            I => \N__19378\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__19378\,
            I => \N__19375\
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__19375\,
            I => \tok.n242_adj_885\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__19372\,
            I => \tok.n200_adj_886_cascade_\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__19369\,
            I => \tok.n6_adj_889_cascade_\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__19366\,
            I => \tok.n8_cascade_\
        );

    \I__3178\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19360\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__19360\,
            I => \N__19357\
        );

    \I__3176\ : Odrv12
    port map (
            O => \N__19357\,
            I => \tok.n6368\
        );

    \I__3175\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19351\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__19351\,
            I => \tok.n197_adj_668\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__19348\,
            I => \tok.n248_adj_669_cascade_\
        );

    \I__3172\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19342\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__19342\,
            I => \tok.n242_adj_670\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__19339\,
            I => \tok.n200_adj_671_cascade_\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__19336\,
            I => \N__19330\
        );

    \I__3168\ : InMux
    port map (
            O => \N__19335\,
            I => \N__19325\
        );

    \I__3167\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19325\
        );

    \I__3166\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19322\
        );

    \I__3165\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19317\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__19325\,
            I => \N__19314\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__19322\,
            I => \N__19311\
        );

    \I__3162\ : InMux
    port map (
            O => \N__19321\,
            I => \N__19308\
        );

    \I__3161\ : InMux
    port map (
            O => \N__19320\,
            I => \N__19305\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__19317\,
            I => \N__19301\
        );

    \I__3159\ : Span4Mux_v
    port map (
            O => \N__19314\,
            I => \N__19292\
        );

    \I__3158\ : Span4Mux_v
    port map (
            O => \N__19311\,
            I => \N__19292\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__19308\,
            I => \N__19292\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__19305\,
            I => \N__19292\
        );

    \I__3155\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19289\
        );

    \I__3154\ : Span4Mux_v
    port map (
            O => \N__19301\,
            I => \N__19286\
        );

    \I__3153\ : Span4Mux_v
    port map (
            O => \N__19292\,
            I => \N__19283\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__19289\,
            I => \N__19278\
        );

    \I__3151\ : Span4Mux_v
    port map (
            O => \N__19286\,
            I => \N__19278\
        );

    \I__3150\ : Span4Mux_h
    port map (
            O => \N__19283\,
            I => \N__19275\
        );

    \I__3149\ : Odrv4
    port map (
            O => \N__19278\,
            I => \tok.S_14\
        );

    \I__3148\ : Odrv4
    port map (
            O => \N__19275\,
            I => \tok.S_14\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__19270\,
            I => \tok.n6_adj_674_cascade_\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__19267\,
            I => \N__19264\
        );

    \I__3145\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19261\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__19261\,
            I => \N__19258\
        );

    \I__3143\ : Span4Mux_v
    port map (
            O => \N__19258\,
            I => \N__19255\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__19255\,
            I => \tok.table_rd_8\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__19252\,
            I => \N__19248\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__19251\,
            I => \N__19241\
        );

    \I__3139\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19237\
        );

    \I__3138\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19234\
        );

    \I__3137\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19231\
        );

    \I__3136\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19228\
        );

    \I__3135\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19225\
        );

    \I__3134\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19222\
        );

    \I__3133\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19219\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__19237\,
            I => \N__19215\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__19234\,
            I => \N__19209\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__19231\,
            I => \N__19209\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__19228\,
            I => \N__19206\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__19225\,
            I => \N__19199\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__19222\,
            I => \N__19199\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__19219\,
            I => \N__19199\
        );

    \I__3125\ : InMux
    port map (
            O => \N__19218\,
            I => \N__19196\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__19215\,
            I => \N__19193\
        );

    \I__3123\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19190\
        );

    \I__3122\ : Span4Mux_v
    port map (
            O => \N__19209\,
            I => \N__19187\
        );

    \I__3121\ : Span4Mux_s2_v
    port map (
            O => \N__19206\,
            I => \N__19180\
        );

    \I__3120\ : Span4Mux_v
    port map (
            O => \N__19199\,
            I => \N__19180\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__19196\,
            I => \N__19180\
        );

    \I__3118\ : Span4Mux_v
    port map (
            O => \N__19193\,
            I => \N__19177\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__19190\,
            I => \tok.n7269\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__19187\,
            I => \tok.n7269\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__19180\,
            I => \tok.n7269\
        );

    \I__3114\ : Odrv4
    port map (
            O => \N__19177\,
            I => \tok.n7269\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__19168\,
            I => \tok.n203_adj_822_cascade_\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__19165\,
            I => \tok.n212_adj_824_cascade_\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__19162\,
            I => \tok.n6457_cascade_\
        );

    \I__3110\ : InMux
    port map (
            O => \N__19159\,
            I => \N__19156\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__19156\,
            I => \N__19153\
        );

    \I__3108\ : Odrv12
    port map (
            O => \N__19153\,
            I => \tok.n208_adj_857\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__19150\,
            I => \N__19147\
        );

    \I__3106\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19144\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__19144\,
            I => \tok.n6328\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__19141\,
            I => \N__19138\
        );

    \I__3103\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19135\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__19135\,
            I => \N__19132\
        );

    \I__3101\ : Odrv12
    port map (
            O => \N__19132\,
            I => \tok.n250\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__19129\,
            I => \tok.n190_adj_774_cascade_\
        );

    \I__3099\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19123\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__19123\,
            I => \N__19120\
        );

    \I__3097\ : Span4Mux_h
    port map (
            O => \N__19120\,
            I => \N__19117\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__19117\,
            I => \tok.n6514\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__19114\,
            I => \tok.n833_cascade_\
        );

    \I__3094\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19108\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__19105\,
            I => \tok.n6515\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__19102\,
            I => \tok.n6534_cascade_\
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__19099\,
            I => \tok.n252_adj_783_cascade_\
        );

    \I__3089\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19093\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__19093\,
            I => \tok.n255_adj_775\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__19090\,
            I => \N__19087\
        );

    \I__3086\ : InMux
    port map (
            O => \N__19087\,
            I => \N__19084\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__19084\,
            I => \tok.n190_adj_774\
        );

    \I__3084\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19078\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__19078\,
            I => \tok.n258_adj_780\
        );

    \I__3082\ : InMux
    port map (
            O => \N__19075\,
            I => \N__19072\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__19072\,
            I => \tok.n177_adj_779\
        );

    \I__3080\ : InMux
    port map (
            O => \N__19069\,
            I => \N__19066\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__19066\,
            I => \tok.n22_adj_847\
        );

    \I__3078\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19060\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__19060\,
            I => \tok.n27_adj_782\
        );

    \I__3076\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19054\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__19054\,
            I => \tok.n298\
        );

    \I__3074\ : InMux
    port map (
            O => \N__19051\,
            I => \N__19048\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__19048\,
            I => \tok.n161_adj_870\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__19045\,
            I => \tok.n6429_cascade_\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__19042\,
            I => \tok.n197_adj_872_cascade_\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__19039\,
            I => \N__19036\
        );

    \I__3069\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19033\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__19033\,
            I => \N__19030\
        );

    \I__3067\ : Span4Mux_s3_h
    port map (
            O => \N__19030\,
            I => \N__19027\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__19027\,
            I => \tok.n248_adj_873\
        );

    \I__3065\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19021\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__19021\,
            I => \tok.n296\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__19018\,
            I => \tok.n6400_cascade_\
        );

    \I__3062\ : InMux
    port map (
            O => \N__19015\,
            I => \N__19012\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__19012\,
            I => \tok.n161\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__19009\,
            I => \N__19006\
        );

    \I__3059\ : InMux
    port map (
            O => \N__19006\,
            I => \N__19003\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__19003\,
            I => \N__19000\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__19000\,
            I => \tok.n6406\
        );

    \I__3056\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18994\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__18994\,
            I => \tok.n6415\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__18991\,
            I => \tok.n161_adj_882_cascade_\
        );

    \I__3053\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18985\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__18985\,
            I => \tok.n26_adj_781\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__18982\,
            I => \tok.n28_adj_778_cascade_\
        );

    \I__3050\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18976\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__18976\,
            I => \tok.n25_adj_788\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__18973\,
            I => \N__18969\
        );

    \I__3047\ : InMux
    port map (
            O => \N__18972\,
            I => \N__18964\
        );

    \I__3046\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18964\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__18964\,
            I => \N__18959\
        );

    \I__3044\ : InMux
    port map (
            O => \N__18963\,
            I => \N__18956\
        );

    \I__3043\ : InMux
    port map (
            O => \N__18962\,
            I => \N__18952\
        );

    \I__3042\ : Span4Mux_s3_v
    port map (
            O => \N__18959\,
            I => \N__18945\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__18956\,
            I => \N__18945\
        );

    \I__3040\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18942\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__18952\,
            I => \N__18939\
        );

    \I__3038\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18936\
        );

    \I__3037\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18933\
        );

    \I__3036\ : Sp12to4
    port map (
            O => \N__18945\,
            I => \N__18928\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__18942\,
            I => \N__18928\
        );

    \I__3034\ : Span4Mux_s3_v
    port map (
            O => \N__18939\,
            I => \N__18923\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__18936\,
            I => \N__18923\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__18933\,
            I => \N__18920\
        );

    \I__3031\ : Span12Mux_s6_v
    port map (
            O => \N__18928\,
            I => \N__18917\
        );

    \I__3030\ : Span4Mux_v
    port map (
            O => \N__18923\,
            I => \N__18912\
        );

    \I__3029\ : Span4Mux_h
    port map (
            O => \N__18920\,
            I => \N__18912\
        );

    \I__3028\ : Odrv12
    port map (
            O => \N__18917\,
            I => \tok.S_15\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__18912\,
            I => \tok.S_15\
        );

    \I__3026\ : InMux
    port map (
            O => \N__18907\,
            I => \N__18904\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__18904\,
            I => \tok.n6634\
        );

    \I__3024\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18898\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__18898\,
            I => \tok.n23_adj_848\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__18895\,
            I => \tok.n21_adj_849_cascade_\
        );

    \I__3021\ : InMux
    port map (
            O => \N__18892\,
            I => \N__18889\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__18889\,
            I => \tok.n24_adj_846\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__18886\,
            I => \N__18883\
        );

    \I__3018\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18880\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__18880\,
            I => \N__18877\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__18877\,
            I => \tok.n30_adj_852\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__18874\,
            I => \N__18871\
        );

    \I__3014\ : InMux
    port map (
            O => \N__18871\,
            I => \N__18868\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__18868\,
            I => \tok.n323\
        );

    \I__3012\ : InMux
    port map (
            O => \N__18865\,
            I => \N__18862\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__18862\,
            I => \tok.n163\
        );

    \I__3010\ : InMux
    port map (
            O => \N__18859\,
            I => \N__18856\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__18856\,
            I => \tok.n256_adj_862\
        );

    \I__3008\ : InMux
    port map (
            O => \N__18853\,
            I => \N__18850\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__18850\,
            I => \N__18847\
        );

    \I__3006\ : Span4Mux_v
    port map (
            O => \N__18847\,
            I => \N__18844\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__18844\,
            I => \N__18841\
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__18841\,
            I => \tok.n5_adj_871\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__18838\,
            I => \tok.n6_adj_868_cascade_\
        );

    \I__3002\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18829\
        );

    \I__3001\ : InMux
    port map (
            O => \N__18834\,
            I => \N__18823\
        );

    \I__3000\ : InMux
    port map (
            O => \N__18833\,
            I => \N__18823\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__18832\,
            I => \N__18820\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__18829\,
            I => \N__18817\
        );

    \I__2997\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18814\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__18823\,
            I => \N__18809\
        );

    \I__2995\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18806\
        );

    \I__2994\ : Span4Mux_v
    port map (
            O => \N__18817\,
            I => \N__18801\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__18814\,
            I => \N__18801\
        );

    \I__2992\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18798\
        );

    \I__2991\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18795\
        );

    \I__2990\ : Span4Mux_v
    port map (
            O => \N__18809\,
            I => \N__18792\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__18806\,
            I => \N__18789\
        );

    \I__2988\ : Span4Mux_v
    port map (
            O => \N__18801\,
            I => \N__18786\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__18798\,
            I => \N__18783\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__18795\,
            I => \N__18776\
        );

    \I__2985\ : Span4Mux_h
    port map (
            O => \N__18792\,
            I => \N__18776\
        );

    \I__2984\ : Span4Mux_h
    port map (
            O => \N__18789\,
            I => \N__18776\
        );

    \I__2983\ : Span4Mux_h
    port map (
            O => \N__18786\,
            I => \N__18773\
        );

    \I__2982\ : Odrv12
    port map (
            O => \N__18783\,
            I => \S_0\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__18776\,
            I => \S_0\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__18773\,
            I => \S_0\
        );

    \I__2979\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18763\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__18763\,
            I => \N__18760\
        );

    \I__2977\ : Span4Mux_h
    port map (
            O => \N__18760\,
            I => \N__18757\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__18757\,
            I => \tok.n28\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__18754\,
            I => \N__18750\
        );

    \I__2974\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18745\
        );

    \I__2973\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18745\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__18745\,
            I => \N__18742\
        );

    \I__2971\ : Span4Mux_v
    port map (
            O => \N__18742\,
            I => \N__18739\
        );

    \I__2970\ : Span4Mux_h
    port map (
            O => \N__18739\,
            I => \N__18736\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__18736\,
            I => \tok.key_rd_11\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__18733\,
            I => \N__18730\
        );

    \I__2967\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18724\
        );

    \I__2966\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18724\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__18724\,
            I => \N__18721\
        );

    \I__2964\ : Span4Mux_h
    port map (
            O => \N__18721\,
            I => \N__18718\
        );

    \I__2963\ : Odrv4
    port map (
            O => \N__18718\,
            I => \tok.key_rd_14\
        );

    \I__2962\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18712\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__18712\,
            I => \N__18709\
        );

    \I__2960\ : Odrv12
    port map (
            O => \N__18709\,
            I => \tok.n23_adj_638\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__18706\,
            I => \N__18702\
        );

    \I__2958\ : InMux
    port map (
            O => \N__18705\,
            I => \N__18697\
        );

    \I__2957\ : InMux
    port map (
            O => \N__18702\,
            I => \N__18697\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__18697\,
            I => \N__18694\
        );

    \I__2955\ : Span4Mux_v
    port map (
            O => \N__18694\,
            I => \N__18691\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__18691\,
            I => \tok.key_rd_15\
        );

    \I__2953\ : InMux
    port map (
            O => \N__18688\,
            I => \N__18682\
        );

    \I__2952\ : InMux
    port map (
            O => \N__18687\,
            I => \N__18682\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__18682\,
            I => \N__18679\
        );

    \I__2950\ : Span4Mux_h
    port map (
            O => \N__18679\,
            I => \N__18676\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__18676\,
            I => \tok.key_rd_9\
        );

    \I__2948\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18670\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__18670\,
            I => \N__18667\
        );

    \I__2946\ : Odrv12
    port map (
            O => \N__18667\,
            I => \tok.n24\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__18664\,
            I => \tok.n283_cascade_\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__18661\,
            I => \tok.n223_cascade_\
        );

    \I__2943\ : InMux
    port map (
            O => \N__18658\,
            I => \N__18655\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__18655\,
            I => \tok.n4_adj_752\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__18652\,
            I => \tok.n6586_cascade_\
        );

    \I__2940\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18646\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__18646\,
            I => \tok.n226_adj_744\
        );

    \I__2938\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18640\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__18640\,
            I => \tok.n254\
        );

    \I__2936\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18634\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__18634\,
            I => \N__18631\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__18631\,
            I => \tok.n319\
        );

    \I__2933\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18625\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__18625\,
            I => \N__18622\
        );

    \I__2931\ : Span4Mux_h
    port map (
            O => \N__18622\,
            I => \N__18619\
        );

    \I__2930\ : Odrv4
    port map (
            O => \N__18619\,
            I => \tok.n6326\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__18616\,
            I => \tok.n387_cascade_\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__18613\,
            I => \tok.n254_adj_860_cascade_\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__18610\,
            I => \N__18607\
        );

    \I__2926\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18603\
        );

    \I__2925\ : InMux
    port map (
            O => \N__18606\,
            I => \N__18600\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__18603\,
            I => \N__18597\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__18600\,
            I => \tok.n5_adj_675\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__18597\,
            I => \tok.n5_adj_675\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__18592\,
            I => \tok.n6205_cascade_\
        );

    \I__2920\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18578\
        );

    \I__2919\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18573\
        );

    \I__2918\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18573\
        );

    \I__2917\ : InMux
    port map (
            O => \N__18586\,
            I => \N__18570\
        );

    \I__2916\ : InMux
    port map (
            O => \N__18585\,
            I => \N__18566\
        );

    \I__2915\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18559\
        );

    \I__2914\ : InMux
    port map (
            O => \N__18583\,
            I => \N__18556\
        );

    \I__2913\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18551\
        );

    \I__2912\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18551\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__18578\,
            I => \N__18543\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18543\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__18570\,
            I => \N__18543\
        );

    \I__2908\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18540\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__18566\,
            I => \N__18537\
        );

    \I__2906\ : InMux
    port map (
            O => \N__18565\,
            I => \N__18530\
        );

    \I__2905\ : InMux
    port map (
            O => \N__18564\,
            I => \N__18530\
        );

    \I__2904\ : InMux
    port map (
            O => \N__18563\,
            I => \N__18530\
        );

    \I__2903\ : InMux
    port map (
            O => \N__18562\,
            I => \N__18527\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__18559\,
            I => \N__18524\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__18556\,
            I => \N__18519\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__18551\,
            I => \N__18519\
        );

    \I__2899\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18516\
        );

    \I__2898\ : Span4Mux_v
    port map (
            O => \N__18543\,
            I => \N__18511\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__18540\,
            I => \N__18511\
        );

    \I__2896\ : Span4Mux_s0_v
    port map (
            O => \N__18537\,
            I => \N__18506\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__18530\,
            I => \N__18506\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__18527\,
            I => \N__18503\
        );

    \I__2893\ : Span4Mux_s3_v
    port map (
            O => \N__18524\,
            I => \N__18496\
        );

    \I__2892\ : Span4Mux_v
    port map (
            O => \N__18519\,
            I => \N__18496\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__18516\,
            I => \N__18496\
        );

    \I__2890\ : Span4Mux_h
    port map (
            O => \N__18511\,
            I => \N__18491\
        );

    \I__2889\ : Span4Mux_v
    port map (
            O => \N__18506\,
            I => \N__18491\
        );

    \I__2888\ : Span4Mux_s3_v
    port map (
            O => \N__18503\,
            I => \N__18486\
        );

    \I__2887\ : Span4Mux_h
    port map (
            O => \N__18496\,
            I => \N__18486\
        );

    \I__2886\ : Odrv4
    port map (
            O => \N__18491\,
            I => \tok.n270\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__18486\,
            I => \tok.n270\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__18481\,
            I => \tok.n270_cascade_\
        );

    \I__2883\ : InMux
    port map (
            O => \N__18478\,
            I => \N__18475\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__18475\,
            I => \N__18472\
        );

    \I__2881\ : Span4Mux_v
    port map (
            O => \N__18472\,
            I => \N__18469\
        );

    \I__2880\ : Span4Mux_h
    port map (
            O => \N__18469\,
            I => \N__18465\
        );

    \I__2879\ : InMux
    port map (
            O => \N__18468\,
            I => \N__18462\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__18465\,
            I => \tok.A_stk.tail_18\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__18462\,
            I => \tok.A_stk.tail_18\
        );

    \I__2876\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18424\
        );

    \I__2875\ : InMux
    port map (
            O => \N__18456\,
            I => \N__18424\
        );

    \I__2874\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18424\
        );

    \I__2873\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18424\
        );

    \I__2872\ : InMux
    port map (
            O => \N__18453\,
            I => \N__18424\
        );

    \I__2871\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18424\
        );

    \I__2870\ : InMux
    port map (
            O => \N__18451\,
            I => \N__18424\
        );

    \I__2869\ : InMux
    port map (
            O => \N__18450\,
            I => \N__18409\
        );

    \I__2868\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18409\
        );

    \I__2867\ : InMux
    port map (
            O => \N__18448\,
            I => \N__18409\
        );

    \I__2866\ : InMux
    port map (
            O => \N__18447\,
            I => \N__18409\
        );

    \I__2865\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18409\
        );

    \I__2864\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18409\
        );

    \I__2863\ : InMux
    port map (
            O => \N__18444\,
            I => \N__18409\
        );

    \I__2862\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18398\
        );

    \I__2861\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18398\
        );

    \I__2860\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18398\
        );

    \I__2859\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18398\
        );

    \I__2858\ : InMux
    port map (
            O => \N__18439\,
            I => \N__18398\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__18424\,
            I => \N__18338\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__18409\,
            I => \N__18338\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__18398\,
            I => \N__18338\
        );

    \I__2854\ : InMux
    port map (
            O => \N__18397\,
            I => \N__18323\
        );

    \I__2853\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18323\
        );

    \I__2852\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18323\
        );

    \I__2851\ : InMux
    port map (
            O => \N__18394\,
            I => \N__18323\
        );

    \I__2850\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18323\
        );

    \I__2849\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18323\
        );

    \I__2848\ : InMux
    port map (
            O => \N__18391\,
            I => \N__18323\
        );

    \I__2847\ : InMux
    port map (
            O => \N__18390\,
            I => \N__18299\
        );

    \I__2846\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18299\
        );

    \I__2845\ : InMux
    port map (
            O => \N__18388\,
            I => \N__18299\
        );

    \I__2844\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18299\
        );

    \I__2843\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18299\
        );

    \I__2842\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18299\
        );

    \I__2841\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18299\
        );

    \I__2840\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18299\
        );

    \I__2839\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18282\
        );

    \I__2838\ : InMux
    port map (
            O => \N__18381\,
            I => \N__18282\
        );

    \I__2837\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18282\
        );

    \I__2836\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18282\
        );

    \I__2835\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18282\
        );

    \I__2834\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18282\
        );

    \I__2833\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18282\
        );

    \I__2832\ : InMux
    port map (
            O => \N__18375\,
            I => \N__18282\
        );

    \I__2831\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18277\
        );

    \I__2830\ : InMux
    port map (
            O => \N__18373\,
            I => \N__18277\
        );

    \I__2829\ : InMux
    port map (
            O => \N__18372\,
            I => \N__18260\
        );

    \I__2828\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18260\
        );

    \I__2827\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18260\
        );

    \I__2826\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18260\
        );

    \I__2825\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18260\
        );

    \I__2824\ : InMux
    port map (
            O => \N__18367\,
            I => \N__18260\
        );

    \I__2823\ : InMux
    port map (
            O => \N__18366\,
            I => \N__18260\
        );

    \I__2822\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18260\
        );

    \I__2821\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18255\
        );

    \I__2820\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18255\
        );

    \I__2819\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18238\
        );

    \I__2818\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18238\
        );

    \I__2817\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18238\
        );

    \I__2816\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18238\
        );

    \I__2815\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18238\
        );

    \I__2814\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18238\
        );

    \I__2813\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18238\
        );

    \I__2812\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18223\
        );

    \I__2811\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18223\
        );

    \I__2810\ : InMux
    port map (
            O => \N__18353\,
            I => \N__18223\
        );

    \I__2809\ : InMux
    port map (
            O => \N__18352\,
            I => \N__18223\
        );

    \I__2808\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18223\
        );

    \I__2807\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18223\
        );

    \I__2806\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18223\
        );

    \I__2805\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18220\
        );

    \I__2804\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18209\
        );

    \I__2803\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18209\
        );

    \I__2802\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18209\
        );

    \I__2801\ : Span4Mux_s3_v
    port map (
            O => \N__18338\,
            I => \N__18204\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__18323\,
            I => \N__18204\
        );

    \I__2799\ : InMux
    port map (
            O => \N__18322\,
            I => \N__18152\
        );

    \I__2798\ : InMux
    port map (
            O => \N__18321\,
            I => \N__18152\
        );

    \I__2797\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18152\
        );

    \I__2796\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18152\
        );

    \I__2795\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18152\
        );

    \I__2794\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18152\
        );

    \I__2793\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18152\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__18299\,
            I => \N__18145\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__18282\,
            I => \N__18145\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__18277\,
            I => \N__18145\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__18260\,
            I => \N__18140\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__18255\,
            I => \N__18140\
        );

    \I__2787\ : InMux
    port map (
            O => \N__18254\,
            I => \N__18137\
        );

    \I__2786\ : InMux
    port map (
            O => \N__18253\,
            I => \N__18134\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__18238\,
            I => \N__18127\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__18223\,
            I => \N__18127\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__18220\,
            I => \N__18127\
        );

    \I__2782\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18118\
        );

    \I__2781\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18118\
        );

    \I__2780\ : InMux
    port map (
            O => \N__18217\,
            I => \N__18118\
        );

    \I__2779\ : InMux
    port map (
            O => \N__18216\,
            I => \N__18118\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18108\
        );

    \I__2777\ : Span4Mux_h
    port map (
            O => \N__18204\,
            I => \N__18108\
        );

    \I__2776\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18101\
        );

    \I__2775\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18101\
        );

    \I__2774\ : InMux
    port map (
            O => \N__18201\,
            I => \N__18101\
        );

    \I__2773\ : InMux
    port map (
            O => \N__18200\,
            I => \N__18088\
        );

    \I__2772\ : InMux
    port map (
            O => \N__18199\,
            I => \N__18088\
        );

    \I__2771\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18088\
        );

    \I__2770\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18088\
        );

    \I__2769\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18088\
        );

    \I__2768\ : InMux
    port map (
            O => \N__18195\,
            I => \N__18088\
        );

    \I__2767\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18073\
        );

    \I__2766\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18073\
        );

    \I__2765\ : InMux
    port map (
            O => \N__18192\,
            I => \N__18073\
        );

    \I__2764\ : InMux
    port map (
            O => \N__18191\,
            I => \N__18073\
        );

    \I__2763\ : InMux
    port map (
            O => \N__18190\,
            I => \N__18073\
        );

    \I__2762\ : InMux
    port map (
            O => \N__18189\,
            I => \N__18073\
        );

    \I__2761\ : InMux
    port map (
            O => \N__18188\,
            I => \N__18073\
        );

    \I__2760\ : InMux
    port map (
            O => \N__18187\,
            I => \N__18058\
        );

    \I__2759\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18058\
        );

    \I__2758\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18058\
        );

    \I__2757\ : InMux
    port map (
            O => \N__18184\,
            I => \N__18058\
        );

    \I__2756\ : InMux
    port map (
            O => \N__18183\,
            I => \N__18058\
        );

    \I__2755\ : InMux
    port map (
            O => \N__18182\,
            I => \N__18058\
        );

    \I__2754\ : InMux
    port map (
            O => \N__18181\,
            I => \N__18058\
        );

    \I__2753\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18045\
        );

    \I__2752\ : InMux
    port map (
            O => \N__18179\,
            I => \N__18045\
        );

    \I__2751\ : InMux
    port map (
            O => \N__18178\,
            I => \N__18045\
        );

    \I__2750\ : InMux
    port map (
            O => \N__18177\,
            I => \N__18045\
        );

    \I__2749\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18045\
        );

    \I__2748\ : InMux
    port map (
            O => \N__18175\,
            I => \N__18045\
        );

    \I__2747\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18028\
        );

    \I__2746\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18028\
        );

    \I__2745\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18028\
        );

    \I__2744\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18028\
        );

    \I__2743\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18028\
        );

    \I__2742\ : InMux
    port map (
            O => \N__18169\,
            I => \N__18028\
        );

    \I__2741\ : InMux
    port map (
            O => \N__18168\,
            I => \N__18028\
        );

    \I__2740\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18028\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__18152\,
            I => \N__18021\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__18145\,
            I => \N__18021\
        );

    \I__2737\ : Span4Mux_s1_v
    port map (
            O => \N__18140\,
            I => \N__18021\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__18137\,
            I => \N__18016\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__18134\,
            I => \N__18016\
        );

    \I__2734\ : Span4Mux_v
    port map (
            O => \N__18127\,
            I => \N__18011\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__18118\,
            I => \N__18011\
        );

    \I__2732\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18008\
        );

    \I__2731\ : InMux
    port map (
            O => \N__18116\,
            I => \N__17999\
        );

    \I__2730\ : InMux
    port map (
            O => \N__18115\,
            I => \N__17999\
        );

    \I__2729\ : InMux
    port map (
            O => \N__18114\,
            I => \N__17999\
        );

    \I__2728\ : InMux
    port map (
            O => \N__18113\,
            I => \N__17999\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__18108\,
            I => \A_stk_delta_1\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__18101\,
            I => \A_stk_delta_1\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__18088\,
            I => \A_stk_delta_1\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__18073\,
            I => \A_stk_delta_1\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__18058\,
            I => \A_stk_delta_1\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__18045\,
            I => \A_stk_delta_1\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__18028\,
            I => \A_stk_delta_1\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__18021\,
            I => \A_stk_delta_1\
        );

    \I__2719\ : Odrv12
    port map (
            O => \N__18016\,
            I => \A_stk_delta_1\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__18011\,
            I => \A_stk_delta_1\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__18008\,
            I => \A_stk_delta_1\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__17999\,
            I => \A_stk_delta_1\
        );

    \I__2715\ : InMux
    port map (
            O => \N__17974\,
            I => \N__17971\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__17971\,
            I => \N__17968\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__17968\,
            I => \N__17964\
        );

    \I__2712\ : InMux
    port map (
            O => \N__17967\,
            I => \N__17961\
        );

    \I__2711\ : Odrv4
    port map (
            O => \N__17964\,
            I => \tok.A_stk.tail_2\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__17961\,
            I => \tok.A_stk.tail_2\
        );

    \I__2709\ : CEMux
    port map (
            O => \N__17956\,
            I => \N__17952\
        );

    \I__2708\ : CEMux
    port map (
            O => \N__17955\,
            I => \N__17949\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__17952\,
            I => \N__17943\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__17949\,
            I => \N__17940\
        );

    \I__2705\ : CEMux
    port map (
            O => \N__17948\,
            I => \N__17937\
        );

    \I__2704\ : CEMux
    port map (
            O => \N__17947\,
            I => \N__17928\
        );

    \I__2703\ : CEMux
    port map (
            O => \N__17946\,
            I => \N__17920\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__17943\,
            I => \N__17916\
        );

    \I__2701\ : Span4Mux_h
    port map (
            O => \N__17940\,
            I => \N__17911\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__17937\,
            I => \N__17911\
        );

    \I__2699\ : CEMux
    port map (
            O => \N__17936\,
            I => \N__17908\
        );

    \I__2698\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17905\
        );

    \I__2697\ : CEMux
    port map (
            O => \N__17934\,
            I => \N__17897\
        );

    \I__2696\ : CEMux
    port map (
            O => \N__17933\,
            I => \N__17894\
        );

    \I__2695\ : CEMux
    port map (
            O => \N__17932\,
            I => \N__17891\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__17931\,
            I => \N__17888\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__17928\,
            I => \N__17881\
        );

    \I__2692\ : CEMux
    port map (
            O => \N__17927\,
            I => \N__17878\
        );

    \I__2691\ : CEMux
    port map (
            O => \N__17926\,
            I => \N__17875\
        );

    \I__2690\ : CEMux
    port map (
            O => \N__17925\,
            I => \N__17871\
        );

    \I__2689\ : CEMux
    port map (
            O => \N__17924\,
            I => \N__17868\
        );

    \I__2688\ : CEMux
    port map (
            O => \N__17923\,
            I => \N__17865\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__17920\,
            I => \N__17862\
        );

    \I__2686\ : CEMux
    port map (
            O => \N__17919\,
            I => \N__17859\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__17916\,
            I => \N__17852\
        );

    \I__2684\ : Span4Mux_v
    port map (
            O => \N__17911\,
            I => \N__17852\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__17908\,
            I => \N__17852\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__17905\,
            I => \N__17849\
        );

    \I__2681\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17846\
        );

    \I__2680\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17841\
        );

    \I__2679\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17841\
        );

    \I__2678\ : CEMux
    port map (
            O => \N__17901\,
            I => \N__17838\
        );

    \I__2677\ : CEMux
    port map (
            O => \N__17900\,
            I => \N__17835\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__17897\,
            I => \N__17828\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__17894\,
            I => \N__17828\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__17891\,
            I => \N__17828\
        );

    \I__2673\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17823\
        );

    \I__2672\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17823\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__17886\,
            I => \N__17820\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__17885\,
            I => \N__17817\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__17884\,
            I => \N__17814\
        );

    \I__2668\ : Span4Mux_s2_v
    port map (
            O => \N__17881\,
            I => \N__17806\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__17878\,
            I => \N__17806\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__17875\,
            I => \N__17803\
        );

    \I__2665\ : CEMux
    port map (
            O => \N__17874\,
            I => \N__17800\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__17871\,
            I => \N__17795\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__17868\,
            I => \N__17795\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__17865\,
            I => \N__17792\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__17862\,
            I => \N__17787\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__17859\,
            I => \N__17787\
        );

    \I__2659\ : Span4Mux_s2_h
    port map (
            O => \N__17852\,
            I => \N__17782\
        );

    \I__2658\ : Span4Mux_s2_h
    port map (
            O => \N__17849\,
            I => \N__17782\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__17846\,
            I => \N__17779\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__17841\,
            I => \N__17776\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__17838\,
            I => \N__17767\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__17835\,
            I => \N__17767\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__17828\,
            I => \N__17767\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__17823\,
            I => \N__17767\
        );

    \I__2651\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17758\
        );

    \I__2650\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17758\
        );

    \I__2649\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17758\
        );

    \I__2648\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17758\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__17812\,
            I => \N__17754\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__17811\,
            I => \N__17750\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__17806\,
            I => \N__17746\
        );

    \I__2644\ : Span4Mux_h
    port map (
            O => \N__17803\,
            I => \N__17741\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__17800\,
            I => \N__17741\
        );

    \I__2642\ : Span4Mux_v
    port map (
            O => \N__17795\,
            I => \N__17734\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__17792\,
            I => \N__17734\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__17787\,
            I => \N__17734\
        );

    \I__2639\ : Span4Mux_v
    port map (
            O => \N__17782\,
            I => \N__17729\
        );

    \I__2638\ : Span4Mux_h
    port map (
            O => \N__17779\,
            I => \N__17729\
        );

    \I__2637\ : Span4Mux_h
    port map (
            O => \N__17776\,
            I => \N__17722\
        );

    \I__2636\ : Span4Mux_s1_v
    port map (
            O => \N__17767\,
            I => \N__17722\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17722\
        );

    \I__2634\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17719\
        );

    \I__2633\ : InMux
    port map (
            O => \N__17754\,
            I => \N__17710\
        );

    \I__2632\ : InMux
    port map (
            O => \N__17753\,
            I => \N__17710\
        );

    \I__2631\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17710\
        );

    \I__2630\ : InMux
    port map (
            O => \N__17749\,
            I => \N__17710\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__17746\,
            I => \rd_15__N_300\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__17741\,
            I => \rd_15__N_300\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__17734\,
            I => \rd_15__N_300\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__17729\,
            I => \rd_15__N_300\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__17722\,
            I => \rd_15__N_300\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__17719\,
            I => \rd_15__N_300\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__17710\,
            I => \rd_15__N_300\
        );

    \I__2622\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17692\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__17692\,
            I => n10_adj_905
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__17689\,
            I => \tok.n83_adj_764_cascade_\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__17686\,
            I => \tok.ram.n6277_cascade_\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__17683\,
            I => \n10_cascade_\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__17680\,
            I => \N__17677\
        );

    \I__2616\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17674\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__17674\,
            I => \N__17671\
        );

    \I__2614\ : Span4Mux_h
    port map (
            O => \N__17671\,
            I => \N__17668\
        );

    \I__2613\ : Span4Mux_v
    port map (
            O => \N__17668\,
            I => \N__17665\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__17665\,
            I => \tok.tc_7\
        );

    \I__2611\ : InMux
    port map (
            O => \N__17662\,
            I => \N__17659\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__17659\,
            I => \tok.n1635\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__17656\,
            I => \N__17653\
        );

    \I__2608\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17650\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__17650\,
            I => \tok.n6662\
        );

    \I__2606\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17644\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__17644\,
            I => \tok.n13_adj_790\
        );

    \I__2604\ : InMux
    port map (
            O => \N__17641\,
            I => \N__17638\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__17638\,
            I => n10
        );

    \I__2602\ : InMux
    port map (
            O => \N__17635\,
            I => \tok.n4817\
        );

    \I__2601\ : InMux
    port map (
            O => \N__17632\,
            I => \tok.n4818\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__17629\,
            I => \tok.n13_adj_760_cascade_\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__17626\,
            I => \n10_adj_905_cascade_\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__17623\,
            I => \N__17620\
        );

    \I__2597\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17617\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17614\
        );

    \I__2595\ : Span4Mux_v
    port map (
            O => \N__17614\,
            I => \N__17611\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__17611\,
            I => \N__17608\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__17608\,
            I => \tok.tc_5\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__17605\,
            I => \tok.ram.n6263_cascade_\
        );

    \I__2591\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17599\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__17599\,
            I => \tok.n1530\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__17596\,
            I => \tok.n83_adj_759_cascade_\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__17593\,
            I => \N__17590\
        );

    \I__2587\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17587\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__17587\,
            I => \tok.n6660\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__17584\,
            I => \tok.n6_adj_699_cascade_\
        );

    \I__2584\ : InMux
    port map (
            O => \N__17581\,
            I => \bfn_6_2_0_\
        );

    \I__2583\ : InMux
    port map (
            O => \N__17578\,
            I => \tok.n4812\
        );

    \I__2582\ : InMux
    port map (
            O => \N__17575\,
            I => \tok.n4813\
        );

    \I__2581\ : InMux
    port map (
            O => \N__17572\,
            I => \tok.n4814\
        );

    \I__2580\ : InMux
    port map (
            O => \N__17569\,
            I => \tok.n4815\
        );

    \I__2579\ : InMux
    port map (
            O => \N__17566\,
            I => \tok.n4816\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__17563\,
            I => \tok.n262_adj_858_cascade_\
        );

    \I__2577\ : InMux
    port map (
            O => \N__17560\,
            I => \N__17557\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__17557\,
            I => \N__17554\
        );

    \I__2575\ : Span12Mux_s7_v
    port map (
            O => \N__17554\,
            I => \N__17551\
        );

    \I__2574\ : Odrv12
    port map (
            O => \N__17551\,
            I => \tok.n268\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__17548\,
            I => \N__17545\
        );

    \I__2572\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17542\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__17542\,
            I => \N__17539\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__17539\,
            I => \tok.n6315\
        );

    \I__2569\ : DummyBuf
    port map (
            O => \N__17536\,
            I => \N__17532\
        );

    \I__2568\ : DummyBuf
    port map (
            O => \N__17535\,
            I => \N__17529\
        );

    \I__2567\ : InMux
    port map (
            O => \N__17532\,
            I => \N__17525\
        );

    \I__2566\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17522\
        );

    \I__2565\ : SRMux
    port map (
            O => \N__17528\,
            I => \N__17519\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__17525\,
            I => \N__17510\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__17522\,
            I => \N__17510\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__17519\,
            I => \N__17504\
        );

    \I__2561\ : SRMux
    port map (
            O => \N__17518\,
            I => \N__17501\
        );

    \I__2560\ : InMux
    port map (
            O => \N__17517\,
            I => \N__17498\
        );

    \I__2559\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17492\
        );

    \I__2558\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17492\
        );

    \I__2557\ : Span4Mux_s1_h
    port map (
            O => \N__17510\,
            I => \N__17489\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__17509\,
            I => \N__17486\
        );

    \I__2555\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17482\
        );

    \I__2554\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17479\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__17504\,
            I => \N__17472\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__17501\,
            I => \N__17472\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__17498\,
            I => \N__17472\
        );

    \I__2550\ : SRMux
    port map (
            O => \N__17497\,
            I => \N__17469\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__17492\,
            I => \N__17466\
        );

    \I__2548\ : Span4Mux_h
    port map (
            O => \N__17489\,
            I => \N__17463\
        );

    \I__2547\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17460\
        );

    \I__2546\ : InMux
    port map (
            O => \N__17485\,
            I => \N__17457\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__17482\,
            I => \N__17448\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__17479\,
            I => \N__17448\
        );

    \I__2543\ : Span4Mux_h
    port map (
            O => \N__17472\,
            I => \N__17448\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__17469\,
            I => \N__17448\
        );

    \I__2541\ : Span4Mux_v
    port map (
            O => \N__17466\,
            I => \N__17445\
        );

    \I__2540\ : Sp12to4
    port map (
            O => \N__17463\,
            I => \N__17440\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__17460\,
            I => \N__17440\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__17457\,
            I => \N__17437\
        );

    \I__2537\ : Span4Mux_v
    port map (
            O => \N__17448\,
            I => \N__17434\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__17445\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2535\ : Odrv12
    port map (
            O => \N__17440\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__17437\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__17434\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__17425\,
            I => \CONSTANT_ONE_NET_cascade_\
        );

    \I__2531\ : InMux
    port map (
            O => \N__17422\,
            I => \N__17418\
        );

    \I__2530\ : InMux
    port map (
            O => \N__17421\,
            I => \N__17415\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__17418\,
            I => \N__17409\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__17415\,
            I => \N__17409\
        );

    \I__2527\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17406\
        );

    \I__2526\ : Span12Mux_s5_v
    port map (
            O => \N__17409\,
            I => \N__17403\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__17406\,
            I => \tok.n239\
        );

    \I__2524\ : Odrv12
    port map (
            O => \N__17403\,
            I => \tok.n239\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__17398\,
            I => \N__17395\
        );

    \I__2522\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17392\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__17392\,
            I => \N__17389\
        );

    \I__2520\ : Span4Mux_s2_h
    port map (
            O => \N__17389\,
            I => \N__17386\
        );

    \I__2519\ : Span4Mux_h
    port map (
            O => \N__17386\,
            I => \N__17383\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__17383\,
            I => sender_2
        );

    \I__2517\ : InMux
    port map (
            O => \N__17380\,
            I => \N__17377\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__17377\,
            I => \N__17374\
        );

    \I__2515\ : Span4Mux_h
    port map (
            O => \N__17374\,
            I => \N__17371\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__17371\,
            I => \tok.n6347\
        );

    \I__2513\ : InMux
    port map (
            O => \N__17368\,
            I => \N__17365\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__17365\,
            I => \tok.n197_adj_693\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__17362\,
            I => \tok.n248_adj_694_cascade_\
        );

    \I__2510\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17356\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__17356\,
            I => \tok.n242_adj_695\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__17353\,
            I => \tok.n200_adj_696_cascade_\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__17350\,
            I => \tok.n200_adj_655_cascade_\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__17347\,
            I => \tok.n6_adj_658_cascade_\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__17344\,
            I => \tok.n6_adj_832_cascade_\
        );

    \I__2504\ : InMux
    port map (
            O => \N__17341\,
            I => \N__17338\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__17338\,
            I => \N__17335\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__17335\,
            I => \N__17332\
        );

    \I__2501\ : Span4Mux_s2_h
    port map (
            O => \N__17332\,
            I => \N__17329\
        );

    \I__2500\ : Odrv4
    port map (
            O => \N__17329\,
            I => \tok.n6383\
        );

    \I__2499\ : InMux
    port map (
            O => \N__17326\,
            I => \N__17323\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__17323\,
            I => \tok.n242_adj_654\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__17320\,
            I => \N__17315\
        );

    \I__2496\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17310\
        );

    \I__2495\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17307\
        );

    \I__2494\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17304\
        );

    \I__2493\ : InMux
    port map (
            O => \N__17314\,
            I => \N__17299\
        );

    \I__2492\ : InMux
    port map (
            O => \N__17313\,
            I => \N__17299\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__17310\,
            I => \N__17289\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__17307\,
            I => \N__17289\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__17304\,
            I => \N__17289\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__17299\,
            I => \N__17289\
        );

    \I__2487\ : InMux
    port map (
            O => \N__17298\,
            I => \N__17285\
        );

    \I__2486\ : Span4Mux_v
    port map (
            O => \N__17289\,
            I => \N__17282\
        );

    \I__2485\ : InMux
    port map (
            O => \N__17288\,
            I => \N__17279\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__17285\,
            I => \N__17276\
        );

    \I__2483\ : Span4Mux_h
    port map (
            O => \N__17282\,
            I => \N__17273\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__17279\,
            I => \tok.S_13\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__17276\,
            I => \tok.S_13\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__17273\,
            I => \tok.S_13\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__17266\,
            I => \N__17262\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__17265\,
            I => \N__17258\
        );

    \I__2477\ : InMux
    port map (
            O => \N__17262\,
            I => \N__17255\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__17261\,
            I => \N__17252\
        );

    \I__2475\ : InMux
    port map (
            O => \N__17258\,
            I => \N__17246\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__17255\,
            I => \N__17243\
        );

    \I__2473\ : InMux
    port map (
            O => \N__17252\,
            I => \N__17240\
        );

    \I__2472\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17235\
        );

    \I__2471\ : InMux
    port map (
            O => \N__17250\,
            I => \N__17235\
        );

    \I__2470\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17232\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__17246\,
            I => \N__17229\
        );

    \I__2468\ : Span4Mux_s3_v
    port map (
            O => \N__17243\,
            I => \N__17224\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__17240\,
            I => \N__17224\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__17235\,
            I => \N__17221\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__17232\,
            I => \N__17217\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__17229\,
            I => \N__17214\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__17224\,
            I => \N__17209\
        );

    \I__2462\ : Span4Mux_s3_v
    port map (
            O => \N__17221\,
            I => \N__17209\
        );

    \I__2461\ : InMux
    port map (
            O => \N__17220\,
            I => \N__17206\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__17217\,
            I => \N__17203\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__17214\,
            I => \N__17198\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__17209\,
            I => \N__17198\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__17206\,
            I => \tok.S_8\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__17203\,
            I => \tok.S_8\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__17198\,
            I => \tok.S_8\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__17191\,
            I => \tok.n14_adj_844_cascade_\
        );

    \I__2453\ : InMux
    port map (
            O => \N__17188\,
            I => \N__17185\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__17185\,
            I => \N__17182\
        );

    \I__2451\ : Odrv12
    port map (
            O => \N__17182\,
            I => \tok.n20_adj_845\
        );

    \I__2450\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17176\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__17176\,
            I => \tok.n26_adj_851\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__17173\,
            I => \tok.n6324_cascade_\
        );

    \I__2447\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17167\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__17167\,
            I => \tok.n6460\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__17164\,
            I => \N__17161\
        );

    \I__2444\ : InMux
    port map (
            O => \N__17161\,
            I => \N__17158\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__17158\,
            I => \tok.n161_adj_825\
        );

    \I__2442\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17152\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__17152\,
            I => \tok.n197_adj_826\
        );

    \I__2440\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17146\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__17146\,
            I => \N__17143\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__17143\,
            I => \N__17140\
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__17140\,
            I => \tok.n18_adj_850\
        );

    \I__2436\ : InMux
    port map (
            O => \N__17137\,
            I => \N__17134\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__17134\,
            I => \tok.n17_adj_853\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__17131\,
            I => \tok.n31_cascade_\
        );

    \I__2433\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17125\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__17125\,
            I => \N__17122\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__17122\,
            I => \tok.n299\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__17119\,
            I => \N__17116\
        );

    \I__2429\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17113\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__17113\,
            I => \tok.n6446\
        );

    \I__2427\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17107\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__17107\,
            I => \N__17104\
        );

    \I__2425\ : Odrv12
    port map (
            O => \N__17104\,
            I => \tok.n308\
        );

    \I__2424\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17098\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__17098\,
            I => \N__17095\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__17095\,
            I => \tok.n294\
        );

    \I__2421\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17089\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__17089\,
            I => \tok.n161_adj_667\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__17086\,
            I => \tok.n6371_cascade_\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__17083\,
            I => \N__17080\
        );

    \I__2417\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17077\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__17077\,
            I => \tok.n248_adj_653\
        );

    \I__2415\ : InMux
    port map (
            O => \N__17074\,
            I => \tok.n4795\
        );

    \I__2414\ : InMux
    port map (
            O => \N__17071\,
            I => \bfn_5_10_0_\
        );

    \I__2413\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17065\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__17065\,
            I => \N__17062\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__17062\,
            I => \tok.n293\
        );

    \I__2410\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17056\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__17056\,
            I => \tok.n297\
        );

    \I__2408\ : InMux
    port map (
            O => \N__17053\,
            I => \N__17050\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__17050\,
            I => \tok.n310\
        );

    \I__2406\ : InMux
    port map (
            O => \N__17047\,
            I => \N__17044\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__17044\,
            I => \tok.n6452\
        );

    \I__2404\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17038\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__17038\,
            I => \tok.n2579\
        );

    \I__2402\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17032\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__17032\,
            I => \tok.n6392\
        );

    \I__2400\ : InMux
    port map (
            O => \N__17029\,
            I => \N__17026\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__17026\,
            I => \tok.n6421\
        );

    \I__2398\ : InMux
    port map (
            O => \N__17023\,
            I => \N__17020\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__17020\,
            I => \tok.n300\
        );

    \I__2396\ : InMux
    port map (
            O => \N__17017\,
            I => \tok.n4787\
        );

    \I__2395\ : InMux
    port map (
            O => \N__17014\,
            I => \N__17008\
        );

    \I__2394\ : InMux
    port map (
            O => \N__17013\,
            I => \N__17005\
        );

    \I__2393\ : InMux
    port map (
            O => \N__17012\,
            I => \N__17000\
        );

    \I__2392\ : InMux
    port map (
            O => \N__17011\,
            I => \N__17000\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__17008\,
            I => \N__16997\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__17005\,
            I => \N__16992\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__17000\,
            I => \N__16992\
        );

    \I__2388\ : Span4Mux_v
    port map (
            O => \N__16997\,
            I => \N__16989\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__16992\,
            I => \N__16986\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__16989\,
            I => \tok.n21_adj_660\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__16986\,
            I => \tok.n21_adj_660\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__16981\,
            I => \N__16978\
        );

    \I__2383\ : InMux
    port map (
            O => \N__16978\,
            I => \N__16975\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__16975\,
            I => \N__16972\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__16972\,
            I => \tok.n318\
        );

    \I__2380\ : InMux
    port map (
            O => \N__16969\,
            I => \bfn_5_9_0_\
        );

    \I__2379\ : InMux
    port map (
            O => \N__16966\,
            I => \tok.n4789\
        );

    \I__2378\ : InMux
    port map (
            O => \N__16963\,
            I => \tok.n4790\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__16960\,
            I => \N__16957\
        );

    \I__2376\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16954\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__16954\,
            I => \N__16951\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__16951\,
            I => \tok.n315\
        );

    \I__2373\ : InMux
    port map (
            O => \N__16948\,
            I => \tok.n4791\
        );

    \I__2372\ : InMux
    port map (
            O => \N__16945\,
            I => \tok.n4792\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__16942\,
            I => \N__16939\
        );

    \I__2370\ : InMux
    port map (
            O => \N__16939\,
            I => \N__16936\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__16936\,
            I => \N__16933\
        );

    \I__2368\ : Odrv4
    port map (
            O => \N__16933\,
            I => \tok.n313\
        );

    \I__2367\ : InMux
    port map (
            O => \N__16930\,
            I => \tok.n4793\
        );

    \I__2366\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16923\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__16926\,
            I => \N__16920\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__16923\,
            I => \N__16917\
        );

    \I__2363\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16914\
        );

    \I__2362\ : Span4Mux_s2_h
    port map (
            O => \N__16917\,
            I => \N__16909\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__16914\,
            I => \N__16909\
        );

    \I__2360\ : Span4Mux_h
    port map (
            O => \N__16909\,
            I => \N__16906\
        );

    \I__2359\ : Sp12to4
    port map (
            O => \N__16906\,
            I => \N__16903\
        );

    \I__2358\ : Odrv12
    port map (
            O => \N__16903\,
            I => \tok.n312\
        );

    \I__2357\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16897\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__16897\,
            I => \N__16894\
        );

    \I__2355\ : Span4Mux_h
    port map (
            O => \N__16894\,
            I => \N__16891\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__16891\,
            I => \tok.n295\
        );

    \I__2353\ : InMux
    port map (
            O => \N__16888\,
            I => \tok.n4794\
        );

    \I__2352\ : InMux
    port map (
            O => \N__16885\,
            I => \N__16881\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__16884\,
            I => \N__16878\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__16881\,
            I => \N__16875\
        );

    \I__2349\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16872\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__16875\,
            I => \tok.key_rd_8\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__16872\,
            I => \tok.key_rd_8\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__16867\,
            I => \tok.n20_cascade_\
        );

    \I__2345\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16861\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__16861\,
            I => \N__16858\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__16858\,
            I => \tok.n26_adj_645\
        );

    \I__2342\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16851\
        );

    \I__2341\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16848\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__16851\,
            I => \N__16845\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__16848\,
            I => \tok.key_rd_13\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__16845\,
            I => \tok.key_rd_13\
        );

    \I__2337\ : InMux
    port map (
            O => \N__16840\,
            I => \N__16837\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__16837\,
            I => \tok.n14_adj_644\
        );

    \I__2335\ : InMux
    port map (
            O => \N__16834\,
            I => \bfn_5_8_0_\
        );

    \I__2334\ : InMux
    port map (
            O => \N__16831\,
            I => \tok.n4782\
        );

    \I__2333\ : InMux
    port map (
            O => \N__16828\,
            I => \tok.n4783\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__16825\,
            I => \N__16822\
        );

    \I__2331\ : InMux
    port map (
            O => \N__16822\,
            I => \N__16819\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__16819\,
            I => \tok.n127\
        );

    \I__2329\ : InMux
    port map (
            O => \N__16816\,
            I => \tok.n4784\
        );

    \I__2328\ : InMux
    port map (
            O => \N__16813\,
            I => \N__16810\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__16810\,
            I => \tok.n6557\
        );

    \I__2326\ : InMux
    port map (
            O => \N__16807\,
            I => \tok.n4785\
        );

    \I__2325\ : InMux
    port map (
            O => \N__16804\,
            I => \N__16801\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__16801\,
            I => \tok.n320\
        );

    \I__2323\ : InMux
    port map (
            O => \N__16798\,
            I => \tok.n4786\
        );

    \I__2322\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16789\
        );

    \I__2321\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16789\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__16789\,
            I => \tok.n12\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__16786\,
            I => \N__16783\
        );

    \I__2318\ : InMux
    port map (
            O => \N__16783\,
            I => \N__16776\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__16782\,
            I => \N__16772\
        );

    \I__2316\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16766\
        );

    \I__2315\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16761\
        );

    \I__2314\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16761\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__16776\,
            I => \N__16758\
        );

    \I__2312\ : InMux
    port map (
            O => \N__16775\,
            I => \N__16755\
        );

    \I__2311\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16748\
        );

    \I__2310\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16748\
        );

    \I__2309\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16748\
        );

    \I__2308\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16745\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__16766\,
            I => \N__16740\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__16761\,
            I => \N__16740\
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__16758\,
            I => \tok.n796\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__16755\,
            I => \tok.n796\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__16748\,
            I => \tok.n796\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__16745\,
            I => \tok.n796\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__16740\,
            I => \tok.n796\
        );

    \I__2300\ : InMux
    port map (
            O => \N__16729\,
            I => \N__16720\
        );

    \I__2299\ : InMux
    port map (
            O => \N__16728\,
            I => \N__16720\
        );

    \I__2298\ : InMux
    port map (
            O => \N__16727\,
            I => \N__16720\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__16720\,
            I => \tok.n2702\
        );

    \I__2296\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16711\
        );

    \I__2295\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16704\
        );

    \I__2294\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16704\
        );

    \I__2293\ : InMux
    port map (
            O => \N__16714\,
            I => \N__16704\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__16711\,
            I => \tok.uart_stall\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__16704\,
            I => \tok.uart_stall\
        );

    \I__2290\ : InMux
    port map (
            O => \N__16699\,
            I => \N__16696\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__16696\,
            I => \tok.n6203\
        );

    \I__2288\ : InMux
    port map (
            O => \N__16693\,
            I => \N__16690\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__16690\,
            I => \tok.search_clk_N_137\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__16687\,
            I => \tok.n31_adj_637_cascade_\
        );

    \I__2285\ : InMux
    port map (
            O => \N__16684\,
            I => \N__16681\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__16681\,
            I => \tok.n6170\
        );

    \I__2283\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16672\
        );

    \I__2282\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16672\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__16672\,
            I => \N__16663\
        );

    \I__2280\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16660\
        );

    \I__2279\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16657\
        );

    \I__2278\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16648\
        );

    \I__2277\ : InMux
    port map (
            O => \N__16668\,
            I => \N__16648\
        );

    \I__2276\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16648\
        );

    \I__2275\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16648\
        );

    \I__2274\ : Span12Mux_s5_v
    port map (
            O => \N__16663\,
            I => \N__16643\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__16660\,
            I => \N__16643\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__16657\,
            I => \tok.n30\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__16648\,
            I => \tok.n30\
        );

    \I__2270\ : Odrv12
    port map (
            O => \N__16643\,
            I => \tok.n30\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__16636\,
            I => \tok.n221_adj_753_cascade_\
        );

    \I__2268\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16630\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__16630\,
            I => \N__16626\
        );

    \I__2266\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16623\
        );

    \I__2265\ : Span4Mux_h
    port map (
            O => \N__16626\,
            I => \N__16620\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__16623\,
            I => \tok.key_rd_3\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__16620\,
            I => \tok.key_rd_3\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__16615\,
            I => \N__16612\
        );

    \I__2261\ : InMux
    port map (
            O => \N__16612\,
            I => \N__16609\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__16609\,
            I => \N__16605\
        );

    \I__2259\ : InMux
    port map (
            O => \N__16608\,
            I => \N__16602\
        );

    \I__2258\ : Span4Mux_h
    port map (
            O => \N__16605\,
            I => \N__16599\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__16602\,
            I => \tok.key_rd_5\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__16599\,
            I => \tok.key_rd_5\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__16594\,
            I => \tok.n9_adj_651_cascade_\
        );

    \I__2254\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16588\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__16588\,
            I => \N__16585\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__16585\,
            I => \tok.n13\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__16582\,
            I => \n15_cascade_\
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__16579\,
            I => \tok.n6_adj_687_cascade_\
        );

    \I__2249\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16572\
        );

    \I__2248\ : InMux
    port map (
            O => \N__16575\,
            I => \N__16569\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__16572\,
            I => \N__16565\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__16569\,
            I => \N__16562\
        );

    \I__2245\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16559\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__16565\,
            I => \tok.n4_adj_641\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__16562\,
            I => \tok.n4_adj_641\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__16559\,
            I => \tok.n4_adj_641\
        );

    \I__2241\ : InMux
    port map (
            O => \N__16552\,
            I => \N__16549\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__16549\,
            I => \tok.n5\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__16546\,
            I => \tok.n796_cascade_\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__16543\,
            I => \tok.n80_cascade_\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__16540\,
            I => \tok.n89_cascade_\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__16537\,
            I => \tok.n83_adj_734_cascade_\
        );

    \I__2235\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16531\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__16531\,
            I => \tok.n6279\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__16528\,
            I => \N__16524\
        );

    \I__2232\ : InMux
    port map (
            O => \N__16527\,
            I => \N__16519\
        );

    \I__2231\ : InMux
    port map (
            O => \N__16524\,
            I => \N__16519\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__16519\,
            I => \N__16516\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__16516\,
            I => \N__16513\
        );

    \I__2228\ : Span4Mux_v
    port map (
            O => \N__16513\,
            I => \N__16510\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__16510\,
            I => \tok.table_rd_0\
        );

    \I__2226\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16504\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__16504\,
            I => \N__16501\
        );

    \I__2224\ : Span4Mux_h
    port map (
            O => \N__16501\,
            I => \N__16498\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__16498\,
            I => \N__16495\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__16495\,
            I => \tok.table_wr_data_14\
        );

    \I__2221\ : InMux
    port map (
            O => \N__16492\,
            I => \N__16489\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__16489\,
            I => \N__16486\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__16486\,
            I => \N__16483\
        );

    \I__2218\ : Span4Mux_v
    port map (
            O => \N__16483\,
            I => \N__16480\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__16480\,
            I => \tok.table_wr_data_11\
        );

    \I__2216\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16474\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__16474\,
            I => \N__16471\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__16471\,
            I => \N__16468\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__16468\,
            I => \tok.table_wr_data_12\
        );

    \I__2212\ : InMux
    port map (
            O => \N__16465\,
            I => \N__16462\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__16462\,
            I => \tok.n2696\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__16459\,
            I => \tok.ram.n6266_cascade_\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__16456\,
            I => \tok.n1495_cascade_\
        );

    \I__2208\ : InMux
    port map (
            O => \N__16453\,
            I => \N__16450\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__16450\,
            I => \tok.n13_adj_766\
        );

    \I__2206\ : InMux
    port map (
            O => \N__16447\,
            I => \N__16444\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__16444\,
            I => n10_adj_907
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__16441\,
            I => \n10_adj_907_cascade_\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__16438\,
            I => \N__16435\
        );

    \I__2202\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16432\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__16432\,
            I => \N__16429\
        );

    \I__2200\ : Span4Mux_v
    port map (
            O => \N__16429\,
            I => \N__16426\
        );

    \I__2199\ : Span4Mux_v
    port map (
            O => \N__16426\,
            I => \N__16423\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__16423\,
            I => \tok.tc_6\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__16420\,
            I => \tok.n83_adj_765_cascade_\
        );

    \I__2196\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16414\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__16414\,
            I => \tok.n6435\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__16411\,
            I => \tok.n6283_cascade_\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__16408\,
            I => \N__16405\
        );

    \I__2192\ : InMux
    port map (
            O => \N__16405\,
            I => \N__16399\
        );

    \I__2191\ : InMux
    port map (
            O => \N__16404\,
            I => \N__16399\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__16399\,
            I => \tok.A_stk.tail_7\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__16396\,
            I => \N__16393\
        );

    \I__2188\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16390\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__16390\,
            I => \N__16386\
        );

    \I__2186\ : InMux
    port map (
            O => \N__16389\,
            I => \N__16383\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__16386\,
            I => tail_97
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__16383\,
            I => tail_97
        );

    \I__2183\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16374\
        );

    \I__2182\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16371\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__16374\,
            I => tail_113
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__16371\,
            I => tail_113
        );

    \I__2179\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16362\
        );

    \I__2178\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16359\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__16362\,
            I => tail_108
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__16359\,
            I => tail_108
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__16354\,
            I => \N__16351\
        );

    \I__2174\ : InMux
    port map (
            O => \N__16351\,
            I => \N__16347\
        );

    \I__2173\ : InMux
    port map (
            O => \N__16350\,
            I => \N__16344\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__16347\,
            I => tail_124
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__16344\,
            I => tail_124
        );

    \I__2170\ : InMux
    port map (
            O => \N__16339\,
            I => \N__16336\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__16336\,
            I => \N__16333\
        );

    \I__2168\ : Span4Mux_v
    port map (
            O => \N__16333\,
            I => \N__16330\
        );

    \I__2167\ : Span4Mux_v
    port map (
            O => \N__16330\,
            I => \N__16327\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__16327\,
            I => \tok.table_wr_data_3\
        );

    \I__2165\ : InMux
    port map (
            O => \N__16324\,
            I => \N__16321\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__16321\,
            I => \N__16318\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__16318\,
            I => \N__16315\
        );

    \I__2162\ : Span4Mux_v
    port map (
            O => \N__16315\,
            I => \N__16312\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__16312\,
            I => table_wr_data_1
        );

    \I__2160\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16306\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__16306\,
            I => \N__16303\
        );

    \I__2158\ : Span4Mux_v
    port map (
            O => \N__16303\,
            I => \N__16300\
        );

    \I__2157\ : Span4Mux_v
    port map (
            O => \N__16300\,
            I => \N__16297\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__16297\,
            I => \tok.table_wr_data_6\
        );

    \I__2155\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16291\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__16291\,
            I => \N__16288\
        );

    \I__2153\ : Span12Mux_v
    port map (
            O => \N__16288\,
            I => \N__16285\
        );

    \I__2152\ : Odrv12
    port map (
            O => \N__16285\,
            I => \tok.table_wr_data_4\
        );

    \I__2151\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16279\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__16279\,
            I => \N__16276\
        );

    \I__2149\ : Span4Mux_v
    port map (
            O => \N__16276\,
            I => \N__16273\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__16273\,
            I => \N__16270\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__16270\,
            I => \tok.table_wr_data_2\
        );

    \I__2146\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16264\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__16264\,
            I => \tok.n6412\
        );

    \I__2144\ : InMux
    port map (
            O => \N__16261\,
            I => \N__16257\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__16260\,
            I => \N__16254\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__16257\,
            I => \N__16251\
        );

    \I__2141\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16248\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__16251\,
            I => tail_119
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__16248\,
            I => tail_119
        );

    \I__2138\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16240\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__16240\,
            I => \N__16236\
        );

    \I__2136\ : InMux
    port map (
            O => \N__16239\,
            I => \N__16233\
        );

    \I__2135\ : Odrv12
    port map (
            O => \N__16236\,
            I => tail_103
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__16233\,
            I => tail_103
        );

    \I__2133\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16222\
        );

    \I__2132\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16222\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__16222\,
            I => \tok.A_stk.tail_87\
        );

    \I__2130\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16213\
        );

    \I__2129\ : InMux
    port map (
            O => \N__16218\,
            I => \N__16213\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__16213\,
            I => \tok.A_stk.tail_71\
        );

    \I__2127\ : InMux
    port map (
            O => \N__16210\,
            I => \N__16204\
        );

    \I__2126\ : InMux
    port map (
            O => \N__16209\,
            I => \N__16204\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__16204\,
            I => \tok.A_stk.tail_55\
        );

    \I__2124\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16195\
        );

    \I__2123\ : InMux
    port map (
            O => \N__16200\,
            I => \N__16195\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__16195\,
            I => \tok.A_stk.tail_39\
        );

    \I__2121\ : InMux
    port map (
            O => \N__16192\,
            I => \N__16188\
        );

    \I__2120\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16185\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__16188\,
            I => \tok.A_stk.tail_23\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__16185\,
            I => \tok.A_stk.tail_23\
        );

    \I__2117\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16177\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__16177\,
            I => \N__16174\
        );

    \I__2115\ : Span4Mux_s3_v
    port map (
            O => \N__16174\,
            I => \N__16171\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__16171\,
            I => \tok.table_rd_11\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__16168\,
            I => \tok.n228_cascade_\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__16165\,
            I => \tok.n203_adj_879_cascade_\
        );

    \I__2111\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16159\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__16159\,
            I => \tok.n228\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__16156\,
            I => \tok.n212_adj_880_cascade_\
        );

    \I__2108\ : InMux
    port map (
            O => \N__16153\,
            I => \N__16150\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__16150\,
            I => \N__16147\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__16147\,
            I => \tok.n6339\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__16144\,
            I => \tok.n161_adj_692_cascade_\
        );

    \I__2104\ : InMux
    port map (
            O => \N__16141\,
            I => \N__16138\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__16138\,
            I => \N__16135\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__16135\,
            I => \tok.n6356\
        );

    \I__2101\ : InMux
    port map (
            O => \N__16132\,
            I => \N__16129\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__16129\,
            I => \tok.n6417\
        );

    \I__2099\ : InMux
    port map (
            O => \N__16126\,
            I => \N__16123\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__16123\,
            I => \tok.n206_adj_881\
        );

    \I__2097\ : InMux
    port map (
            O => \N__16120\,
            I => \N__16108\
        );

    \I__2096\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16108\
        );

    \I__2095\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16101\
        );

    \I__2094\ : InMux
    port map (
            O => \N__16117\,
            I => \N__16101\
        );

    \I__2093\ : InMux
    port map (
            O => \N__16116\,
            I => \N__16101\
        );

    \I__2092\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16094\
        );

    \I__2091\ : InMux
    port map (
            O => \N__16114\,
            I => \N__16094\
        );

    \I__2090\ : InMux
    port map (
            O => \N__16113\,
            I => \N__16094\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__16108\,
            I => \tok.n83\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__16101\,
            I => \tok.n83\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__16094\,
            I => \tok.n83\
        );

    \I__2086\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16084\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__16084\,
            I => \N__16081\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__16081\,
            I => \N__16078\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__16078\,
            I => \tok.n161_adj_836\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__16075\,
            I => \tok.n197_adj_837_cascade_\
        );

    \I__2081\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16069\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__16069\,
            I => \N__16066\
        );

    \I__2079\ : Span4Mux_v
    port map (
            O => \N__16066\,
            I => \N__16063\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__16063\,
            I => \tok.n248_adj_838\
        );

    \I__2077\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16057\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__16057\,
            I => \N__16054\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__16054\,
            I => \N__16051\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__16051\,
            I => \tok.n161_adj_650\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__16048\,
            I => \tok.n6386_cascade_\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__16045\,
            I => \tok.n197_adj_652_cascade_\
        );

    \I__2071\ : InMux
    port map (
            O => \N__16042\,
            I => \tok.n4807\
        );

    \I__2070\ : InMux
    port map (
            O => \N__16039\,
            I => \tok.n4808\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__16036\,
            I => \N__16033\
        );

    \I__2068\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16030\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__16030\,
            I => \N__16027\
        );

    \I__2066\ : Odrv12
    port map (
            O => \N__16027\,
            I => \tok.n6377\
        );

    \I__2065\ : InMux
    port map (
            O => \N__16024\,
            I => \tok.n4809\
        );

    \I__2064\ : InMux
    port map (
            O => \N__16021\,
            I => \bfn_4_11_0_\
        );

    \I__2063\ : InMux
    port map (
            O => \N__16018\,
            I => \tok.n4811\
        );

    \I__2062\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16012\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__16012\,
            I => \tok.n6362\
        );

    \I__2060\ : InMux
    port map (
            O => \N__16009\,
            I => \tok.n4799\
        );

    \I__2059\ : InMux
    port map (
            O => \N__16006\,
            I => \N__16003\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__16003\,
            I => \tok.n6556\
        );

    \I__2057\ : InMux
    port map (
            O => \N__16000\,
            I => \tok.n4800\
        );

    \I__2056\ : InMux
    port map (
            O => \N__15997\,
            I => \tok.n4801\
        );

    \I__2055\ : InMux
    port map (
            O => \N__15994\,
            I => \tok.n4802\
        );

    \I__2054\ : InMux
    port map (
            O => \N__15991\,
            I => \bfn_4_10_0_\
        );

    \I__2053\ : InMux
    port map (
            O => \N__15988\,
            I => \tok.n4804\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__15985\,
            I => \N__15982\
        );

    \I__2051\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15979\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__15979\,
            I => \N__15976\
        );

    \I__2049\ : Odrv12
    port map (
            O => \N__15976\,
            I => \tok.n6437\
        );

    \I__2048\ : InMux
    port map (
            O => \N__15973\,
            I => \tok.n4805\
        );

    \I__2047\ : InMux
    port map (
            O => \N__15970\,
            I => \tok.n4806\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__15967\,
            I => \N__15964\
        );

    \I__2045\ : InMux
    port map (
            O => \N__15964\,
            I => \N__15958\
        );

    \I__2044\ : InMux
    port map (
            O => \N__15963\,
            I => \N__15958\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__15958\,
            I => \tok.key_rd_6\
        );

    \I__2042\ : InMux
    port map (
            O => \N__15955\,
            I => \N__15949\
        );

    \I__2041\ : InMux
    port map (
            O => \N__15954\,
            I => \N__15949\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__15949\,
            I => \tok.key_rd_0\
        );

    \I__2039\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15943\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__15943\,
            I => \N__15940\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__15940\,
            I => \tok.n25\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__15937\,
            I => \N__15934\
        );

    \I__2035\ : InMux
    port map (
            O => \N__15934\,
            I => \N__15928\
        );

    \I__2034\ : InMux
    port map (
            O => \N__15933\,
            I => \N__15928\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__15928\,
            I => \tok.key_rd_4\
        );

    \I__2032\ : InMux
    port map (
            O => \N__15925\,
            I => \N__15919\
        );

    \I__2031\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15919\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__15919\,
            I => \tok.key_rd_1\
        );

    \I__2029\ : InMux
    port map (
            O => \N__15916\,
            I => \N__15913\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__15913\,
            I => \N__15910\
        );

    \I__2027\ : Span4Mux_h
    port map (
            O => \N__15910\,
            I => \N__15907\
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__15907\,
            I => \tok.n18\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__15904\,
            I => \tok.n6575_cascade_\
        );

    \I__2024\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15898\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__15898\,
            I => \tok.n177\
        );

    \I__2022\ : InMux
    port map (
            O => \N__15895\,
            I => \tok.n4797\
        );

    \I__2021\ : InMux
    port map (
            O => \N__15892\,
            I => \tok.n4798\
        );

    \I__2020\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15886\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__15886\,
            I => \N__15883\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__15883\,
            I => \tok.n33\
        );

    \I__2017\ : InMux
    port map (
            O => \N__15880\,
            I => \N__15877\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__15877\,
            I => \tok.n27_adj_707\
        );

    \I__2015\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15871\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__15871\,
            I => \N__15868\
        );

    \I__2013\ : Odrv12
    port map (
            O => \N__15868\,
            I => \tok.n33_adj_663\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__15865\,
            I => \tok.n27_adj_708_cascade_\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__15862\,
            I => \N__15858\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__15861\,
            I => \N__15855\
        );

    \I__2009\ : CascadeBuf
    port map (
            O => \N__15858\,
            I => \N__15852\
        );

    \I__2008\ : CascadeBuf
    port map (
            O => \N__15855\,
            I => \N__15849\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__15852\,
            I => \N__15846\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__15849\,
            I => \N__15841\
        );

    \I__2005\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15837\
        );

    \I__2004\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15834\
        );

    \I__2003\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15831\
        );

    \I__2002\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15828\
        );

    \I__2001\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15825\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__15837\,
            I => \N__15822\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__15834\,
            I => \N__15817\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__15831\,
            I => \N__15817\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__15828\,
            I => \N__15814\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__15825\,
            I => \N__15809\
        );

    \I__1995\ : Span4Mux_h
    port map (
            O => \N__15822\,
            I => \N__15809\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__15817\,
            I => \tok.n29\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__15814\,
            I => \tok.n29\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__15809\,
            I => \tok.n29\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__15802\,
            I => \N__15798\
        );

    \I__1990\ : InMux
    port map (
            O => \N__15801\,
            I => \N__15789\
        );

    \I__1989\ : InMux
    port map (
            O => \N__15798\,
            I => \N__15789\
        );

    \I__1988\ : InMux
    port map (
            O => \N__15797\,
            I => \N__15789\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__15796\,
            I => \N__15784\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__15789\,
            I => \N__15780\
        );

    \I__1985\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15773\
        );

    \I__1984\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15773\
        );

    \I__1983\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15773\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__15783\,
            I => \N__15768\
        );

    \I__1981\ : Span4Mux_h
    port map (
            O => \N__15780\,
            I => \N__15763\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__15773\,
            I => \N__15760\
        );

    \I__1979\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15749\
        );

    \I__1978\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15749\
        );

    \I__1977\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15749\
        );

    \I__1976\ : InMux
    port map (
            O => \N__15767\,
            I => \N__15749\
        );

    \I__1975\ : InMux
    port map (
            O => \N__15766\,
            I => \N__15749\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__15763\,
            I => \tok.search_clk\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__15760\,
            I => \tok.search_clk\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__15749\,
            I => \tok.search_clk\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__15742\,
            I => \N__15736\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__15741\,
            I => \N__15733\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__15740\,
            I => \N__15730\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__15739\,
            I => \N__15727\
        );

    \I__1967\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15714\
        );

    \I__1966\ : InMux
    port map (
            O => \N__15733\,
            I => \N__15714\
        );

    \I__1965\ : InMux
    port map (
            O => \N__15730\,
            I => \N__15714\
        );

    \I__1964\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15714\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__15726\,
            I => \N__15710\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__15725\,
            I => \N__15707\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__15724\,
            I => \N__15704\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__15723\,
            I => \N__15701\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__15714\,
            I => \N__15698\
        );

    \I__1958\ : InMux
    port map (
            O => \N__15713\,
            I => \N__15695\
        );

    \I__1957\ : InMux
    port map (
            O => \N__15710\,
            I => \N__15686\
        );

    \I__1956\ : InMux
    port map (
            O => \N__15707\,
            I => \N__15686\
        );

    \I__1955\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15686\
        );

    \I__1954\ : InMux
    port map (
            O => \N__15701\,
            I => \N__15686\
        );

    \I__1953\ : Span4Mux_s2_h
    port map (
            O => \N__15698\,
            I => \N__15681\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__15695\,
            I => \N__15681\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__15686\,
            I => \tok.found_slot\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__15681\,
            I => \tok.found_slot\
        );

    \I__1949\ : InMux
    port map (
            O => \N__15676\,
            I => \N__15673\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__15673\,
            I => \N__15670\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__15670\,
            I => \N__15667\
        );

    \I__1946\ : Span4Mux_s2_h
    port map (
            O => \N__15667\,
            I => \N__15664\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__15664\,
            I => \tok.n6670\
        );

    \I__1944\ : InMux
    port map (
            O => \N__15661\,
            I => \N__15658\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__15658\,
            I => \N__15655\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__15655\,
            I => \N__15652\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__15652\,
            I => \tok.n33_adj_633\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__15649\,
            I => \tok.n27_adj_704_cascade_\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__15646\,
            I => \N__15642\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__15645\,
            I => \N__15639\
        );

    \I__1937\ : CascadeBuf
    port map (
            O => \N__15642\,
            I => \N__15636\
        );

    \I__1936\ : CascadeBuf
    port map (
            O => \N__15639\,
            I => \N__15633\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__15636\,
            I => \N__15628\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__15633\,
            I => \N__15625\
        );

    \I__1933\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15622\
        );

    \I__1932\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15619\
        );

    \I__1931\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15616\
        );

    \I__1930\ : InMux
    port map (
            O => \N__15625\,
            I => \N__15613\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__15622\,
            I => \N__15608\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__15619\,
            I => \N__15608\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__15616\,
            I => \N__15603\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__15613\,
            I => \N__15603\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__15608\,
            I => \N__15599\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__15603\,
            I => \N__15596\
        );

    \I__1923\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15593\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__15599\,
            I => \N__15590\
        );

    \I__1921\ : Span4Mux_s3_h
    port map (
            O => \N__15596\,
            I => \N__15587\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__15593\,
            I => \tok.n38\
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__15590\,
            I => \tok.n38\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__15587\,
            I => \tok.n38\
        );

    \I__1917\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15577\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__15577\,
            I => \N__15574\
        );

    \I__1915\ : Span4Mux_v
    port map (
            O => \N__15574\,
            I => \N__15571\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__15571\,
            I => \tok.n33_adj_632\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__15568\,
            I => \N__15565\
        );

    \I__1912\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15562\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__15562\,
            I => \N__15559\
        );

    \I__1910\ : Span4Mux_h
    port map (
            O => \N__15559\,
            I => \N__15556\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__15556\,
            I => \tok.n33_adj_661\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__15553\,
            I => \tok.n27_adj_705_cascade_\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__15550\,
            I => \N__15546\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__15549\,
            I => \N__15543\
        );

    \I__1905\ : CascadeBuf
    port map (
            O => \N__15546\,
            I => \N__15539\
        );

    \I__1904\ : CascadeBuf
    port map (
            O => \N__15543\,
            I => \N__15536\
        );

    \I__1903\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15533\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__15539\,
            I => \N__15529\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__15536\,
            I => \N__15526\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__15533\,
            I => \N__15523\
        );

    \I__1899\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15520\
        );

    \I__1898\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15517\
        );

    \I__1897\ : InMux
    port map (
            O => \N__15526\,
            I => \N__15514\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__15523\,
            I => \N__15510\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__15520\,
            I => \N__15507\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__15517\,
            I => \N__15502\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__15514\,
            I => \N__15502\
        );

    \I__1892\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15499\
        );

    \I__1891\ : Span4Mux_s1_h
    port map (
            O => \N__15510\,
            I => \N__15494\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__15507\,
            I => \N__15494\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__15502\,
            I => \N__15491\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__15499\,
            I => \tok.n36\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__15494\,
            I => \tok.n36\
        );

    \I__1886\ : Odrv4
    port map (
            O => \N__15491\,
            I => \tok.n36\
        );

    \I__1885\ : InMux
    port map (
            O => \N__15484\,
            I => \N__15481\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__15481\,
            I => \tok.n27_adj_703\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__15478\,
            I => \N__15474\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__15477\,
            I => \N__15471\
        );

    \I__1881\ : CascadeBuf
    port map (
            O => \N__15474\,
            I => \N__15468\
        );

    \I__1880\ : CascadeBuf
    port map (
            O => \N__15471\,
            I => \N__15465\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__15468\,
            I => \N__15462\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__15465\,
            I => \N__15457\
        );

    \I__1877\ : InMux
    port map (
            O => \N__15462\,
            I => \N__15454\
        );

    \I__1876\ : InMux
    port map (
            O => \N__15461\,
            I => \N__15451\
        );

    \I__1875\ : InMux
    port map (
            O => \N__15460\,
            I => \N__15448\
        );

    \I__1874\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15445\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__15454\,
            I => \N__15442\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__15451\,
            I => \N__15436\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__15448\,
            I => \N__15436\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__15445\,
            I => \N__15433\
        );

    \I__1869\ : Span4Mux_h
    port map (
            O => \N__15442\,
            I => \N__15430\
        );

    \I__1868\ : InMux
    port map (
            O => \N__15441\,
            I => \N__15427\
        );

    \I__1867\ : Span4Mux_h
    port map (
            O => \N__15436\,
            I => \N__15424\
        );

    \I__1866\ : Span4Mux_v
    port map (
            O => \N__15433\,
            I => \N__15419\
        );

    \I__1865\ : Span4Mux_v
    port map (
            O => \N__15430\,
            I => \N__15419\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__15427\,
            I => \tok.n40\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__15424\,
            I => \tok.n40\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__15419\,
            I => \tok.n40\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__15412\,
            I => \N__15408\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__15411\,
            I => \N__15405\
        );

    \I__1859\ : CascadeBuf
    port map (
            O => \N__15408\,
            I => \N__15402\
        );

    \I__1858\ : CascadeBuf
    port map (
            O => \N__15405\,
            I => \N__15399\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__15402\,
            I => \N__15394\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__15399\,
            I => \N__15391\
        );

    \I__1855\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15388\
        );

    \I__1854\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15385\
        );

    \I__1853\ : InMux
    port map (
            O => \N__15394\,
            I => \N__15382\
        );

    \I__1852\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15379\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__15388\,
            I => \N__15373\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__15385\,
            I => \N__15373\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__15382\,
            I => \N__15368\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__15379\,
            I => \N__15368\
        );

    \I__1847\ : InMux
    port map (
            O => \N__15378\,
            I => \N__15365\
        );

    \I__1846\ : Span12Mux_s8_v
    port map (
            O => \N__15373\,
            I => \N__15362\
        );

    \I__1845\ : Sp12to4
    port map (
            O => \N__15368\,
            I => \N__15359\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__15365\,
            I => \tok.n32\
        );

    \I__1843\ : Odrv12
    port map (
            O => \N__15362\,
            I => \tok.n32\
        );

    \I__1842\ : Odrv12
    port map (
            O => \N__15359\,
            I => \tok.n32\
        );

    \I__1841\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15346\
        );

    \I__1840\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15346\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__15346\,
            I => \tok.A_stk.tail_19\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__15343\,
            I => \N__15340\
        );

    \I__1837\ : InMux
    port map (
            O => \N__15340\,
            I => \N__15334\
        );

    \I__1836\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15334\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__15334\,
            I => \tok.A_stk.tail_3\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__15331\,
            I => \tok.n4_cascade_\
        );

    \I__1833\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15325\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__15325\,
            I => \N__15322\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__15322\,
            I => \tok.n6273\
        );

    \I__1830\ : InMux
    port map (
            O => \N__15319\,
            I => \N__15316\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__15316\,
            I => \N__15313\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__15313\,
            I => \N__15310\
        );

    \I__1827\ : Odrv4
    port map (
            O => \N__15310\,
            I => \tok.table_wr_data_9\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__15307\,
            I => \N__15304\
        );

    \I__1825\ : InMux
    port map (
            O => \N__15304\,
            I => \N__15301\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__15301\,
            I => \tok.n4\
        );

    \I__1823\ : InMux
    port map (
            O => \N__15298\,
            I => \N__15295\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__15295\,
            I => \N__15292\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__15292\,
            I => \tok.n6252\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__15289\,
            I => \tok.n6253_cascade_\
        );

    \I__1819\ : InMux
    port map (
            O => \N__15286\,
            I => \N__15282\
        );

    \I__1818\ : InMux
    port map (
            O => \N__15285\,
            I => \N__15279\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__15282\,
            I => tail_99
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__15279\,
            I => tail_99
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__15274\,
            I => \N__15270\
        );

    \I__1814\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15267\
        );

    \I__1813\ : InMux
    port map (
            O => \N__15270\,
            I => \N__15264\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__15267\,
            I => tail_115
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__15264\,
            I => tail_115
        );

    \I__1810\ : InMux
    port map (
            O => \N__15259\,
            I => \N__15255\
        );

    \I__1809\ : InMux
    port map (
            O => \N__15258\,
            I => \N__15252\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__15255\,
            I => \tok.A_stk.tail_92\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__15252\,
            I => \tok.A_stk.tail_92\
        );

    \I__1806\ : InMux
    port map (
            O => \N__15247\,
            I => \N__15241\
        );

    \I__1805\ : InMux
    port map (
            O => \N__15246\,
            I => \N__15241\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__15241\,
            I => \tok.A_stk.tail_60\
        );

    \I__1803\ : InMux
    port map (
            O => \N__15238\,
            I => \N__15234\
        );

    \I__1802\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15231\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__15234\,
            I => \tok.A_stk.tail_76\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__15231\,
            I => \tok.A_stk.tail_76\
        );

    \I__1799\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15222\
        );

    \I__1798\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15219\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__15222\,
            I => \tok.A_stk.tail_6\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__15219\,
            I => \tok.A_stk.tail_6\
        );

    \I__1795\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15210\
        );

    \I__1794\ : InMux
    port map (
            O => \N__15213\,
            I => \N__15207\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__15210\,
            I => \tok.A_stk.tail_12\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__15207\,
            I => \tok.A_stk.tail_12\
        );

    \I__1791\ : InMux
    port map (
            O => \N__15202\,
            I => \N__15198\
        );

    \I__1790\ : InMux
    port map (
            O => \N__15201\,
            I => \N__15195\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__15198\,
            I => \N__15192\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__15195\,
            I => \N__15189\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__15192\,
            I => \N__15184\
        );

    \I__1786\ : Span4Mux_h
    port map (
            O => \N__15189\,
            I => \N__15184\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__15184\,
            I => \tok.A_stk.tail_10\
        );

    \I__1784\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15175\
        );

    \I__1783\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15175\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__15175\,
            I => \tok.A_stk.tail_83\
        );

    \I__1781\ : InMux
    port map (
            O => \N__15172\,
            I => \N__15166\
        );

    \I__1780\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15166\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__15166\,
            I => \tok.A_stk.tail_67\
        );

    \I__1778\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15157\
        );

    \I__1777\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15157\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__15157\,
            I => \tok.A_stk.tail_51\
        );

    \I__1775\ : InMux
    port map (
            O => \N__15154\,
            I => \N__15148\
        );

    \I__1774\ : InMux
    port map (
            O => \N__15153\,
            I => \N__15148\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__15148\,
            I => \tok.A_stk.tail_35\
        );

    \I__1772\ : InMux
    port map (
            O => \N__15145\,
            I => \N__15139\
        );

    \I__1771\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15139\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__15139\,
            I => \tok.A_stk.tail_70\
        );

    \I__1769\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15130\
        );

    \I__1768\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15130\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__15130\,
            I => \tok.A_stk.tail_54\
        );

    \I__1766\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15121\
        );

    \I__1765\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15121\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__15121\,
            I => \tok.A_stk.tail_38\
        );

    \I__1763\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15114\
        );

    \I__1762\ : InMux
    port map (
            O => \N__15117\,
            I => \N__15111\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__15114\,
            I => \tok.A_stk.tail_22\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__15111\,
            I => \tok.A_stk.tail_22\
        );

    \I__1759\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15100\
        );

    \I__1758\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15100\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__15100\,
            I => \tok.A_stk.tail_28\
        );

    \I__1756\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15091\
        );

    \I__1755\ : InMux
    port map (
            O => \N__15096\,
            I => \N__15091\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__15091\,
            I => \tok.A_stk.tail_44\
        );

    \I__1753\ : InMux
    port map (
            O => \N__15088\,
            I => \N__15082\
        );

    \I__1752\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15082\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__15082\,
            I => \tok.A_stk.tail_65\
        );

    \I__1750\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15073\
        );

    \I__1749\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15073\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__15073\,
            I => tail_49
        );

    \I__1747\ : InMux
    port map (
            O => \N__15070\,
            I => \N__15064\
        );

    \I__1746\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15064\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__15064\,
            I => tail_81
        );

    \I__1744\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15055\
        );

    \I__1743\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15055\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__15055\,
            I => \tok.A_stk.tail_33\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__15052\,
            I => \N__15049\
        );

    \I__1740\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15043\
        );

    \I__1739\ : InMux
    port map (
            O => \N__15048\,
            I => \N__15043\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__15043\,
            I => tail_17
        );

    \I__1737\ : InMux
    port map (
            O => \N__15040\,
            I => \N__15034\
        );

    \I__1736\ : InMux
    port map (
            O => \N__15039\,
            I => \N__15034\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__15034\,
            I => \tok.A_stk.tail_1\
        );

    \I__1734\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15027\
        );

    \I__1733\ : InMux
    port map (
            O => \N__15030\,
            I => \N__15024\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__15027\,
            I => \N__15021\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__15024\,
            I => tail_102
        );

    \I__1730\ : Odrv12
    port map (
            O => \N__15021\,
            I => tail_102
        );

    \I__1729\ : InMux
    port map (
            O => \N__15016\,
            I => \N__15012\
        );

    \I__1728\ : InMux
    port map (
            O => \N__15015\,
            I => \N__15009\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__15012\,
            I => \N__15006\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__15009\,
            I => \tok.A_stk.tail_86\
        );

    \I__1725\ : Odrv12
    port map (
            O => \N__15006\,
            I => \tok.A_stk.tail_86\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__15001\,
            I => \tok.n281_cascade_\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__14998\,
            I => \tok.n236_adj_864_cascade_\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__14995\,
            I => \tok.n2648_cascade_\
        );

    \I__1721\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14989\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__14989\,
            I => \tok.n226_adj_865\
        );

    \I__1719\ : InMux
    port map (
            O => \N__14986\,
            I => \N__14983\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__14983\,
            I => \tok.n6334\
        );

    \I__1717\ : InMux
    port map (
            O => \N__14980\,
            I => \N__14977\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__14977\,
            I => \tok.n4_adj_762\
        );

    \I__1715\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14971\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__14971\,
            I => \tok.n6316\
        );

    \I__1713\ : InMux
    port map (
            O => \N__14968\,
            I => \N__14965\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__14965\,
            I => \N__14961\
        );

    \I__1711\ : InMux
    port map (
            O => \N__14964\,
            I => \N__14958\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__14961\,
            I => sender_1
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__14958\,
            I => sender_1
        );

    \I__1708\ : IoInMux
    port map (
            O => \N__14953\,
            I => \N__14950\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__14950\,
            I => \N__14947\
        );

    \I__1706\ : Span4Mux_s0_v
    port map (
            O => \N__14947\,
            I => \N__14944\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__14944\,
            I => tx_c
        );

    \I__1704\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14938\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__14938\,
            I => \N__14935\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__14935\,
            I => \N__14932\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__14932\,
            I => \tok.table_rd_14\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__14929\,
            I => \tok.n225_cascade_\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__14926\,
            I => \tok.n203_adj_664_cascade_\
        );

    \I__1698\ : InMux
    port map (
            O => \N__14923\,
            I => \N__14920\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__14920\,
            I => \tok.n225\
        );

    \I__1696\ : InMux
    port map (
            O => \N__14917\,
            I => \N__14914\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__14914\,
            I => \tok.n224\
        );

    \I__1694\ : InMux
    port map (
            O => \N__14911\,
            I => \N__14908\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__14908\,
            I => \N__14905\
        );

    \I__1692\ : Span4Mux_s3_v
    port map (
            O => \N__14905\,
            I => \N__14902\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__14902\,
            I => \tok.table_rd_15\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__14899\,
            I => \tok.n224_cascade_\
        );

    \I__1689\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14893\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__14893\,
            I => \tok.n203_adj_688\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__14890\,
            I => \tok.n6373_cascade_\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__14887\,
            I => \tok.n206_adj_666_cascade_\
        );

    \I__1685\ : InMux
    port map (
            O => \N__14884\,
            I => \N__14881\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__14881\,
            I => \tok.n212_adj_665\
        );

    \I__1683\ : InMux
    port map (
            O => \N__14878\,
            I => \tok.n4779\
        );

    \I__1682\ : InMux
    port map (
            O => \N__14875\,
            I => \tok.n4780\
        );

    \I__1681\ : InMux
    port map (
            O => \N__14872\,
            I => \bfn_2_11_0_\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__14869\,
            I => \tok.n214_cascade_\
        );

    \I__1679\ : InMux
    port map (
            O => \N__14866\,
            I => \N__14863\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__14863\,
            I => \N__14860\
        );

    \I__1677\ : Span4Mux_v
    port map (
            O => \N__14860\,
            I => \N__14857\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__14857\,
            I => \tok.n6358\
        );

    \I__1675\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14851\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__14851\,
            I => \N__14848\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__14848\,
            I => \tok.n6402\
        );

    \I__1672\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14842\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__14842\,
            I => \N__14839\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__14839\,
            I => \tok.table_rd_12\
        );

    \I__1669\ : InMux
    port map (
            O => \N__14836\,
            I => \N__14830\
        );

    \I__1668\ : InMux
    port map (
            O => \N__14835\,
            I => \N__14830\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__14830\,
            I => \tok.n227\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__14827\,
            I => \tok.n203_cascade_\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__14824\,
            I => \tok.n212_cascade_\
        );

    \I__1664\ : InMux
    port map (
            O => \N__14821\,
            I => \N__14818\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__14818\,
            I => \tok.n206\
        );

    \I__1662\ : InMux
    port map (
            O => \N__14815\,
            I => \tok.n4774\
        );

    \I__1661\ : InMux
    port map (
            O => \N__14812\,
            I => \tok.n4775\
        );

    \I__1660\ : InMux
    port map (
            O => \N__14809\,
            I => \tok.n4776\
        );

    \I__1659\ : InMux
    port map (
            O => \N__14806\,
            I => \tok.n4777\
        );

    \I__1658\ : InMux
    port map (
            O => \N__14803\,
            I => \tok.n4778\
        );

    \I__1657\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14794\
        );

    \I__1656\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14794\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__14794\,
            I => \tok.key_rd_10\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__14791\,
            I => \N__14787\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__14790\,
            I => \N__14784\
        );

    \I__1652\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14779\
        );

    \I__1651\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14779\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__14779\,
            I => \tok.key_rd_12\
        );

    \I__1649\ : InMux
    port map (
            O => \N__14776\,
            I => \N__14773\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__14773\,
            I => \tok.n26\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__14770\,
            I => \tok.n27_adj_639_cascade_\
        );

    \I__1646\ : InMux
    port map (
            O => \N__14767\,
            I => \N__14764\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__14764\,
            I => \tok.found_slot_N_144\
        );

    \I__1644\ : InMux
    port map (
            O => \N__14761\,
            I => \N__14758\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__14758\,
            I => \tok.n6322\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__14755\,
            I => \tok.n313_cascade_\
        );

    \I__1641\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14748\
        );

    \I__1640\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14745\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__14748\,
            I => \tok.key_rd_2\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__14745\,
            I => \tok.key_rd_2\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__14740\,
            I => \N__14736\
        );

    \I__1636\ : InMux
    port map (
            O => \N__14739\,
            I => \N__14733\
        );

    \I__1635\ : InMux
    port map (
            O => \N__14736\,
            I => \N__14730\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__14733\,
            I => \tok.key_rd_7\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__14730\,
            I => \tok.key_rd_7\
        );

    \I__1632\ : InMux
    port map (
            O => \N__14725\,
            I => \N__14722\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__14722\,
            I => \tok.n22\
        );

    \I__1630\ : InMux
    port map (
            O => \N__14719\,
            I => \N__14716\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__14716\,
            I => \tok.n33_adj_634\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__14713\,
            I => \tok.n27_adj_706_cascade_\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__14710\,
            I => \N__14706\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__14709\,
            I => \N__14703\
        );

    \I__1625\ : CascadeBuf
    port map (
            O => \N__14706\,
            I => \N__14700\
        );

    \I__1624\ : CascadeBuf
    port map (
            O => \N__14703\,
            I => \N__14697\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__14700\,
            I => \N__14694\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__14697\,
            I => \N__14691\
        );

    \I__1621\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14688\
        );

    \I__1620\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14685\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__14688\,
            I => \N__14677\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__14685\,
            I => \N__14677\
        );

    \I__1617\ : InMux
    port map (
            O => \N__14684\,
            I => \N__14674\
        );

    \I__1616\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14671\
        );

    \I__1615\ : InMux
    port map (
            O => \N__14682\,
            I => \N__14668\
        );

    \I__1614\ : Span12Mux_s8_v
    port map (
            O => \N__14677\,
            I => \N__14665\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__14674\,
            I => \tok.n35\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__14671\,
            I => \tok.n35\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__14668\,
            I => \tok.n35\
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__14665\,
            I => \tok.n35\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__14656\,
            I => \tok.n6667_cascade_\
        );

    \I__1608\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14650\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__14650\,
            I => \N__14647\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__14647\,
            I => \tok.n2532\
        );

    \I__1605\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14641\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__14641\,
            I => \N__14638\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__14638\,
            I => \tok.n4_adj_642\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__14635\,
            I => \tok.found_slot_cascade_\
        );

    \I__1601\ : SRMux
    port map (
            O => \N__14632\,
            I => \N__14628\
        );

    \I__1600\ : SRMux
    port map (
            O => \N__14631\,
            I => \N__14625\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__14628\,
            I => \N__14622\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__14625\,
            I => \N__14619\
        );

    \I__1597\ : Span4Mux_h
    port map (
            O => \N__14622\,
            I => \N__14616\
        );

    \I__1596\ : Span4Mux_h
    port map (
            O => \N__14619\,
            I => \N__14613\
        );

    \I__1595\ : Span4Mux_s2_h
    port map (
            O => \N__14616\,
            I => \N__14610\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__14613\,
            I => \tok.write_slot\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__14610\,
            I => \tok.write_slot\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__14605\,
            I => \tok.n21_cascade_\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__14602\,
            I => \N__14599\
        );

    \I__1590\ : InMux
    port map (
            O => \N__14599\,
            I => \N__14596\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__14596\,
            I => \tok.n30_adj_647\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__14593\,
            I => \tok.n4_adj_642_cascade_\
        );

    \I__1587\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14587\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__14587\,
            I => \N__14584\
        );

    \I__1585\ : Span4Mux_v
    port map (
            O => \N__14584\,
            I => \N__14581\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__14581\,
            I => \tok.table_wr_data_13\
        );

    \I__1583\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14575\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__14575\,
            I => \N__14572\
        );

    \I__1581\ : Span4Mux_h
    port map (
            O => \N__14572\,
            I => \N__14569\
        );

    \I__1580\ : Span4Mux_v
    port map (
            O => \N__14569\,
            I => \N__14566\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__14566\,
            I => \tok.table_wr_data_10\
        );

    \I__1578\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14560\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__14560\,
            I => \N__14557\
        );

    \I__1576\ : Span4Mux_v
    port map (
            O => \N__14557\,
            I => \N__14554\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__14554\,
            I => \tok.table_wr_data_15\
        );

    \I__1574\ : InMux
    port map (
            O => \N__14551\,
            I => \N__14548\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__14548\,
            I => \tok.n33_adj_631\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__14545\,
            I => \tok.n27_cascade_\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__14542\,
            I => \N__14538\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__14541\,
            I => \N__14535\
        );

    \I__1569\ : CascadeBuf
    port map (
            O => \N__14538\,
            I => \N__14532\
        );

    \I__1568\ : CascadeBuf
    port map (
            O => \N__14535\,
            I => \N__14529\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__14532\,
            I => \N__14526\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__14529\,
            I => \N__14523\
        );

    \I__1565\ : InMux
    port map (
            O => \N__14526\,
            I => \N__14520\
        );

    \I__1564\ : InMux
    port map (
            O => \N__14523\,
            I => \N__14517\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__14520\,
            I => \N__14509\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__14517\,
            I => \N__14509\
        );

    \I__1561\ : InMux
    port map (
            O => \N__14516\,
            I => \N__14506\
        );

    \I__1560\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14503\
        );

    \I__1559\ : InMux
    port map (
            O => \N__14514\,
            I => \N__14500\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__14509\,
            I => \N__14497\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__14506\,
            I => \tok.n41\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__14503\,
            I => \tok.n41\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__14500\,
            I => \tok.n41\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__14497\,
            I => \tok.n41\
        );

    \I__1553\ : InMux
    port map (
            O => \N__14488\,
            I => \N__14485\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__14485\,
            I => \tok.n33_adj_662\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__14482\,
            I => \tok.n27_adj_709_cascade_\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__14479\,
            I => \N__14475\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__14478\,
            I => \N__14472\
        );

    \I__1548\ : CascadeBuf
    port map (
            O => \N__14475\,
            I => \N__14469\
        );

    \I__1547\ : CascadeBuf
    port map (
            O => \N__14472\,
            I => \N__14466\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__14469\,
            I => \N__14463\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__14466\,
            I => \N__14460\
        );

    \I__1544\ : InMux
    port map (
            O => \N__14463\,
            I => \N__14457\
        );

    \I__1543\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14454\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__14457\,
            I => \N__14446\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__14454\,
            I => \N__14446\
        );

    \I__1540\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14443\
        );

    \I__1539\ : InMux
    port map (
            O => \N__14452\,
            I => \N__14440\
        );

    \I__1538\ : InMux
    port map (
            O => \N__14451\,
            I => \N__14437\
        );

    \I__1537\ : Span4Mux_v
    port map (
            O => \N__14446\,
            I => \N__14434\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__14443\,
            I => \tok.n19\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__14440\,
            I => \tok.n19\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__14437\,
            I => \tok.n19\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__14434\,
            I => \tok.n19\
        );

    \I__1532\ : InMux
    port map (
            O => \N__14425\,
            I => \N__14419\
        );

    \I__1531\ : InMux
    port map (
            O => \N__14424\,
            I => \N__14419\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__14419\,
            I => \tok.A_stk.tail_34\
        );

    \I__1529\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14410\
        );

    \I__1528\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14410\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__14410\,
            I => \tok.A_stk.tail_50\
        );

    \I__1526\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14401\
        );

    \I__1525\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14401\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__14401\,
            I => \tok.A_stk.tail_66\
        );

    \I__1523\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14392\
        );

    \I__1522\ : InMux
    port map (
            O => \N__14397\,
            I => \N__14392\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__14392\,
            I => \tok.A_stk.tail_82\
        );

    \I__1520\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14386\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__14386\,
            I => \N__14383\
        );

    \I__1518\ : Span4Mux_v
    port map (
            O => \N__14383\,
            I => \N__14380\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__14380\,
            I => table_wr_data_0
        );

    \I__1516\ : InMux
    port map (
            O => \N__14377\,
            I => \N__14373\
        );

    \I__1515\ : InMux
    port map (
            O => \N__14376\,
            I => \N__14370\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__14373\,
            I => tail_98
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__14370\,
            I => tail_98
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__14365\,
            I => \N__14361\
        );

    \I__1511\ : InMux
    port map (
            O => \N__14364\,
            I => \N__14358\
        );

    \I__1510\ : InMux
    port map (
            O => \N__14361\,
            I => \N__14355\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__14358\,
            I => tail_114
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__14355\,
            I => tail_114
        );

    \I__1507\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14347\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__14347\,
            I => \N__14343\
        );

    \I__1505\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14340\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__14343\,
            I => \tok.A_stk.tail_26\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__14340\,
            I => \tok.A_stk.tail_26\
        );

    \I__1502\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14332\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__14332\,
            I => \N__14328\
        );

    \I__1500\ : InMux
    port map (
            O => \N__14331\,
            I => \N__14325\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__14328\,
            I => tail_126
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__14325\,
            I => tail_126
        );

    \I__1497\ : InMux
    port map (
            O => \N__14320\,
            I => \N__14317\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__14317\,
            I => \N__14314\
        );

    \I__1495\ : Span4Mux_s2_h
    port map (
            O => \N__14314\,
            I => \N__14310\
        );

    \I__1494\ : InMux
    port map (
            O => \N__14313\,
            I => \N__14307\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__14310\,
            I => tail_110
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__14307\,
            I => tail_110
        );

    \I__1491\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14298\
        );

    \I__1490\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14295\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__14298\,
            I => \tok.A_stk.tail_94\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__14295\,
            I => \tok.A_stk.tail_94\
        );

    \I__1487\ : InMux
    port map (
            O => \N__14290\,
            I => \N__14284\
        );

    \I__1486\ : InMux
    port map (
            O => \N__14289\,
            I => \N__14284\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__14284\,
            I => \tok.A_stk.tail_78\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__14281\,
            I => \N__14278\
        );

    \I__1483\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14272\
        );

    \I__1482\ : InMux
    port map (
            O => \N__14277\,
            I => \N__14272\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__14272\,
            I => \tok.A_stk.tail_62\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__14269\,
            I => \N__14266\
        );

    \I__1479\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14260\
        );

    \I__1478\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14260\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__14260\,
            I => \tok.A_stk.tail_46\
        );

    \I__1476\ : InMux
    port map (
            O => \N__14257\,
            I => \N__14251\
        );

    \I__1475\ : InMux
    port map (
            O => \N__14256\,
            I => \N__14251\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__14251\,
            I => \tok.A_stk.tail_30\
        );

    \I__1473\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14244\
        );

    \I__1472\ : InMux
    port map (
            O => \N__14247\,
            I => \N__14241\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__14244\,
            I => \tok.A_stk.tail_14\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__14241\,
            I => \tok.A_stk.tail_14\
        );

    \I__1469\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14232\
        );

    \I__1468\ : InMux
    port map (
            O => \N__14235\,
            I => \N__14229\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__14232\,
            I => tail_127
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__14229\,
            I => tail_127
        );

    \I__1465\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14220\
        );

    \I__1464\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14217\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__14220\,
            I => tail_111
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__14217\,
            I => tail_111
        );

    \I__1461\ : InMux
    port map (
            O => \N__14212\,
            I => \N__14206\
        );

    \I__1460\ : InMux
    port map (
            O => \N__14211\,
            I => \N__14206\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__14206\,
            I => \tok.A_stk.tail_95\
        );

    \I__1458\ : InMux
    port map (
            O => \N__14203\,
            I => \N__14197\
        );

    \I__1457\ : InMux
    port map (
            O => \N__14202\,
            I => \N__14197\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__14197\,
            I => \tok.A_stk.tail_79\
        );

    \I__1455\ : InMux
    port map (
            O => \N__14194\,
            I => \N__14188\
        );

    \I__1454\ : InMux
    port map (
            O => \N__14193\,
            I => \N__14188\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__14188\,
            I => \tok.A_stk.tail_63\
        );

    \I__1452\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14179\
        );

    \I__1451\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14179\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__14179\,
            I => \tok.A_stk.tail_47\
        );

    \I__1449\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14170\
        );

    \I__1448\ : InMux
    port map (
            O => \N__14175\,
            I => \N__14170\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__14170\,
            I => \tok.A_stk.tail_31\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__14167\,
            I => \N__14164\
        );

    \I__1445\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14161\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__14161\,
            I => \N__14158\
        );

    \I__1443\ : Span12Mux_s2_h
    port map (
            O => \N__14158\,
            I => \N__14154\
        );

    \I__1442\ : InMux
    port map (
            O => \N__14157\,
            I => \N__14151\
        );

    \I__1441\ : Odrv12
    port map (
            O => \N__14154\,
            I => \tok.A_stk.tail_15\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__14151\,
            I => \tok.A_stk.tail_15\
        );

    \I__1439\ : InMux
    port map (
            O => \N__14146\,
            I => \N__14142\
        );

    \I__1438\ : InMux
    port map (
            O => \N__14145\,
            I => \N__14139\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__14142\,
            I => \tok.uart.txclkcounter_1\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__14139\,
            I => \tok.uart.txclkcounter_1\
        );

    \I__1435\ : InMux
    port map (
            O => \N__14134\,
            I => \tok.uart.n4830\
        );

    \I__1434\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14127\
        );

    \I__1433\ : InMux
    port map (
            O => \N__14130\,
            I => \N__14124\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__14127\,
            I => \tok.uart.txclkcounter_2\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__14124\,
            I => \tok.uart.txclkcounter_2\
        );

    \I__1430\ : InMux
    port map (
            O => \N__14119\,
            I => \tok.uart.n4831\
        );

    \I__1429\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14112\
        );

    \I__1428\ : InMux
    port map (
            O => \N__14115\,
            I => \N__14109\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__14112\,
            I => \tok.uart.txclkcounter_3\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__14109\,
            I => \tok.uart.txclkcounter_3\
        );

    \I__1425\ : InMux
    port map (
            O => \N__14104\,
            I => \tok.uart.n4832\
        );

    \I__1424\ : InMux
    port map (
            O => \N__14101\,
            I => \N__14097\
        );

    \I__1423\ : InMux
    port map (
            O => \N__14100\,
            I => \N__14094\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__14097\,
            I => \tok.uart.txclkcounter_4\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__14094\,
            I => \tok.uart.txclkcounter_4\
        );

    \I__1420\ : InMux
    port map (
            O => \N__14089\,
            I => \tok.uart.n4833\
        );

    \I__1419\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14082\
        );

    \I__1418\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14079\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__14082\,
            I => \tok.uart.txclkcounter_5\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__14079\,
            I => \tok.uart.txclkcounter_5\
        );

    \I__1415\ : InMux
    port map (
            O => \N__14074\,
            I => \tok.uart.n4834\
        );

    \I__1414\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14067\
        );

    \I__1413\ : InMux
    port map (
            O => \N__14070\,
            I => \N__14064\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__14067\,
            I => \tok.uart.txclkcounter_6\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__14064\,
            I => \tok.uart.txclkcounter_6\
        );

    \I__1410\ : InMux
    port map (
            O => \N__14059\,
            I => \tok.uart.n4835\
        );

    \I__1409\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14052\
        );

    \I__1408\ : InMux
    port map (
            O => \N__14055\,
            I => \N__14049\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__14052\,
            I => \tok.uart.txclkcounter_7\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__14049\,
            I => \tok.uart.txclkcounter_7\
        );

    \I__1405\ : InMux
    port map (
            O => \N__14044\,
            I => \tok.uart.n4836\
        );

    \I__1404\ : InMux
    port map (
            O => \N__14041\,
            I => \bfn_1_14_0_\
        );

    \I__1403\ : InMux
    port map (
            O => \N__14038\,
            I => \N__14034\
        );

    \I__1402\ : InMux
    port map (
            O => \N__14037\,
            I => \N__14031\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__14034\,
            I => \N__14028\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__14031\,
            I => \tok.uart.txclkcounter_8\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__14028\,
            I => \tok.uart.txclkcounter_8\
        );

    \I__1398\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14020\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__14020\,
            I => \tok.n206_adj_691\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__14017\,
            I => \tok.n212_adj_689_cascade_\
        );

    \I__1395\ : InMux
    port map (
            O => \N__14014\,
            I => \N__14008\
        );

    \I__1394\ : InMux
    port map (
            O => \N__14013\,
            I => \N__14008\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__14008\,
            I => \tok.n229_adj_863\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__14005\,
            I => \tok.uart.n6223_cascade_\
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__14002\,
            I => \txtick_cascade_\
        );

    \I__1390\ : InMux
    port map (
            O => \N__13999\,
            I => \N__13996\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__13996\,
            I => \tok.uart.n12\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__13993\,
            I => \N__13989\
        );

    \I__1387\ : InMux
    port map (
            O => \N__13992\,
            I => \N__13986\
        );

    \I__1386\ : InMux
    port map (
            O => \N__13989\,
            I => \N__13983\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__13986\,
            I => \tok.uart.txclkcounter_0\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__13983\,
            I => \tok.uart.txclkcounter_0\
        );

    \I__1383\ : InMux
    port map (
            O => \N__13978\,
            I => \bfn_1_13_0_\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__13975\,
            I => \tok.n203_adj_833_cascade_\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__13972\,
            I => \tok.n212_adj_835_cascade_\
        );

    \I__1380\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13966\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__13966\,
            I => \tok.n206_adj_834\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__13963\,
            I => \tok.n6443_cascade_\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__13960\,
            I => \tok.n242_adj_839_cascade_\
        );

    \I__1376\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13951\
        );

    \I__1375\ : InMux
    port map (
            O => \N__13956\,
            I => \N__13951\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__13951\,
            I => \tok.n230\
        );

    \I__1373\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13945\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__13945\,
            I => \tok.n242_adj_874\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__13942\,
            I => \tok.n6431_cascade_\
        );

    \I__1370\ : InMux
    port map (
            O => \N__13939\,
            I => \N__13936\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__13936\,
            I => \tok.n206_adj_869\
        );

    \I__1368\ : InMux
    port map (
            O => \N__13933\,
            I => \N__13930\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__13930\,
            I => \N__13927\
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__13927\,
            I => \tok.table_rd_13\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__13924\,
            I => \tok.n226_cascade_\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__13921\,
            I => \tok.n203_adj_643_cascade_\
        );

    \I__1363\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13915\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__13915\,
            I => \tok.n226\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__13912\,
            I => \tok.n212_adj_646_cascade_\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__13909\,
            I => \tok.n6448_cascade_\
        );

    \I__1359\ : InMux
    port map (
            O => \N__13906\,
            I => \N__13903\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__13903\,
            I => \tok.n6388\
        );

    \I__1357\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13897\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__13897\,
            I => \tok.n206_adj_649\
        );

    \I__1355\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13891\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__13891\,
            I => \N__13888\
        );

    \I__1353\ : Span4Mux_v
    port map (
            O => \N__13888\,
            I => \N__13885\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__13885\,
            I => \tok.table_rd_9\
        );

    \I__1351\ : InMux
    port map (
            O => \N__13882\,
            I => \tok.n4773\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__13879\,
            I => \N__13875\
        );

    \I__1349\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13872\
        );

    \I__1348\ : InMux
    port map (
            O => \N__13875\,
            I => \N__13869\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__13872\,
            I => tail_120
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__13869\,
            I => tail_120
        );

    \I__1345\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13860\
        );

    \I__1344\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13857\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__13860\,
            I => tail_104
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__13857\,
            I => tail_104
        );

    \I__1341\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13848\
        );

    \I__1340\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13845\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__13848\,
            I => \tok.A_stk.tail_88\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__13845\,
            I => \tok.A_stk.tail_88\
        );

    \I__1337\ : InMux
    port map (
            O => \N__13840\,
            I => \N__13834\
        );

    \I__1336\ : InMux
    port map (
            O => \N__13839\,
            I => \N__13834\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__13834\,
            I => \tok.A_stk.tail_72\
        );

    \I__1334\ : InMux
    port map (
            O => \N__13831\,
            I => \N__13825\
        );

    \I__1333\ : InMux
    port map (
            O => \N__13830\,
            I => \N__13825\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__13825\,
            I => \tok.A_stk.tail_56\
        );

    \I__1331\ : InMux
    port map (
            O => \N__13822\,
            I => \N__13816\
        );

    \I__1330\ : InMux
    port map (
            O => \N__13821\,
            I => \N__13816\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__13816\,
            I => \tok.A_stk.tail_40\
        );

    \I__1328\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13807\
        );

    \I__1327\ : InMux
    port map (
            O => \N__13812\,
            I => \N__13807\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__13807\,
            I => \tok.A_stk.tail_24\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__13804\,
            I => \N__13801\
        );

    \I__1324\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13795\
        );

    \I__1323\ : InMux
    port map (
            O => \N__13800\,
            I => \N__13795\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__13795\,
            I => \tok.A_stk.tail_8\
        );

    \I__1321\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13789\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__13789\,
            I => \N__13785\
        );

    \I__1319\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13782\
        );

    \I__1318\ : Odrv12
    port map (
            O => \N__13785\,
            I => \tok.A_stk.tail_0\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__13782\,
            I => \tok.A_stk.tail_0\
        );

    \I__1316\ : InMux
    port map (
            O => \N__13777\,
            I => \N__13771\
        );

    \I__1315\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13771\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__13771\,
            I => \tok.A_stk.tail_4\
        );

    \I__1313\ : InMux
    port map (
            O => \N__13768\,
            I => \bfn_1_7_0_\
        );

    \I__1312\ : InMux
    port map (
            O => \N__13765\,
            I => \tok.n4767\
        );

    \I__1311\ : InMux
    port map (
            O => \N__13762\,
            I => \tok.n4768\
        );

    \I__1310\ : InMux
    port map (
            O => \N__13759\,
            I => \tok.n4769\
        );

    \I__1309\ : InMux
    port map (
            O => \N__13756\,
            I => \tok.n4770\
        );

    \I__1308\ : InMux
    port map (
            O => \N__13753\,
            I => \tok.n4771\
        );

    \I__1307\ : InMux
    port map (
            O => \N__13750\,
            I => \tok.n4772\
        );

    \I__1306\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13744\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13741\
        );

    \I__1304\ : Span4Mux_h
    port map (
            O => \N__13741\,
            I => \N__13737\
        );

    \I__1303\ : InMux
    port map (
            O => \N__13740\,
            I => \N__13734\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__13737\,
            I => tail_101
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__13734\,
            I => tail_101
        );

    \I__1300\ : InMux
    port map (
            O => \N__13729\,
            I => \N__13726\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__13726\,
            I => \N__13722\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__13725\,
            I => \N__13719\
        );

    \I__1297\ : Span4Mux_s2_h
    port map (
            O => \N__13722\,
            I => \N__13716\
        );

    \I__1296\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13713\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__13716\,
            I => tail_117
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__13713\,
            I => tail_117
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__13708\,
            I => \N__13705\
        );

    \I__1292\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13702\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__13702\,
            I => \tok.n34\
        );

    \I__1290\ : InMux
    port map (
            O => \N__13699\,
            I => \N__13696\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__13696\,
            I => \N__13692\
        );

    \I__1288\ : InMux
    port map (
            O => \N__13695\,
            I => \N__13689\
        );

    \I__1287\ : Span4Mux_v
    port map (
            O => \N__13692\,
            I => \N__13686\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__13689\,
            I => tail_100
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__13686\,
            I => tail_100
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__13681\,
            I => \rd_15__N_300_cascade_\
        );

    \I__1283\ : InMux
    port map (
            O => \N__13678\,
            I => \N__13674\
        );

    \I__1282\ : InMux
    port map (
            O => \N__13677\,
            I => \N__13671\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__13674\,
            I => tail_116
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__13671\,
            I => tail_116
        );

    \I__1279\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13662\
        );

    \I__1278\ : InMux
    port map (
            O => \N__13665\,
            I => \N__13659\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__13662\,
            I => \tok.A_stk.tail_91\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__13659\,
            I => \tok.A_stk.tail_91\
        );

    \I__1275\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13650\
        );

    \I__1274\ : InMux
    port map (
            O => \N__13653\,
            I => \N__13647\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__13650\,
            I => tail_123
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__13647\,
            I => tail_123
        );

    \I__1271\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13638\
        );

    \I__1270\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13635\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__13638\,
            I => tail_107
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__13635\,
            I => tail_107
        );

    \I__1267\ : InMux
    port map (
            O => \N__13630\,
            I => \N__13626\
        );

    \I__1266\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13623\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__13626\,
            I => \N__13620\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__13623\,
            I => \N__13617\
        );

    \I__1263\ : Span4Mux_h
    port map (
            O => \N__13620\,
            I => \N__13614\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__13617\,
            I => \tok.A_stk.tail_84\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__13614\,
            I => \tok.A_stk.tail_84\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__13609\,
            I => \N__13605\
        );

    \I__1259\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13602\
        );

    \I__1258\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13599\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__13602\,
            I => \tok.A_stk.tail_68\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__13599\,
            I => \tok.A_stk.tail_68\
        );

    \I__1255\ : InMux
    port map (
            O => \N__13594\,
            I => \N__13588\
        );

    \I__1254\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13588\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__13588\,
            I => \tok.A_stk.tail_52\
        );

    \I__1252\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13579\
        );

    \I__1251\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13579\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__13579\,
            I => \tok.A_stk.tail_36\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__13576\,
            I => \N__13573\
        );

    \I__1248\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13567\
        );

    \I__1247\ : InMux
    port map (
            O => \N__13572\,
            I => \N__13567\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__13567\,
            I => \tok.A_stk.tail_20\
        );

    \I__1245\ : InMux
    port map (
            O => \N__13564\,
            I => \N__13560\
        );

    \I__1244\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13557\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__13560\,
            I => \N__13554\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__13557\,
            I => tail_106
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__13554\,
            I => tail_106
        );

    \I__1240\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13543\
        );

    \I__1239\ : InMux
    port map (
            O => \N__13548\,
            I => \N__13543\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__13543\,
            I => \tok.A_stk.tail_90\
        );

    \I__1237\ : InMux
    port map (
            O => \N__13540\,
            I => \N__13536\
        );

    \I__1236\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13533\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__13536\,
            I => \tok.A_stk.tail_74\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__13533\,
            I => \tok.A_stk.tail_74\
        );

    \I__1233\ : InMux
    port map (
            O => \N__13528\,
            I => \N__13522\
        );

    \I__1232\ : InMux
    port map (
            O => \N__13527\,
            I => \N__13522\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__13522\,
            I => \tok.A_stk.tail_58\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__13519\,
            I => \N__13516\
        );

    \I__1229\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13510\
        );

    \I__1228\ : InMux
    port map (
            O => \N__13515\,
            I => \N__13510\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__13510\,
            I => \tok.A_stk.tail_42\
        );

    \I__1226\ : InMux
    port map (
            O => \N__13507\,
            I => \N__13503\
        );

    \I__1225\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13500\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__13503\,
            I => tail_109
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__13500\,
            I => tail_109
        );

    \I__1222\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13491\
        );

    \I__1221\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13488\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__13491\,
            I => tail_125
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__13488\,
            I => tail_125
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__13483\,
            I => \N__13480\
        );

    \I__1217\ : InMux
    port map (
            O => \N__13480\,
            I => \N__13477\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__13477\,
            I => \N__13474\
        );

    \I__1215\ : Odrv4
    port map (
            O => \N__13474\,
            I => \tok.n6274\
        );

    \I__1214\ : CascadeMux
    port map (
            O => \N__13471\,
            I => \tok.n34_cascade_\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__13468\,
            I => \A_stk_delta_1_cascade_\
        );

    \I__1212\ : InMux
    port map (
            O => \N__13465\,
            I => \N__13461\
        );

    \I__1211\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13458\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__13461\,
            I => \N__13455\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__13458\,
            I => \N__13452\
        );

    \I__1208\ : Odrv4
    port map (
            O => \N__13455\,
            I => tail_105
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__13452\,
            I => tail_105
        );

    \I__1206\ : InMux
    port map (
            O => \N__13447\,
            I => \N__13444\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__13444\,
            I => \N__13440\
        );

    \I__1204\ : InMux
    port map (
            O => \N__13443\,
            I => \N__13437\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__13440\,
            I => tail_121
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__13437\,
            I => tail_121
        );

    \I__1201\ : InMux
    port map (
            O => \N__13432\,
            I => \N__13428\
        );

    \I__1200\ : InMux
    port map (
            O => \N__13431\,
            I => \N__13425\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__13428\,
            I => tail_96
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__13425\,
            I => tail_96
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__13420\,
            I => \N__13416\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__13419\,
            I => \N__13413\
        );

    \I__1195\ : InMux
    port map (
            O => \N__13416\,
            I => \N__13410\
        );

    \I__1194\ : InMux
    port map (
            O => \N__13413\,
            I => \N__13407\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__13410\,
            I => tail_112
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__13407\,
            I => tail_112
        );

    \I__1191\ : InMux
    port map (
            O => \N__13402\,
            I => \N__13398\
        );

    \I__1190\ : InMux
    port map (
            O => \N__13401\,
            I => \N__13395\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__13398\,
            I => \N__13392\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__13395\,
            I => \N__13389\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__13392\,
            I => tail_118
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__13389\,
            I => tail_118
        );

    \I__1185\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13381\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__13381\,
            I => \N__13378\
        );

    \I__1183\ : Span4Mux_v
    port map (
            O => \N__13378\,
            I => \N__13375\
        );

    \I__1182\ : Span4Mux_v
    port map (
            O => \N__13375\,
            I => \N__13372\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__13372\,
            I => \tok.table_wr_data_8\
        );

    \I__1180\ : InMux
    port map (
            O => \N__13369\,
            I => \N__13365\
        );

    \I__1179\ : InMux
    port map (
            O => \N__13368\,
            I => \N__13362\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__13365\,
            I => \N__13359\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__13362\,
            I => \tok.A_stk.tail_89\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__13359\,
            I => \tok.A_stk.tail_89\
        );

    \I__1175\ : InMux
    port map (
            O => \N__13354\,
            I => \N__13350\
        );

    \I__1174\ : InMux
    port map (
            O => \N__13353\,
            I => \N__13347\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__13350\,
            I => tail_122
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__13347\,
            I => tail_122
        );

    \I__1171\ : InMux
    port map (
            O => \N__13342\,
            I => \N__13336\
        );

    \I__1170\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13336\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__13336\,
            I => tail_80
        );

    \I__1168\ : InMux
    port map (
            O => \N__13333\,
            I => \N__13327\
        );

    \I__1167\ : InMux
    port map (
            O => \N__13332\,
            I => \N__13327\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__13327\,
            I => \tok.A_stk.tail_64\
        );

    \I__1165\ : InMux
    port map (
            O => \N__13324\,
            I => \N__13318\
        );

    \I__1164\ : InMux
    port map (
            O => \N__13323\,
            I => \N__13318\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__13318\,
            I => tail_48
        );

    \I__1162\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13309\
        );

    \I__1161\ : InMux
    port map (
            O => \N__13314\,
            I => \N__13309\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__13309\,
            I => \tok.A_stk.tail_32\
        );

    \I__1159\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13300\
        );

    \I__1158\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13300\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__13300\,
            I => tail_16
        );

    \I__1156\ : InMux
    port map (
            O => \N__13297\,
            I => \N__13291\
        );

    \I__1155\ : InMux
    port map (
            O => \N__13296\,
            I => \N__13291\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__13291\,
            I => \tok.A_stk.tail_9\
        );

    \I__1153\ : InMux
    port map (
            O => \N__13288\,
            I => \N__13282\
        );

    \I__1152\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13282\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__13282\,
            I => \tok.A_stk.tail_25\
        );

    \I__1150\ : InMux
    port map (
            O => \N__13279\,
            I => \N__13276\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__13276\,
            I => \N__13273\
        );

    \I__1148\ : Span4Mux_v
    port map (
            O => \N__13273\,
            I => \N__13269\
        );

    \I__1147\ : InMux
    port map (
            O => \N__13272\,
            I => \N__13266\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__13269\,
            I => \tok.A_stk.tail_57\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__13266\,
            I => \tok.A_stk.tail_57\
        );

    \I__1144\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13257\
        );

    \I__1143\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13254\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__13257\,
            I => \N__13251\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__13254\,
            I => \N__13248\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__13251\,
            I => \N__13245\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__13248\,
            I => \tok.A_stk.tail_41\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__13245\,
            I => \tok.A_stk.tail_41\
        );

    \I__1137\ : InMux
    port map (
            O => \N__13240\,
            I => \N__13237\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__13237\,
            I => \N__13234\
        );

    \I__1135\ : Span4Mux_v
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__13231\,
            I => \tok.table_rd_10\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__13228\,
            I => \tok.n203_adj_866_cascade_\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__13225\,
            I => \tok.n212_adj_867_cascade_\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__13222\,
            I => \tok.n6426_cascade_\
        );

    \I__1130\ : InMux
    port map (
            O => \N__13219\,
            I => \N__13213\
        );

    \I__1129\ : InMux
    port map (
            O => \N__13218\,
            I => \N__13213\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__13213\,
            I => \tok.A_stk.tail_85\
        );

    \I__1127\ : InMux
    port map (
            O => \N__13210\,
            I => \N__13204\
        );

    \I__1126\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13204\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__13204\,
            I => \tok.A_stk.tail_69\
        );

    \I__1124\ : InMux
    port map (
            O => \N__13201\,
            I => \N__13195\
        );

    \I__1123\ : InMux
    port map (
            O => \N__13200\,
            I => \N__13195\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__13195\,
            I => \tok.A_stk.tail_53\
        );

    \I__1121\ : InMux
    port map (
            O => \N__13192\,
            I => \N__13186\
        );

    \I__1120\ : InMux
    port map (
            O => \N__13191\,
            I => \N__13186\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__13186\,
            I => \tok.A_stk.tail_37\
        );

    \I__1118\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13179\
        );

    \I__1117\ : InMux
    port map (
            O => \N__13182\,
            I => \N__13176\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__13179\,
            I => \tok.A_stk.tail_21\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__13176\,
            I => \tok.A_stk.tail_21\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__13171\,
            I => \N__13168\
        );

    \I__1113\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13162\
        );

    \I__1112\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13162\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__13162\,
            I => \tok.A_stk.tail_5\
        );

    \I__1110\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13156\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__13156\,
            I => \N__13152\
        );

    \I__1108\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13149\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__13152\,
            I => \tok.A_stk.tail_11\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__13149\,
            I => \tok.A_stk.tail_11\
        );

    \I__1105\ : InMux
    port map (
            O => \N__13144\,
            I => \N__13138\
        );

    \I__1104\ : InMux
    port map (
            O => \N__13143\,
            I => \N__13138\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__13138\,
            I => \tok.A_stk.tail_29\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__13135\,
            I => \N__13132\
        );

    \I__1101\ : InMux
    port map (
            O => \N__13132\,
            I => \N__13126\
        );

    \I__1100\ : InMux
    port map (
            O => \N__13131\,
            I => \N__13126\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__13126\,
            I => \tok.A_stk.tail_13\
        );

    \I__1098\ : InMux
    port map (
            O => \N__13123\,
            I => \N__13117\
        );

    \I__1097\ : InMux
    port map (
            O => \N__13122\,
            I => \N__13117\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__13117\,
            I => \tok.A_stk.tail_75\
        );

    \I__1095\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13108\
        );

    \I__1094\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13108\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__13108\,
            I => \tok.A_stk.tail_59\
        );

    \I__1092\ : InMux
    port map (
            O => \N__13105\,
            I => \N__13099\
        );

    \I__1091\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13099\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__13099\,
            I => \tok.A_stk.tail_43\
        );

    \I__1089\ : InMux
    port map (
            O => \N__13096\,
            I => \N__13090\
        );

    \I__1088\ : InMux
    port map (
            O => \N__13095\,
            I => \N__13090\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__13090\,
            I => \tok.A_stk.tail_27\
        );

    \I__1086\ : InMux
    port map (
            O => \N__13087\,
            I => \N__13081\
        );

    \I__1085\ : InMux
    port map (
            O => \N__13086\,
            I => \N__13081\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__13081\,
            I => \tok.A_stk.tail_73\
        );

    \I__1083\ : InMux
    port map (
            O => \N__13078\,
            I => \N__13074\
        );

    \I__1082\ : InMux
    port map (
            O => \N__13077\,
            I => \N__13071\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__13074\,
            I => \tok.A_stk.tail_93\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__13071\,
            I => \tok.A_stk.tail_93\
        );

    \I__1079\ : InMux
    port map (
            O => \N__13066\,
            I => \N__13060\
        );

    \I__1078\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13060\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__13060\,
            I => \tok.A_stk.tail_77\
        );

    \I__1076\ : InMux
    port map (
            O => \N__13057\,
            I => \N__13051\
        );

    \I__1075\ : InMux
    port map (
            O => \N__13056\,
            I => \N__13051\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__13051\,
            I => \tok.A_stk.tail_61\
        );

    \I__1073\ : InMux
    port map (
            O => \N__13048\,
            I => \N__13042\
        );

    \I__1072\ : InMux
    port map (
            O => \N__13047\,
            I => \N__13042\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__13042\,
            I => \tok.A_stk.tail_45\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.uart.n4837\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4788_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4796\,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4781\,
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_6_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_2_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4803_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4810_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_4_11_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \OSCInst0\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b01"
        )
    port map (
            CLKHFPU => \N__17536\,
            CLKHFEN => \N__17535\,
            CLKHF => clk
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i57_LC_0_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13261\,
            in1 => \N__13087\,
            in2 => \_gnd_net_\,
            in3 => \N__18201\,
            lcout => \tok.A_stk.tail_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38428\,
            ce => \N__17919\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i89_LC_0_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13464\,
            in1 => \N__13086\,
            in2 => \_gnd_net_\,
            in3 => \N__18203\,
            lcout => \tok.A_stk.tail_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38428\,
            ce => \N__17919\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i73_LC_0_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18202\,
            in1 => \N__13368\,
            in2 => \_gnd_net_\,
            in3 => \N__13272\,
            lcout => \tok.A_stk.tail_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38428\,
            ce => \N__17919\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i109_LC_0_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13494\,
            in1 => \N__13077\,
            in2 => \_gnd_net_\,
            in3 => \N__18181\,
            lcout => tail_109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38431\,
            ce => \N__17936\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i93_LC_0_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18187\,
            in1 => \N__13506\,
            in2 => \_gnd_net_\,
            in3 => \N__13065\,
            lcout => \tok.A_stk.tail_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38431\,
            ce => \N__17936\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i77_LC_0_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13078\,
            in1 => \N__13056\,
            in2 => \_gnd_net_\,
            in3 => \N__18186\,
            lcout => \tok.A_stk.tail_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38431\,
            ce => \N__17936\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i61_LC_0_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18185\,
            in1 => \N__13047\,
            in2 => \_gnd_net_\,
            in3 => \N__13066\,
            lcout => \tok.A_stk.tail_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38431\,
            ce => \N__17936\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i45_LC_0_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13143\,
            in1 => \N__13057\,
            in2 => \_gnd_net_\,
            in3 => \N__18184\,
            lcout => \tok.A_stk.tail_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38431\,
            ce => \N__17936\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i29_LC_0_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__18183\,
            in1 => \_gnd_net_\,
            in2 => \N__13135\,
            in3 => \N__13048\,
            lcout => \tok.A_stk.tail_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38431\,
            ce => \N__17936\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i13_LC_0_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13144\,
            in1 => \N__18182\,
            in2 => \_gnd_net_\,
            in3 => \N__17288\,
            lcout => \tok.A_stk.tail_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38431\,
            ce => \N__17936\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i13_LC_0_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13131\,
            in1 => \N__18569\,
            in2 => \_gnd_net_\,
            in3 => \N__32232\,
            lcout => \tok.S_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38431\,
            ce => \N__17936\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i91_LC_0_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18194\,
            in1 => \N__13641\,
            in2 => \_gnd_net_\,
            in3 => \N__13122\,
            lcout => \tok.A_stk.tail_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38435\,
            ce => \N__17874\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i75_LC_0_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13666\,
            in1 => \N__13113\,
            in2 => \_gnd_net_\,
            in3 => \N__18192\,
            lcout => \tok.A_stk.tail_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38435\,
            ce => \N__17874\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i59_LC_0_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18191\,
            in1 => \N__13104\,
            in2 => \_gnd_net_\,
            in3 => \N__13123\,
            lcout => \tok.A_stk.tail_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38435\,
            ce => \N__17874\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i43_LC_0_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13095\,
            in1 => \N__13114\,
            in2 => \_gnd_net_\,
            in3 => \N__18190\,
            lcout => \tok.A_stk.tail_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38435\,
            ce => \N__17874\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i27_LC_0_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18189\,
            in1 => \N__13155\,
            in2 => \_gnd_net_\,
            in3 => \N__13105\,
            lcout => \tok.A_stk.tail_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38435\,
            ce => \N__17874\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i11_LC_0_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13096\,
            in1 => \N__18188\,
            in2 => \_gnd_net_\,
            in3 => \N__19470\,
            lcout => \tok.A_stk.tail_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38435\,
            ce => \N__17874\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i84_LC_0_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__18193\,
            in1 => \_gnd_net_\,
            in2 => \N__13609\,
            in3 => \N__13699\,
            lcout => \tok.A_stk.tail_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38435\,
            ce => \N__17874\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i101_LC_0_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13729\,
            in1 => \N__13218\,
            in2 => \_gnd_net_\,
            in3 => \N__18356\,
            lcout => tail_101,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38440\,
            ce => \N__17946\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i85_LC_0_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18362\,
            in1 => \N__13740\,
            in2 => \_gnd_net_\,
            in3 => \N__13209\,
            lcout => \tok.A_stk.tail_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38440\,
            ce => \N__17946\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i69_LC_0_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13200\,
            in1 => \N__13219\,
            in2 => \_gnd_net_\,
            in3 => \N__18361\,
            lcout => \tok.A_stk.tail_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38440\,
            ce => \N__17946\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i53_LC_0_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18359\,
            in1 => \N__13210\,
            in2 => \_gnd_net_\,
            in3 => \N__13191\,
            lcout => \tok.A_stk.tail_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38440\,
            ce => \N__17946\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i37_LC_0_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13201\,
            in1 => \N__13182\,
            in2 => \_gnd_net_\,
            in3 => \N__18358\,
            lcout => \tok.A_stk.tail_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38440\,
            ce => \N__17946\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i21_LC_0_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__18357\,
            in1 => \_gnd_net_\,
            in2 => \N__13171\,
            in3 => \N__13192\,
            lcout => \tok.A_stk.tail_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38440\,
            ce => \N__17946\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i5_LC_0_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13183\,
            in1 => \N__18360\,
            in2 => \_gnd_net_\,
            in3 => \N__21986\,
            lcout => \tok.A_stk.tail_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38440\,
            ce => \N__17946\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i5_LC_0_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13167\,
            in1 => \N__18586\,
            in2 => \_gnd_net_\,
            in3 => \N__30343\,
            lcout => \tok.S_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38440\,
            ce => \N__17946\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i11_LC_0_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13159\,
            in1 => \N__18587\,
            in2 => \_gnd_net_\,
            in3 => \N__24000\,
            lcout => \tok.S_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38445\,
            ce => \N__17923\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i9_LC_0_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13296\,
            in1 => \N__18588\,
            in2 => \_gnd_net_\,
            in3 => \N__26803\,
            lcout => \tok.S_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38445\,
            ce => \N__17923\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i15_LC_0_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24198\,
            in2 => \N__14167\,
            in3 => \N__18589\,
            lcout => \tok.S_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38445\,
            ce => \N__17923\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i9_LC_0_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18347\,
            in1 => \N__13288\,
            in2 => \_gnd_net_\,
            in3 => \N__21737\,
            lcout => \tok.A_stk.tail_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38445\,
            ce => \N__17923\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i25_LC_0_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13260\,
            in1 => \N__13297\,
            in2 => \_gnd_net_\,
            in3 => \N__18345\,
            lcout => \tok.A_stk.tail_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38445\,
            ce => \N__17923\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i41_LC_0_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18346\,
            in1 => \N__13287\,
            in2 => \_gnd_net_\,
            in3 => \N__13279\,
            lcout => \tok.A_stk.tail_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38445\,
            ce => \N__17923\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i120_LC_0_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__18348\,
            in1 => \N__13864\,
            in2 => \N__13879\,
            in3 => \N__17935\,
            lcout => tail_120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i312_4_lut_adj_301_LC_0_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__13240\,
            in1 => \N__33097\,
            in2 => \N__31214\,
            in3 => \N__14013\,
            lcout => OPEN,
            ltout => \tok.n203_adj_866_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_302_LC_0_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__14014\,
            in1 => \N__19246\,
            in2 => \N__13228\,
            in3 => \N__31940\,
            lcout => OPEN,
            ltout => \tok.n212_adj_867_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6917_4_lut_LC_0_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__31941\,
            in1 => \N__33430\,
            in2 => \N__13225\,
            in3 => \N__13939\,
            lcout => OPEN,
            ltout => \tok.n6426_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_309_LC_0_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__26182\,
            in1 => \N__36981\,
            in2 => \N__13222\,
            in3 => \N__30322\,
            lcout => \tok.n242_adj_874\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i300_4_lut_4_lut_LC_0_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__20689\,
            in1 => \N__35972\,
            in2 => \N__24197\,
            in3 => \N__14866\,
            lcout => \tok.n206_adj_691\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i96_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18372\,
            in1 => \_gnd_net_\,
            in2 => \N__13420\,
            in3 => \N__13341\,
            lcout => tail_96,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38426\,
            ce => \N__17900\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i80_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13431\,
            in1 => \N__13332\,
            in2 => \_gnd_net_\,
            in3 => \N__18371\,
            lcout => tail_80,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38426\,
            ce => \N__17900\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i64_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18370\,
            in1 => \N__13342\,
            in2 => \_gnd_net_\,
            in3 => \N__13323\,
            lcout => \tok.A_stk.tail_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38426\,
            ce => \N__17900\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i48_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13314\,
            in1 => \N__13333\,
            in2 => \_gnd_net_\,
            in3 => \N__18369\,
            lcout => tail_48,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38426\,
            ce => \N__17900\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i32_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18368\,
            in1 => \N__13305\,
            in2 => \_gnd_net_\,
            in3 => \N__13324\,
            lcout => \tok.A_stk.tail_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38426\,
            ce => \N__17900\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i16_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13315\,
            in1 => \N__13788\,
            in2 => \_gnd_net_\,
            in3 => \N__18367\,
            lcout => tail_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38426\,
            ce => \N__17900\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i0_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18365\,
            in1 => \N__13306\,
            in2 => \_gnd_net_\,
            in3 => \N__18813\,
            lcout => \tok.A_stk.tail_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38426\,
            ce => \N__17900\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i102_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13402\,
            in1 => \N__15016\,
            in2 => \_gnd_net_\,
            in3 => \N__18366\,
            lcout => tail_102,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38426\,
            ce => \N__17900\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i112_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__13432\,
            in1 => \N__17813\,
            in2 => \N__13419\,
            in3 => \N__18216\,
            lcout => tail_112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i122_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18218\,
            in1 => \N__13353\,
            in2 => \N__17885\,
            in3 => \N__13563\,
            lcout => tail_122,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7005_4_lut_4_lut_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001100010011"
        )
    port map (
            in0 => \N__31939\,
            in1 => \N__33296\,
            in2 => \N__34840\,
            in3 => \N__31296\,
            lcout => \tok.n6274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i118_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18217\,
            in1 => \N__13401\,
            in2 => \N__17884\,
            in3 => \N__15030\,
            lcout => tail_118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i126_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__18219\,
            in1 => \N__14320\,
            in2 => \N__17886\,
            in3 => \N__14331\,
            lcout => tail_126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2626_2_lut_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28474\,
            in2 => \_gnd_net_\,
            in3 => \N__17249\,
            lcout => \tok.table_wr_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i105_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13447\,
            in1 => \N__13369\,
            in2 => \_gnd_net_\,
            in3 => \N__18168\,
            lcout => tail_105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__17932\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i26_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18170\,
            in1 => \_gnd_net_\,
            in2 => \N__13519\,
            in3 => \N__15202\,
            lcout => \tok.A_stk.tail_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__17932\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i100_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13678\,
            in1 => \N__13630\,
            in2 => \_gnd_net_\,
            in3 => \N__18167\,
            lcout => tail_100,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__17932\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i106_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18169\,
            in1 => \N__13354\,
            in2 => \_gnd_net_\,
            in3 => \N__13548\,
            lcout => tail_106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__17932\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i90_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13564\,
            in1 => \N__13539\,
            in2 => \_gnd_net_\,
            in3 => \N__18174\,
            lcout => \tok.A_stk.tail_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__17932\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i74_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18173\,
            in1 => \N__13549\,
            in2 => \_gnd_net_\,
            in3 => \N__13527\,
            lcout => \tok.A_stk.tail_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__17932\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i58_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13540\,
            in1 => \N__13515\,
            in2 => \_gnd_net_\,
            in3 => \N__18172\,
            lcout => \tok.A_stk.tail_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__17932\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i42_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18171\,
            in1 => \N__14346\,
            in2 => \_gnd_net_\,
            in3 => \N__13528\,
            lcout => \tok.A_stk.tail_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__17932\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i125_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__18116\,
            in1 => \N__13507\,
            in2 => \N__17812\,
            in3 => \N__13495\,
            lcout => tail_125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i49_4_lut_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__15328\,
            in1 => \N__35480\,
            in2 => \N__13483\,
            in3 => \N__36227\,
            lcout => \tok.n34\,
            ltout => \tok.n34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2541_2_lut_4_lut_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21348\,
            in1 => \N__32433\,
            in2 => \N__13471\,
            in3 => \N__25254\,
            lcout => \A_stk_delta_1\,
            ltout => \A_stk_delta_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i123_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__13653\,
            in1 => \N__13642\,
            in2 => \N__13468\,
            in3 => \N__17753\,
            lcout => tail_123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i121_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__18115\,
            in1 => \N__13443\,
            in2 => \N__17811\,
            in3 => \N__13465\,
            lcout => tail_121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i117_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__13747\,
            in1 => \N__17749\,
            in2 => \N__13725\,
            in3 => \N__18114\,
            lcout => tail_117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i426_2_lut_4_lut_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010101"
        )
    port map (
            in0 => \N__21349\,
            in1 => \N__32434\,
            in2 => \N__13708\,
            in3 => \N__25255\,
            lcout => \rd_15__N_300\,
            ltout => \rd_15__N_300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i116_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__13695\,
            in1 => \N__13677\,
            in2 => \N__13681\,
            in3 => \N__18113\,
            lcout => tail_116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i107_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13665\,
            in1 => \N__13654\,
            in2 => \_gnd_net_\,
            in3 => \N__18175\,
            lcout => tail_107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__17933\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i4_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18178\,
            in1 => \_gnd_net_\,
            in2 => \N__13576\,
            in3 => \N__23800\,
            lcout => \tok.A_stk.tail_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__17933\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i68_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13593\,
            in1 => \N__13629\,
            in2 => \_gnd_net_\,
            in3 => \N__18180\,
            lcout => \tok.A_stk.tail_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__17933\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i52_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18179\,
            in1 => \N__13584\,
            in2 => \_gnd_net_\,
            in3 => \N__13608\,
            lcout => \tok.A_stk.tail_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__17933\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i36_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13594\,
            in1 => \N__13572\,
            in2 => \_gnd_net_\,
            in3 => \N__18177\,
            lcout => \tok.A_stk.tail_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__17933\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i20_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18176\,
            in1 => \N__13585\,
            in2 => \_gnd_net_\,
            in3 => \N__13777\,
            lcout => \tok.A_stk.tail_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__17933\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i0_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13792\,
            in1 => \N__18581\,
            in2 => \_gnd_net_\,
            in3 => \N__30526\,
            lcout => \S_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__17933\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i4_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18582\,
            in1 => \N__13776\,
            in2 => \_gnd_net_\,
            in3 => \N__27390\,
            lcout => \tok.S_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__17933\,
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_2_lut_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__14515\,
            in1 => \N__14514\,
            in2 => \N__15739\,
            in3 => \N__13768\,
            lcout => \tok.n33_adj_631\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \tok.n4767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_3_lut_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__15461\,
            in1 => \N__15460\,
            in2 => \N__15723\,
            in3 => \N__13765\,
            lcout => \tok.n33_adj_632\,
            ltout => OPEN,
            carryin => \tok.n4767\,
            carryout => \tok.n4768\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_4_lut_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__15632\,
            in1 => \N__15631\,
            in2 => \N__15740\,
            in3 => \N__13762\,
            lcout => \tok.n33_adj_633\,
            ltout => OPEN,
            carryin => \tok.n4768\,
            carryout => \tok.n4769\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_5_lut_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__15542\,
            in1 => \N__15532\,
            in2 => \N__15724\,
            in3 => \N__13759\,
            lcout => \tok.n33_adj_661\,
            ltout => OPEN,
            carryin => \tok.n4769\,
            carryout => \tok.n4770\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_6_lut_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__14683\,
            in1 => \N__14682\,
            in2 => \N__15741\,
            in3 => \N__13756\,
            lcout => \tok.n33_adj_634\,
            ltout => OPEN,
            carryin => \tok.n4770\,
            carryout => \tok.n4771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_7_lut_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__15397\,
            in1 => \N__15398\,
            in2 => \N__15725\,
            in3 => \N__13753\,
            lcout => \tok.n33\,
            ltout => OPEN,
            carryin => \tok.n4771\,
            carryout => \tok.n4772\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_8_lut_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__15845\,
            in1 => \N__15844\,
            in2 => \N__15742\,
            in3 => \N__13750\,
            lcout => \tok.n33_adj_663\,
            ltout => OPEN,
            carryin => \tok.n4772\,
            carryout => \tok.n4773\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_9_lut_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__14451\,
            in1 => \N__14452\,
            in2 => \N__15726\,
            in3 => \N__13882\,
            lcout => \tok.n33_adj_662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i104_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13878\,
            in1 => \N__13851\,
            in2 => \_gnd_net_\,
            in3 => \N__18349\,
            lcout => tail_104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38450\,
            ce => \N__17926\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i88_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18354\,
            in1 => \N__13863\,
            in2 => \_gnd_net_\,
            in3 => \N__13839\,
            lcout => \tok.A_stk.tail_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38450\,
            ce => \N__17926\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i72_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13852\,
            in1 => \N__13830\,
            in2 => \_gnd_net_\,
            in3 => \N__18353\,
            lcout => \tok.A_stk.tail_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38450\,
            ce => \N__17926\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i56_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18352\,
            in1 => \N__13840\,
            in2 => \_gnd_net_\,
            in3 => \N__13821\,
            lcout => \tok.A_stk.tail_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38450\,
            ce => \N__17926\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i40_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13812\,
            in1 => \N__13831\,
            in2 => \_gnd_net_\,
            in3 => \N__18351\,
            lcout => \tok.A_stk.tail_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38450\,
            ce => \N__17926\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i24_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__18350\,
            in1 => \_gnd_net_\,
            in2 => \N__13804\,
            in3 => \N__13822\,
            lcout => \tok.A_stk.tail_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38450\,
            ce => \N__17926\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i8_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13813\,
            in1 => \N__18355\,
            in2 => \_gnd_net_\,
            in3 => \N__17220\,
            lcout => \tok.A_stk.tail_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38450\,
            ce => \N__17926\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i8_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13800\,
            in1 => \N__18583\,
            in2 => \_gnd_net_\,
            in3 => \N__22251\,
            lcout => \tok.S_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38450\,
            ce => \N__17926\,
            sr => \_gnd_net_\
        );

    \tok.or_100_i14_2_lut_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26797\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20767\,
            lcout => \tok.n226\,
            ltout => \tok.n226_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i312_4_lut_adj_34_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__13933\,
            in1 => \N__33098\,
            in2 => \N__13924\,
            in3 => \N__30972\,
            lcout => OPEN,
            ltout => \tok.n203_adj_643_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_37_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__31919\,
            in1 => \N__19247\,
            in2 => \N__13921\,
            in3 => \N__13918\,
            lcout => OPEN,
            ltout => \tok.n212_adj_646_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6897_4_lut_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__33415\,
            in1 => \N__31920\,
            in2 => \N__13912\,
            in3 => \N__13900\,
            lcout => \tok.n6383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6700_3_lut_4_lut_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__30970\,
            in1 => \N__34537\,
            in2 => \N__26802\,
            in3 => \N__20766\,
            lcout => \tok.n6388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6738_3_lut_4_lut_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__20768\,
            in1 => \N__30344\,
            in2 => \N__34706\,
            in3 => \N__30971\,
            lcout => OPEN,
            ltout => \tok.n6448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i300_4_lut_adj_265_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__36048\,
            in1 => \N__20679\,
            in2 => \N__13909\,
            in3 => \N__26798\,
            lcout => \tok.n206_adj_834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i300_4_lut_adj_39_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__20678\,
            in1 => \N__16927\,
            in2 => \N__36228\,
            in3 => \N__13906\,
            lcout => \tok.n206_adj_649\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i312_4_lut_adj_259_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__13894\,
            in1 => \N__33099\,
            in2 => \N__31215\,
            in3 => \N__13956\,
            lcout => OPEN,
            ltout => \tok.n203_adj_833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_326_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__13957\,
            in1 => \N__31931\,
            in2 => \N__13975\,
            in3 => \N__19244\,
            lcout => OPEN,
            ltout => \tok.n212_adj_835_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6922_4_lut_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__31932\,
            in1 => \N__33372\,
            in2 => \N__13972\,
            in3 => \N__13969\,
            lcout => OPEN,
            ltout => \tok.n6443_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_269_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__26181\,
            in1 => \N__27363\,
            in2 => \N__13963\,
            in3 => \N__36982\,
            lcout => OPEN,
            ltout => \tok.n242_adj_839_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_270_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__36983\,
            in1 => \N__16072\,
            in2 => \N__13960\,
            in3 => \N__35446\,
            lcout => \tok.n200_adj_840\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_100_i10_2_lut_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30321\,
            in2 => \_gnd_net_\,
            in3 => \N__20765\,
            lcout => \tok.n230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_310_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__35445\,
            in1 => \N__36984\,
            in2 => \N__19039\,
            in3 => \N__13948\,
            lcout => \tok.n200_adj_875\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6730_3_lut_4_lut_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__34547\,
            in1 => \N__30973\,
            in2 => \N__20781\,
            in3 => \N__30084\,
            lcout => OPEN,
            ltout => \tok.n6431_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i300_4_lut_adj_304_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__20656\,
            in1 => \N__35778\,
            in2 => \N__13942\,
            in3 => \N__29627\,
            lcout => \tok.n206_adj_869\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_238_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33798\,
            in2 => \_gnd_net_\,
            in3 => \N__36897\,
            lcout => \tok.n9_adj_677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_74_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__31917\,
            in1 => \N__14917\,
            in2 => \N__19251\,
            in3 => \N__14896\,
            lcout => OPEN,
            ltout => \tok.n212_adj_689_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6880_4_lut_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__14023\,
            in1 => \N__33445\,
            in2 => \N__14017\,
            in3 => \N__31918\,
            lcout => \tok.n6347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_100_i11_2_lut_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30083\,
            in2 => \_gnd_net_\,
            in3 => \N__20761\,
            lcout => \tok.n229_adj_863\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i6139_3_lut_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14055\,
            in1 => \N__14070\,
            in2 => \_gnd_net_\,
            in3 => \N__14100\,
            lcout => OPEN,
            ltout => \tok.uart.n6223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i7019_4_lut_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__14115\,
            in1 => \N__14130\,
            in2 => \N__14005\,
            in3 => \N__13999\,
            lcout => txtick,
            ltout => \txtick_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i7027_2_lut_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14002\,
            in3 => \N__37556\,
            lcout => \tok.uart.n950\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i2_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__14964\,
            in1 => \N__37591\,
            in2 => \N__17398\,
            in3 => \N__37557\,
            lcout => sender_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i5_4_lut_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14038\,
            in1 => \N__14145\,
            in2 => \N__13993\,
            in3 => \N__14085\,
            lcout => \tok.uart.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_70_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__35267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30785\,
            lcout => \tok.n4_adj_636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.txclkcounter_141__i0_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13992\,
            in2 => \_gnd_net_\,
            in3 => \N__13978\,
            lcout => \tok.uart.txclkcounter_0\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \tok.uart.n4830\,
            clk => \N__38477\,
            ce => 'H',
            sr => \N__37607\
        );

    \tok.uart.txclkcounter_141__i1_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14146\,
            in2 => \_gnd_net_\,
            in3 => \N__14134\,
            lcout => \tok.uart.txclkcounter_1\,
            ltout => OPEN,
            carryin => \tok.uart.n4830\,
            carryout => \tok.uart.n4831\,
            clk => \N__38477\,
            ce => 'H',
            sr => \N__37607\
        );

    \tok.uart.txclkcounter_141__i2_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14131\,
            in2 => \_gnd_net_\,
            in3 => \N__14119\,
            lcout => \tok.uart.txclkcounter_2\,
            ltout => OPEN,
            carryin => \tok.uart.n4831\,
            carryout => \tok.uart.n4832\,
            clk => \N__38477\,
            ce => 'H',
            sr => \N__37607\
        );

    \tok.uart.txclkcounter_141__i3_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14116\,
            in2 => \_gnd_net_\,
            in3 => \N__14104\,
            lcout => \tok.uart.txclkcounter_3\,
            ltout => OPEN,
            carryin => \tok.uart.n4832\,
            carryout => \tok.uart.n4833\,
            clk => \N__38477\,
            ce => 'H',
            sr => \N__37607\
        );

    \tok.uart.txclkcounter_141__i4_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14101\,
            in2 => \_gnd_net_\,
            in3 => \N__14089\,
            lcout => \tok.uart.txclkcounter_4\,
            ltout => OPEN,
            carryin => \tok.uart.n4833\,
            carryout => \tok.uart.n4834\,
            clk => \N__38477\,
            ce => 'H',
            sr => \N__37607\
        );

    \tok.uart.txclkcounter_141__i5_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14086\,
            in2 => \_gnd_net_\,
            in3 => \N__14074\,
            lcout => \tok.uart.txclkcounter_5\,
            ltout => OPEN,
            carryin => \tok.uart.n4834\,
            carryout => \tok.uart.n4835\,
            clk => \N__38477\,
            ce => 'H',
            sr => \N__37607\
        );

    \tok.uart.txclkcounter_141__i6_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14071\,
            in2 => \_gnd_net_\,
            in3 => \N__14059\,
            lcout => \tok.uart.txclkcounter_6\,
            ltout => OPEN,
            carryin => \tok.uart.n4835\,
            carryout => \tok.uart.n4836\,
            clk => \N__38477\,
            ce => 'H',
            sr => \N__37607\
        );

    \tok.uart.txclkcounter_141__i7_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14056\,
            in2 => \_gnd_net_\,
            in3 => \N__14044\,
            lcout => \tok.uart.txclkcounter_7\,
            ltout => OPEN,
            carryin => \tok.uart.n4836\,
            carryout => \tok.uart.n4837\,
            clk => \N__38477\,
            ce => 'H',
            sr => \N__37607\
        );

    \tok.uart.txclkcounter_141__i8_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14037\,
            in2 => \_gnd_net_\,
            in3 => \N__14041\,
            lcout => \tok.uart.txclkcounter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38482\,
            ce => 'H',
            sr => \N__37601\
        );

    \tok.A_stk.tail_i0_i119_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__16243\,
            in1 => \N__17887\,
            in2 => \N__16260\,
            in3 => \N__18363\,
            lcout => tail_119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i127_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__18364\,
            in1 => \N__14224\,
            in2 => \N__17931\,
            in3 => \N__14235\,
            lcout => tail_127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i111_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18376\,
            in1 => \N__14236\,
            in2 => \_gnd_net_\,
            in3 => \N__14211\,
            lcout => tail_111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38430\,
            ce => \N__17901\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i95_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14223\,
            in1 => \N__18382\,
            in2 => \_gnd_net_\,
            in3 => \N__14202\,
            lcout => \tok.A_stk.tail_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38430\,
            ce => \N__17901\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i79_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18381\,
            in1 => \N__14212\,
            in2 => \_gnd_net_\,
            in3 => \N__14193\,
            lcout => \tok.A_stk.tail_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38430\,
            ce => \N__17901\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i63_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14184\,
            in1 => \N__18380\,
            in2 => \_gnd_net_\,
            in3 => \N__14203\,
            lcout => \tok.A_stk.tail_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38430\,
            ce => \N__17901\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i47_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18379\,
            in1 => \N__14175\,
            in2 => \_gnd_net_\,
            in3 => \N__14194\,
            lcout => \tok.A_stk.tail_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38430\,
            ce => \N__17901\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i31_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14185\,
            in1 => \N__18378\,
            in2 => \_gnd_net_\,
            in3 => \N__14157\,
            lcout => \tok.A_stk.tail_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38430\,
            ce => \N__17901\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i15_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18377\,
            in1 => \N__14176\,
            in2 => \_gnd_net_\,
            in3 => \N__18962\,
            lcout => \tok.A_stk.tail_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38430\,
            ce => \N__17901\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i10_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14350\,
            in1 => \N__18375\,
            in2 => \_gnd_net_\,
            in3 => \N__20178\,
            lcout => \tok.A_stk.tail_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38430\,
            ce => \N__17901\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i110_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14335\,
            in1 => \N__14301\,
            in2 => \_gnd_net_\,
            in3 => \N__18316\,
            lcout => tail_110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38433\,
            ce => \N__17948\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i94_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18322\,
            in1 => \N__14313\,
            in2 => \_gnd_net_\,
            in3 => \N__14289\,
            lcout => \tok.A_stk.tail_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38433\,
            ce => \N__17948\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i78_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14302\,
            in1 => \N__14277\,
            in2 => \_gnd_net_\,
            in3 => \N__18321\,
            lcout => \tok.A_stk.tail_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38433\,
            ce => \N__17948\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i46_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18319\,
            in1 => \_gnd_net_\,
            in2 => \N__14281\,
            in3 => \N__14256\,
            lcout => \tok.A_stk.tail_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38433\,
            ce => \N__17948\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i62_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14290\,
            in1 => \N__14265\,
            in2 => \_gnd_net_\,
            in3 => \N__18320\,
            lcout => \tok.A_stk.tail_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38433\,
            ce => \N__17948\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i30_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18318\,
            in1 => \_gnd_net_\,
            in2 => \N__14269\,
            in3 => \N__14248\,
            lcout => \tok.A_stk.tail_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38433\,
            ce => \N__17948\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i14_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14257\,
            in1 => \N__18317\,
            in2 => \_gnd_net_\,
            in3 => \N__19304\,
            lcout => \tok.A_stk.tail_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38433\,
            ce => \N__17948\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i14_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14247\,
            in1 => \N__18584\,
            in2 => \_gnd_net_\,
            in3 => \N__32380\,
            lcout => \tok.S_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38433\,
            ce => \N__17948\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i18_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14425\,
            in1 => \N__17974\,
            in2 => \_gnd_net_\,
            in3 => \N__18195\,
            lcout => \tok.A_stk.tail_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38437\,
            ce => \N__17934\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i34_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18196\,
            in1 => \N__18468\,
            in2 => \_gnd_net_\,
            in3 => \N__14416\,
            lcout => \tok.A_stk.tail_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38437\,
            ce => \N__17934\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i50_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14424\,
            in1 => \N__14407\,
            in2 => \_gnd_net_\,
            in3 => \N__18197\,
            lcout => \tok.A_stk.tail_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38437\,
            ce => \N__17934\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i66_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18198\,
            in1 => \N__14415\,
            in2 => \_gnd_net_\,
            in3 => \N__14398\,
            lcout => \tok.A_stk.tail_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38437\,
            ce => \N__17934\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i82_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14376\,
            in1 => \N__14406\,
            in2 => \_gnd_net_\,
            in3 => \N__18199\,
            lcout => \tok.A_stk.tail_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38437\,
            ce => \N__17934\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i98_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18200\,
            in1 => \N__14364\,
            in2 => \_gnd_net_\,
            in3 => \N__14397\,
            lcout => tail_98,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38437\,
            ce => \N__17934\,
            sr => \_gnd_net_\
        );

    \tok.i6975_2_lut_3_lut_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36220\,
            in1 => \N__33161\,
            in2 => \_gnd_net_\,
            in3 => \N__31285\,
            lcout => \tok.n6644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1412_3_lut_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__18812\,
            in1 => \_gnd_net_\,
            in2 => \N__28473\,
            in3 => \N__21172\,
            lcout => table_wr_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i114_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__14377\,
            in1 => \N__17757\,
            in2 => \N__14365\,
            in3 => \N__18117\,
            lcout => tail_114,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38442\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_adj_86_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__32967\,
            in1 => \N__31828\,
            in2 => \N__34560\,
            in3 => \N__31092\,
            lcout => \tok.n4_adj_642\,
            ltout => \tok.n4_adj_642_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6118_3_lut_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16568\,
            in2 => \N__14593\,
            in3 => \N__30145\,
            lcout => \tok.n2532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_adj_262_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__32966\,
            in1 => \N__31827\,
            in2 => \N__34559\,
            in3 => \N__31091\,
            lcout => \tok.n4_adj_641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2619_2_lut_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28450\,
            in2 => \_gnd_net_\,
            in3 => \N__17298\,
            lcout => \tok.table_wr_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2622_2_lut_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28451\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20177\,
            lcout => \tok.table_wr_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2617_2_lut_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18951\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28449\,
            lcout => \tok.table_wr_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__25360\,
            in1 => \N__14551\,
            in2 => \N__30535\,
            in3 => \N__15801\,
            lcout => OPEN,
            ltout => \tok.n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__14516\,
            in1 => \N__16779\,
            in2 => \N__14545\,
            in3 => \N__16677\,
            lcout => \tok.n41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38446\,
            ce => 'H',
            sr => \N__29254\
        );

    \tok.i50_4_lut_adj_100_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__14488\,
            in1 => \N__15797\,
            in2 => \N__25375\,
            in3 => \N__37467\,
            lcout => OPEN,
            ltout => \tok.n27_adj_709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i7_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__14453\,
            in1 => \N__16780\,
            in2 => \N__14482\,
            in3 => \N__16678\,
            lcout => \tok.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38446\,
            ce => 'H',
            sr => \N__29254\
        );

    \tok.i50_4_lut_adj_94_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__25353\,
            in1 => \N__14719\,
            in2 => \N__15802\,
            in3 => \N__27389\,
            lcout => OPEN,
            ltout => \tok.n27_adj_706_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i4_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__16671\,
            in1 => \N__14684\,
            in2 => \N__14713\,
            in3 => \N__16781\,
            lcout => \tok.n35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38446\,
            ce => 'H',
            sr => \N__29254\
        );

    \tok.i10_4_lut_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16608\,
            in1 => \N__16629\,
            in2 => \N__16884\,
            in3 => \N__16854\,
            lcout => \tok.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6974_4_lut_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16864\,
            in1 => \N__15676\,
            in2 => \N__14602\,
            in3 => \N__15916\,
            lcout => OPEN,
            ltout => \tok.n6667_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_41_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000101010"
        )
    port map (
            in0 => \N__25367\,
            in1 => \N__14767\,
            in2 => \N__14656\,
            in3 => \N__14653\,
            lcout => \tok.found_slot\,
            ltout => \tok.found_slot_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_4_lut_adj_291_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__14644\,
            in1 => \N__16576\,
            in2 => \N__14635\,
            in3 => \N__30134\,
            lcout => \tok.write_slot\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6632_3_lut_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__35260\,
            in1 => \N__14761\,
            in2 => \_gnd_net_\,
            in3 => \N__31826\,
            lcout => \tok.n6326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__29595\,
            in1 => \N__14799\,
            in2 => \N__14790\,
            in3 => \N__27039\,
            lcout => OPEN,
            ltout => \tok.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i14_4_lut_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14725\,
            in1 => \N__18673\,
            in2 => \N__14605\,
            in3 => \N__18715\,
            lcout => \tok.n30_adj_647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_100_i13_2_lut_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22241\,
            in2 => \_gnd_net_\,
            in3 => \N__20769\,
            lcout => \tok.n227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i11_4_lut_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14752\,
            in1 => \N__14800\,
            in2 => \N__14791\,
            in3 => \N__14739\,
            lcout => OPEN,
            ltout => \tok.n27_adj_639_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i15_4_lut_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15946\,
            in1 => \N__14776\,
            in2 => \N__14770\,
            in3 => \N__18766\,
            lcout => \tok.found_slot_N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6657_4_lut_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100111011"
        )
    port map (
            in0 => \N__36049\,
            in1 => \N__34710\,
            in2 => \N__33163\,
            in3 => \N__22242\,
            lcout => \tok.n6322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i13_1_lut_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27018\,
            lcout => \tok.n313\,
            ltout => \tok.n313_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i300_4_lut_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__20677\,
            in1 => \N__36044\,
            in2 => \N__14755\,
            in3 => \N__14854\,
            lcout => \tok.n206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__14751\,
            in1 => \N__37401\,
            in2 => \N__14740\,
            in3 => \N__33625\,
            lcout => \tok.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i11_1_lut_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29620\,
            lcout => \tok.n315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i8_1_lut_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37402\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i312_4_lut_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__14845\,
            in1 => \N__32851\,
            in2 => \N__31111\,
            in3 => \N__14835\,
            lcout => OPEN,
            ltout => \tok.n203_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__14836\,
            in1 => \N__19240\,
            in2 => \N__14827\,
            in3 => \N__31921\,
            lcout => OPEN,
            ltout => \tok.n212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6903_4_lut_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__31922\,
            in1 => \N__33414\,
            in2 => \N__14824\,
            in3 => \N__14821\,
            lcout => \tok.n6397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_224_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__36698\,
            in1 => \_gnd_net_\,
            in2 => \N__30857\,
            in3 => \_gnd_net_\,
            lcout => \tok.n5_adj_713\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \tok.n4774\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_99_add_2_3_lut_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32827\,
            in2 => \_gnd_net_\,
            in3 => \N__14815\,
            lcout => \tok.n238\,
            ltout => OPEN,
            carryin => \tok.n4774\,
            carryout => \tok.n4775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_99_add_2_4_lut_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31572\,
            in2 => \_gnd_net_\,
            in3 => \N__14812\,
            lcout => \tok.n237\,
            ltout => OPEN,
            carryin => \tok.n4775\,
            carryout => \tok.n4776\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_99_add_2_5_lut_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17515\,
            in2 => \N__34428\,
            in3 => \N__14809\,
            lcout => \tok.n236\,
            ltout => OPEN,
            carryin => \tok.n4776\,
            carryout => \tok.n4777\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_99_add_2_6_lut_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__30503\,
            in1 => \N__35612\,
            in2 => \_gnd_net_\,
            in3 => \N__14806\,
            lcout => \tok.n235\,
            ltout => OPEN,
            carryin => \tok.n4777\,
            carryout => \tok.n4778\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_99_add_2_7_lut_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__27560\,
            in1 => \N__36697\,
            in2 => \_gnd_net_\,
            in3 => \N__14803\,
            lcout => \tok.n234\,
            ltout => OPEN,
            carryin => \tok.n4778\,
            carryout => \tok.n4779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_99_add_2_8_lut_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__33633\,
            in1 => \N__17508\,
            in2 => \N__35057\,
            in3 => \N__14878\,
            lcout => \tok.n233\,
            ltout => OPEN,
            carryin => \tok.n4779\,
            carryout => \tok.n4780\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_99_add_2_9_lut_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__36528\,
            in1 => \N__17516\,
            in2 => \N__33797\,
            in3 => \N__14875\,
            lcout => \tok.n232\,
            ltout => OPEN,
            carryin => \tok.n4780\,
            carryout => \tok.n4781\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_99_add_2_10_lut_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__17507\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14872\,
            lcout => \tok.n214\,
            ltout => \tok.n214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6679_3_lut_4_lut_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__30716\,
            in1 => \N__34269\,
            in2 => \N__14869\,
            in3 => \N__23994\,
            lcout => \tok.n6358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_258_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__34268\,
            in1 => \N__32781\,
            in2 => \_gnd_net_\,
            in3 => \N__30715\,
            lcout => \tok.n786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_49_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35611\,
            in2 => \_gnd_net_\,
            in3 => \N__34267\,
            lcout => \tok.n289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_adj_117_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__35610\,
            in1 => \N__34917\,
            in2 => \N__36727\,
            in3 => \N__33711\,
            lcout => \tok.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6710_3_lut_4_lut_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__34270\,
            in1 => \N__30717\,
            in2 => \N__22250\,
            in3 => \N__20740\,
            lcout => \tok.n6402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i14_1_lut_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32210\,
            lcout => \tok.n312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_100_i15_2_lut_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__29621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20758\,
            lcout => \tok.n225\,
            ltout => \tok.n225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i312_4_lut_adj_50_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__14941\,
            in1 => \N__32785\,
            in2 => \N__14929\,
            in3 => \N__30721\,
            lcout => OPEN,
            ltout => \tok.n203_adj_664_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_51_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__31538\,
            in1 => \N__19218\,
            in2 => \N__14926\,
            in3 => \N__14923\,
            lcout => \tok.n212_adj_665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_100_i16_2_lut_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__20759\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23995\,
            lcout => \tok.n224\,
            ltout => \tok.n224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i312_4_lut_adj_73_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__30720\,
            in1 => \N__14911\,
            in2 => \N__14899\,
            in3 => \N__32786\,
            lcout => \tok.n203_adj_688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6689_3_lut_4_lut_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__20760\,
            in1 => \N__34397\,
            in2 => \N__30974\,
            in3 => \N__29622\,
            lcout => OPEN,
            ltout => \tok.n6373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i300_4_lut_adj_52_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20670\,
            in1 => \N__32281\,
            in2 => \N__14890\,
            in3 => \N__35722\,
            lcout => OPEN,
            ltout => \tok.n206_adj_666_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6890_4_lut_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__31547\,
            in1 => \N__33371\,
            in2 => \N__14887\,
            in3 => \N__14884\,
            lcout => \tok.n6368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_294_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__36946\,
            in1 => \N__14974\,
            in2 => \N__17548\,
            in3 => \N__34004\,
            lcout => OPEN,
            ltout => \tok.n281_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_300_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101000"
        )
    port map (
            in0 => \N__35272\,
            in1 => \N__14980\,
            in2 => \N__15001\,
            in3 => \N__30510\,
            lcout => OPEN,
            ltout => \tok.n236_adj_864_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_306_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__30729\,
            in1 => \N__14992\,
            in2 => \N__14998\,
            in3 => \N__31546\,
            lcout => \tok.n5_adj_871\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2624_4_lut_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36051\,
            in1 => \N__30509\,
            in2 => \N__35444\,
            in3 => \N__34275\,
            lcout => OPEN,
            ltout => \tok.n2648_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i360_4_lut_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100100010"
        )
    port map (
            in0 => \N__14986\,
            in1 => \N__34003\,
            in2 => \N__14995\,
            in3 => \N__32789\,
            lcout => \tok.n226_adj_865\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6994_3_lut_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35268\,
            in1 => \N__36945\,
            in2 => \_gnd_net_\,
            in3 => \N__30727\,
            lcout => \tok.n6334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__34274\,
            in1 => \N__31545\,
            in2 => \N__33135\,
            in3 => \N__36052\,
            lcout => \tok.n4_adj_762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6661_4_lut_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__36050\,
            in1 => \N__34273\,
            in2 => \_gnd_net_\,
            in3 => \N__30728\,
            lcout => \tok.n6316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i1_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14968\,
            lcout => tx_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38485\,
            ce => \N__27163\,
            sr => \N__37566\
        );

    \tok.A_stk.tail_i0_i65_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18448\,
            in1 => \N__15078\,
            in2 => \_gnd_net_\,
            in3 => \N__15070\,
            lcout => \tok.A_stk.tail_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38434\,
            ce => \N__17955\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i49_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15088\,
            in1 => \N__15060\,
            in2 => \_gnd_net_\,
            in3 => \N__18447\,
            lcout => tail_49,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38434\,
            ce => \N__17955\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i81_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18449\,
            in1 => \N__16389\,
            in2 => \_gnd_net_\,
            in3 => \N__15087\,
            lcout => tail_81,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38434\,
            ce => \N__17955\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i33_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15079\,
            in1 => \N__15048\,
            in2 => \_gnd_net_\,
            in3 => \N__18446\,
            lcout => \tok.A_stk.tail_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38434\,
            ce => \N__17955\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i97_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18450\,
            in1 => \N__16378\,
            in2 => \_gnd_net_\,
            in3 => \N__15069\,
            lcout => tail_97,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38434\,
            ce => \N__17955\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i17_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15040\,
            in1 => \N__15061\,
            in2 => \_gnd_net_\,
            in3 => \N__18444\,
            lcout => tail_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38434\,
            ce => \N__17955\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i1_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18445\,
            in1 => \_gnd_net_\,
            in2 => \N__15052\,
            in3 => \N__23496\,
            lcout => \tok.A_stk.tail_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38434\,
            ce => \N__17955\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i1_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15039\,
            in1 => \N__18585\,
            in2 => \_gnd_net_\,
            in3 => \N__27562\,
            lcout => \S_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38434\,
            ce => \N__17955\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i108_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16350\,
            in1 => \N__15258\,
            in2 => \_gnd_net_\,
            in3 => \N__18383\,
            lcout => tail_108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38438\,
            ce => \N__17925\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i86_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18389\,
            in1 => \N__15031\,
            in2 => \_gnd_net_\,
            in3 => \N__15144\,
            lcout => \tok.A_stk.tail_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38438\,
            ce => \N__17925\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i70_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15135\,
            in1 => \N__15015\,
            in2 => \_gnd_net_\,
            in3 => \N__18388\,
            lcout => \tok.A_stk.tail_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38438\,
            ce => \N__17925\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i54_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18386\,
            in1 => \N__15145\,
            in2 => \_gnd_net_\,
            in3 => \N__15126\,
            lcout => \tok.A_stk.tail_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38438\,
            ce => \N__17925\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i38_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15136\,
            in1 => \N__15117\,
            in2 => \_gnd_net_\,
            in3 => \N__18385\,
            lcout => \tok.A_stk.tail_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38438\,
            ce => \N__17925\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i22_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18384\,
            in1 => \N__15127\,
            in2 => \_gnd_net_\,
            in3 => \N__15225\,
            lcout => \tok.A_stk.tail_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38438\,
            ce => \N__17925\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i6_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15118\,
            in1 => \N__18387\,
            in2 => \_gnd_net_\,
            in3 => \N__25937\,
            lcout => \tok.A_stk.tail_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38438\,
            ce => \N__17925\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i92_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18390\,
            in1 => \N__16365\,
            in2 => \_gnd_net_\,
            in3 => \N__15237\,
            lcout => \tok.A_stk.tail_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38438\,
            ce => \N__17925\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i12_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18439\,
            in1 => \N__15106\,
            in2 => \_gnd_net_\,
            in3 => \N__20226\,
            lcout => \tok.A_stk.tail_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38443\,
            ce => \N__17927\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i28_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15214\,
            in1 => \N__15097\,
            in2 => \_gnd_net_\,
            in3 => \N__18440\,
            lcout => \tok.A_stk.tail_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38443\,
            ce => \N__17927\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i44_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18441\,
            in1 => \N__15105\,
            in2 => \_gnd_net_\,
            in3 => \N__15247\,
            lcout => \tok.A_stk.tail_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38443\,
            ce => \N__17927\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i60_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15238\,
            in1 => \N__15096\,
            in2 => \_gnd_net_\,
            in3 => \N__18442\,
            lcout => \tok.A_stk.tail_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38443\,
            ce => \N__17927\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i76_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18443\,
            in1 => \N__15259\,
            in2 => \_gnd_net_\,
            in3 => \N__15246\,
            lcout => \tok.A_stk.tail_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38443\,
            ce => \N__17927\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i6_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18565\,
            in1 => \N__15226\,
            in2 => \_gnd_net_\,
            in3 => \N__30073\,
            lcout => \tok.S_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38443\,
            ce => \N__17927\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i12_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15213\,
            in1 => \N__18564\,
            in2 => \_gnd_net_\,
            in3 => \N__27038\,
            lcout => \tok.S_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38443\,
            ce => \N__17927\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i10_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18563\,
            in1 => \N__15201\,
            in2 => \_gnd_net_\,
            in3 => \N__29628\,
            lcout => \tok.S_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38443\,
            ce => \N__17927\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i99_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18397\,
            in1 => \N__15273\,
            in2 => \_gnd_net_\,
            in3 => \N__15180\,
            lcout => tail_99,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38447\,
            ce => \N__17924\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i83_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15285\,
            in1 => \N__15171\,
            in2 => \_gnd_net_\,
            in3 => \N__18396\,
            lcout => \tok.A_stk.tail_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38447\,
            ce => \N__17924\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i67_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18395\,
            in1 => \N__15162\,
            in2 => \_gnd_net_\,
            in3 => \N__15181\,
            lcout => \tok.A_stk.tail_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38447\,
            ce => \N__17924\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i51_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15153\,
            in1 => \N__15172\,
            in2 => \_gnd_net_\,
            in3 => \N__18394\,
            lcout => \tok.A_stk.tail_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38447\,
            ce => \N__17924\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i35_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18392\,
            in1 => \N__15351\,
            in2 => \_gnd_net_\,
            in3 => \N__15163\,
            lcout => \tok.A_stk.tail_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38447\,
            ce => \N__17924\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i19_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__15154\,
            in1 => \_gnd_net_\,
            in2 => \N__15343\,
            in3 => \N__18391\,
            lcout => \tok.A_stk.tail_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38447\,
            ce => \N__17924\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i3_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18393\,
            in1 => \N__15352\,
            in2 => \_gnd_net_\,
            in3 => \N__23178\,
            lcout => \tok.A_stk.tail_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38447\,
            ce => \N__17924\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i3_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15339\,
            in1 => \N__18550\,
            in2 => \_gnd_net_\,
            in3 => \N__36513\,
            lcout => \tok.S_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38447\,
            ce => \N__17924\,
            sr => \_gnd_net_\
        );

    \tok.i6631_4_lut_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__34661\,
            in1 => \N__26512\,
            in2 => \N__18610\,
            in3 => \N__31095\,
            lcout => \tok.n6252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_4_lut_adj_299_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33240\,
            in1 => \N__34660\,
            in2 => \N__36231\,
            in3 => \N__32111\,
            lcout => \tok.n4\,
            ltout => \tok.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6594_2_lut_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15331\,
            in3 => \N__31094\,
            lcout => \tok.n6273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2623_2_lut_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21768\,
            lcout => \tok.table_wr_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6993_4_lut_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010001"
        )
    port map (
            in0 => \N__21514\,
            in1 => \N__37042\,
            in2 => \N__15307\,
            in3 => \N__31096\,
            lcout => OPEN,
            ltout => \tok.n6253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6119_4_lut_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__15298\,
            in1 => \N__16552\,
            in2 => \N__15289\,
            in3 => \N__35199\,
            lcout => \tok.n6203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i115_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__15286\,
            in1 => \N__17904\,
            in2 => \N__15274\,
            in3 => \N__18253\,
            lcout => tail_115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_90_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__25338\,
            in1 => \N__15661\,
            in2 => \N__33646\,
            in3 => \N__15787\,
            lcout => OPEN,
            ltout => \tok.n27_adj_704_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i2_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__15602\,
            in1 => \N__16770\,
            in2 => \N__15649\,
            in3 => \N__16668\,
            lcout => \tok.n38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38457\,
            ce => 'H',
            sr => \N__29216\
        );

    \tok.i314_4_lut_adj_266_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__27553\,
            in1 => \N__34461\,
            in2 => \N__15985\,
            in3 => \N__31907\,
            lcout => \tok.n161_adj_836\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_88_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__25343\,
            in1 => \N__15580\,
            in2 => \N__15796\,
            in3 => \N__27554\,
            lcout => \tok.n27_adj_703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_92_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__25339\,
            in1 => \N__36479\,
            in2 => \N__15568\,
            in3 => \N__15788\,
            lcout => OPEN,
            ltout => \tok.n27_adj_705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i3_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__15513\,
            in1 => \N__16771\,
            in2 => \N__15553\,
            in3 => \N__16669\,
            lcout => \tok.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38457\,
            ce => 'H',
            sr => \N__29216\
        );

    \tok.idx_i1_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__16666\,
            in1 => \N__15441\,
            in2 => \N__16782\,
            in3 => \N__15484\,
            lcout => \tok.n40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38457\,
            ce => 'H',
            sr => \N__29216\
        );

    \tok.idx_i5_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__15378\,
            in1 => \N__16667\,
            in2 => \N__16786\,
            in3 => \N__15880\,
            lcout => \tok.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38457\,
            ce => 'H',
            sr => \N__29216\
        );

    \tok.i314_4_lut_adj_40_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__30328\,
            in1 => \N__34481\,
            in2 => \N__16036\,
            in3 => \N__31908\,
            lcout => \tok.n161_adj_650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i6_1_lut_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30327\,
            lcout => \tok.n320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_96_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__30329\,
            in1 => \N__25329\,
            in2 => \N__15783\,
            in3 => \N__15889\,
            lcout => \tok.n27_adj_707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_98_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__30054\,
            in1 => \N__15771\,
            in2 => \N__25359\,
            in3 => \N__15874\,
            lcout => OPEN,
            ltout => \tok.n27_adj_708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i6_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__15840\,
            in1 => \N__16775\,
            in2 => \N__15865\,
            in3 => \N__16670\,
            lcout => \tok.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38462\,
            ce => 'H',
            sr => \N__29259\
        );

    \tok.search_clk_I_0_1_lut_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15767\,
            lcout => \tok.search_clk_N_137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.search_clk_359_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15772\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.search_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38462\,
            ce => 'H',
            sr => \N__29259\
        );

    \tok.i1_2_lut_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15766\,
            in2 => \_gnd_net_\,
            in3 => \N__15713\,
            lcout => \tok.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_375_i13_2_lut_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33802\,
            in2 => \_gnd_net_\,
            in3 => \N__35237\,
            lcout => \tok.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7002_4_lut_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__15955\,
            in1 => \N__30010\,
            in2 => \N__15967\,
            in3 => \N__30478\,
            lcout => \tok.n6670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15924\,
            in1 => \N__15963\,
            in2 => \N__15937\,
            in3 => \N__15954\,
            lcout => \tok.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_31_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__27524\,
            in1 => \N__15933\,
            in2 => \N__27387\,
            in3 => \N__15925\,
            lcout => \tok.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_281_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23548\,
            in1 => \N__27353\,
            in2 => \N__23843\,
            in3 => \N__27523\,
            lcout => \tok.n18_adj_850\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i317_4_lut_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111000000"
        )
    port map (
            in0 => \N__27357\,
            in1 => \N__36841\,
            in2 => \N__23844\,
            in3 => \N__31041\,
            lcout => \tok.n177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6817_4_lut_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__16006\,
            in1 => \N__23616\,
            in2 => \N__32075\,
            in3 => \N__16813\,
            lcout => OPEN,
            ltout => \tok.n6575_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i303_4_lut_adj_169_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__35238\,
            in1 => \N__25892\,
            in2 => \N__15904\,
            in3 => \N__15901\,
            lcout => \tok.n252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_2_lut_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18828\,
            in2 => \N__30508\,
            in3 => \N__31671\,
            lcout => \tok.n2579\,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \tok.n4797\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_3_lut_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__31672\,
            in1 => \N__27552\,
            in2 => \N__23546\,
            in3 => \N__15895\,
            lcout => \tok.n2635\,
            ltout => OPEN,
            carryin => \tok.n4797\,
            carryout => \tok.n4798\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_4_lut_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34460\,
            in1 => \N__33597\,
            in2 => \N__20095\,
            in3 => \N__15892\,
            lcout => \tok.n6615\,
            ltout => OPEN,
            carryin => \tok.n4798\,
            carryout => \tok.n4799\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_5_lut_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23210\,
            in2 => \N__36541\,
            in3 => \N__16009\,
            lcout => \tok.n288\,
            ltout => OPEN,
            carryin => \tok.n4799\,
            carryout => \tok.n4800\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_6_lut_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__32853\,
            in1 => \N__27386\,
            in2 => \N__23839\,
            in3 => \N__16000\,
            lcout => \tok.n6556\,
            ltout => OPEN,
            carryin => \tok.n4800\,
            carryout => \tok.n4801\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_7_lut_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__32877\,
            in1 => \N__30319\,
            in2 => \N__22027\,
            in3 => \N__15997\,
            lcout => \tok.n6514\,
            ltout => OPEN,
            carryin => \tok.n4801\,
            carryout => \tok.n4802\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_8_lut_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__32852\,
            in1 => \N__30042\,
            in2 => \N__25971\,
            in3 => \N__15994\,
            lcout => \tok.n6490\,
            ltout => OPEN,
            carryin => \tok.n4802\,
            carryout => \tok.n4803\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_8_THRU_CRY_0_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17517\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \tok.n4803\,
            carryout => \tok.n4803_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_9_lut_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__33093\,
            in1 => \N__37443\,
            in2 => \N__28330\,
            in3 => \N__15991\,
            lcout => \tok.n6466\,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \tok.n4804\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_10_lut_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16116\,
            in1 => \N__22233\,
            in2 => \N__17261\,
            in3 => \N__15988\,
            lcout => \tok.n6452\,
            ltout => OPEN,
            carryin => \tok.n4804\,
            carryout => \tok.n4805\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_11_lut_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16113\,
            in1 => \N__26775\,
            in2 => \N__21772\,
            in3 => \N__15973\,
            lcout => \tok.n6437\,
            ltout => OPEN,
            carryin => \tok.n4805\,
            carryout => \tok.n4806\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_12_lut_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16117\,
            in1 => \N__29577\,
            in2 => \N__20173\,
            in3 => \N__15970\,
            lcout => \tok.n6421\,
            ltout => OPEN,
            carryin => \tok.n4806\,
            carryout => \tok.n4807\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_13_lut_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16115\,
            in1 => \N__23992\,
            in2 => \N__19503\,
            in3 => \N__16042\,
            lcout => \tok.n6406\,
            ltout => OPEN,
            carryin => \tok.n4807\,
            carryout => \tok.n4808\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_14_lut_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16118\,
            in1 => \N__27036\,
            in2 => \N__20258\,
            in3 => \N__16039\,
            lcout => \tok.n6392\,
            ltout => OPEN,
            carryin => \tok.n4808\,
            carryout => \tok.n4809\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_15_lut_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16114\,
            in1 => \N__32200\,
            in2 => \N__17320\,
            in3 => \N__16024\,
            lcout => \tok.n6377\,
            ltout => OPEN,
            carryin => \tok.n4809\,
            carryout => \tok.n4810\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_15_THRU_CRY_0_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17485\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \tok.n4810\,
            carryout => \tok.n4810_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_16_lut_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__16119\,
            in1 => \N__32368\,
            in2 => \N__19336\,
            in3 => \N__16021\,
            lcout => \tok.n6362\,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \tok.n4811\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_103_17_lut_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__18963\,
            in1 => \N__16120\,
            in2 => \N__24199\,
            in3 => \N__16018\,
            lcout => \tok.n6339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_adj_53_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__31470\,
            in1 => \N__16015\,
            in2 => \N__30066\,
            in3 => \N__34266\,
            lcout => \tok.n161_adj_667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_4_lut_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__34265\,
            in1 => \N__35715\,
            in2 => \N__36980\,
            in3 => \N__32695\,
            lcout => \tok.n260_adj_717\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_284_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__30043\,
            in1 => \N__18835\,
            in2 => \N__25984\,
            in3 => \N__30531\,
            lcout => \tok.n17_adj_853\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_1_lut_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32694\,
            lcout => \tok.n21_adj_660\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34264\,
            lcout => \tok.n4_adj_635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i402_1_lut_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31468\,
            lcout => \tok.n83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_248_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__20341\,
            in1 => \N__24288\,
            in2 => \N__17266\,
            in3 => \N__17155\,
            lcout => \tok.n248_adj_827\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i299_4_lut_adj_267_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__35716\,
            in1 => \N__16087\,
            in2 => \N__17119\,
            in3 => \N__32779\,
            lcout => OPEN,
            ltout => \tok.n197_adj_837_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_268_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__20342\,
            in1 => \N__24289\,
            in2 => \N__16075\,
            in3 => \N__21761\,
            lcout => \tok.n248_adj_838\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6699_4_lut_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23731\,
            in1 => \N__20396\,
            in2 => \N__35874\,
            in3 => \N__16900\,
            lcout => OPEN,
            ltout => \tok.n6386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i299_4_lut_adj_42_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32780\,
            in1 => \N__16060\,
            in2 => \N__16048\,
            in3 => \N__35721\,
            lcout => OPEN,
            ltout => \tok.n197_adj_652_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_43_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__24290\,
            in1 => \N__20343\,
            in2 => \N__16045\,
            in3 => \N__17319\,
            lcout => \tok.n248_adj_653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6706_4_lut_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011100000"
        )
    port map (
            in0 => \N__17068\,
            in1 => \N__35717\,
            in2 => \N__20412\,
            in3 => \N__23730\,
            lcout => \tok.n6356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i335_rep_143_2_lut_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32778\,
            in2 => \_gnd_net_\,
            in3 => \N__30714\,
            lcout => \tok.n7269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_100_i12_2_lut_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__20785\,
            in1 => \N__37445\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n228\,
            ltout => \tok.n228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i312_4_lut_adj_320_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__30719\,
            in1 => \N__16180\,
            in2 => \N__16168\,
            in3 => \N__32787\,
            lcout => OPEN,
            ltout => \tok.n203_adj_879_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_321_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__31743\,
            in1 => \N__19214\,
            in2 => \N__16165\,
            in3 => \N__16162\,
            lcout => OPEN,
            ltout => \tok.n212_adj_880_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6911_4_lut_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__31548\,
            in1 => \N__33490\,
            in2 => \N__16156\,
            in3 => \N__16126\,
            lcout => \tok.n6412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6719_3_lut_4_lut_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__34271\,
            in1 => \N__30718\,
            in2 => \N__20792\,
            in3 => \N__37444\,
            lcout => \tok.n6417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_adj_76_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__31549\,
            in1 => \N__16153\,
            in2 => \N__37469\,
            in3 => \N__34272\,
            lcout => OPEN,
            ltout => \tok.n161_adj_692_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i299_4_lut_adj_77_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__32788\,
            in1 => \N__36142\,
            in2 => \N__16144\,
            in3 => \N__16141\,
            lcout => \tok.n197_adj_693\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i300_4_lut_adj_322_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__20690\,
            in1 => \N__20610\,
            in2 => \N__36283\,
            in3 => \N__16132\,
            lcout => \tok.n206_adj_881\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2579_2_lut_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33936\,
            in2 => \_gnd_net_\,
            in3 => \N__36548\,
            lcout => \tok.n2602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_327_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__30072\,
            in1 => \N__36852\,
            in2 => \N__26226\,
            in3 => \N__16267\,
            lcout => \tok.n242_adj_885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i103_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16261\,
            in1 => \N__16227\,
            in2 => \_gnd_net_\,
            in3 => \N__18451\,
            lcout => tail_103,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38439\,
            ce => \N__17947\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i87_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18457\,
            in1 => \N__16239\,
            in2 => \_gnd_net_\,
            in3 => \N__16218\,
            lcout => \tok.A_stk.tail_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38439\,
            ce => \N__17947\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i71_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16209\,
            in1 => \N__16228\,
            in2 => \_gnd_net_\,
            in3 => \N__18455\,
            lcout => \tok.A_stk.tail_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38439\,
            ce => \N__17947\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i55_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18454\,
            in1 => \N__16219\,
            in2 => \_gnd_net_\,
            in3 => \N__16200\,
            lcout => \tok.A_stk.tail_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38439\,
            ce => \N__17947\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i39_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16210\,
            in1 => \N__16191\,
            in2 => \_gnd_net_\,
            in3 => \N__18453\,
            lcout => \tok.A_stk.tail_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38439\,
            ce => \N__17947\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i23_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__18452\,
            in1 => \_gnd_net_\,
            in2 => \N__16408\,
            in3 => \N__16201\,
            lcout => \tok.A_stk.tail_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38439\,
            ce => \N__17947\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i7_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16192\,
            in1 => \N__18456\,
            in2 => \_gnd_net_\,
            in3 => \N__28297\,
            lcout => \tok.A_stk.tail_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38439\,
            ce => \N__17947\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i7_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16404\,
            in1 => \N__18562\,
            in2 => \_gnd_net_\,
            in3 => \N__37477\,
            lcout => \tok.S_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38439\,
            ce => \N__17947\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i113_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__18373\,
            in1 => \N__16377\,
            in2 => \N__16396\,
            in3 => \N__17902\,
            lcout => tail_113,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38444\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i124_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__17903\,
            in1 => \N__16366\,
            in2 => \N__16354\,
            in3 => \N__18374\,
            lcout => tail_124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38444\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.S_15__I_0_i4_3_lut_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23218\,
            in1 => \N__22646\,
            in2 => \_gnd_net_\,
            in3 => \N__28476\,
            lcout => \tok.table_wr_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1379_3_lut_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28475\,
            in1 => \N__24986\,
            in2 => \_gnd_net_\,
            in3 => \N__23495\,
            lcout => table_wr_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1464_3_lut_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27738\,
            in1 => \N__28477\,
            in2 => \_gnd_net_\,
            in3 => \N__25936\,
            lcout => \tok.table_wr_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1536_3_lut_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23851\,
            in1 => \N__21057\,
            in2 => \_gnd_net_\,
            in3 => \N__28478\,
            lcout => \tok.table_wr_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1572_3_lut_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28479\,
            in1 => \N__22487\,
            in2 => \_gnd_net_\,
            in3 => \N__20094\,
            lcout => \tok.table_wr_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6634_4_lut_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__22939\,
            in1 => \N__22875\,
            in2 => \N__27685\,
            in3 => \N__27736\,
            lcout => OPEN,
            ltout => \tok.ram.n6266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1456_4_lut_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__22807\,
            in1 => \N__27684\,
            in2 => \N__16459\,
            in3 => \N__31934\,
            lcout => OPEN,
            ltout => \tok.n1495_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_167_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__16417\,
            in1 => \N__35522\,
            in2 => \N__16456\,
            in3 => \N__31331\,
            lcout => \tok.n13_adj_766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i6_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16447\,
            in1 => \N__27707\,
            in2 => \_gnd_net_\,
            in3 => \N__19738\,
            lcout => tc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38448\,
            ce => 'H',
            sr => \N__29220\
        );

    \tok.i1_4_lut_adj_168_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__25809\,
            in1 => \N__16453\,
            in2 => \N__29725\,
            in3 => \N__27737\,
            lcout => n10_adj_907,
            ltout => \n10_adj_907_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_200_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27706\,
            in2 => \N__16441\,
            in3 => \N__19737\,
            lcout => \tok.tc_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_164_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__27680\,
            in1 => \N__33295\,
            in2 => \N__24060\,
            in3 => \N__31330\,
            lcout => OPEN,
            ltout => \tok.n83_adj_765_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6725_2_lut_3_lut_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__36306\,
            in1 => \_gnd_net_\,
            in2 => \N__16420\,
            in3 => \N__31933\,
            lcout => \tok.n6435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6614_4_lut_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__22945\,
            in1 => \N__21102\,
            in2 => \N__21167\,
            in3 => \N__22864\,
            lcout => OPEN,
            ltout => \tok.n6283_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i124_4_lut_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__22806\,
            in1 => \N__21101\,
            in2 => \N__16411\,
            in3 => \N__32022\,
            lcout => OPEN,
            ltout => \tok.n80_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i126_4_lut_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__16534\,
            in1 => \N__35504\,
            in2 => \N__16543\,
            in3 => \N__31252\,
            lcout => OPEN,
            ltout => \tok.n89_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_131_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__29718\,
            in1 => \N__25805\,
            in2 => \N__16540\,
            in3 => \N__21160\,
            lcout => n92_adj_897,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__16527\,
            in1 => \N__33137\,
            in2 => \N__21103\,
            in3 => \N__31251\,
            lcout => OPEN,
            ltout => \tok.n83_adj_734_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6637_2_lut_3_lut_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36183\,
            in2 => \N__16537\,
            in3 => \N__32021\,
            lcout => \tok.n6279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i358_4_lut_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__17421\,
            in1 => \N__33136\,
            in2 => \N__16528\,
            in3 => \N__31250\,
            lcout => \tok.n2696\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2618_2_lut_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28424\,
            in2 => \_gnd_net_\,
            in3 => \N__19333\,
            lcout => \tok.table_wr_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2583_2_lut_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__28448\,
            in1 => \N__19514\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.table_wr_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2542_2_lut_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28447\,
            in2 => \_gnd_net_\,
            in3 => \N__20238\,
            lcout => \tok.table_wr_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_292_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110011"
        )
    port map (
            in0 => \N__17422\,
            in1 => \N__16465\,
            in2 => \N__19252\,
            in3 => \N__32109\,
            lcout => \tok.n268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.stall_I_0_369_i11_2_lut_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31093\,
            in2 => \_gnd_net_\,
            in3 => \N__33236\,
            lcout => \tok.n9_adj_651\,
            ltout => \tok.n9_adj_651_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_4_lut_adj_293_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__30142\,
            in1 => \N__34643\,
            in2 => \N__16594\,
            in3 => \N__32110\,
            lcout => n15,
            ltout => \n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_69_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__16591\,
            in1 => \N__21363\,
            in2 => \N__16582\,
            in3 => \N__19609\,
            lcout => OPEN,
            ltout => \tok.n6_adj_687_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_71_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__30144\,
            in1 => \N__27923\,
            in2 => \N__16579\,
            in3 => \N__16575\,
            lcout => \tok.n2702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_4_lut_adj_275_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__32108\,
            in1 => \N__26129\,
            in2 => \N__34780\,
            in3 => \N__30143\,
            lcout => \tok.n891\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_255_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101111"
        )
    port map (
            in0 => \N__29448\,
            in1 => \_gnd_net_\,
            in2 => \N__37241\,
            in3 => \N__37203\,
            lcout => \tok.uart_stall\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_257_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__37202\,
            in1 => \N__37230\,
            in2 => \_gnd_net_\,
            in3 => \N__29447\,
            lcout => \tok.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_33_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__16728\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16714\,
            lcout => \tok.n6170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_4_lut_adj_312_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__37234\,
            in1 => \N__29449\,
            in2 => \N__37207\,
            in3 => \N__16727\,
            lcout => \tok.n796\,
            ltout => \tok.n796_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_28_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011011100"
        )
    port map (
            in0 => \N__25354\,
            in1 => \N__16715\,
            in2 => \N__16546\,
            in3 => \N__16794\,
            lcout => \stall_\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.stall_361_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001100"
        )
    port map (
            in0 => \N__16795\,
            in1 => \N__16769\,
            in2 => \N__25358\,
            in3 => \N__16717\,
            lcout => \tok.stall\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38463\,
            ce => 'H',
            sr => \N__29242\
        );

    \tok.i36_4_lut_4_lut_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__16729\,
            in1 => \N__16716\,
            in2 => \N__25374\,
            in3 => \N__16699\,
            lcout => OPEN,
            ltout => \tok.n31_adj_637_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_29_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__25325\,
            in1 => \N__16693\,
            in2 => \N__16687\,
            in3 => \N__16684\,
            lcout => \tok.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_276_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__21987\,
            in1 => \N__30324\,
            in2 => \N__23215\,
            in3 => \N__36454\,
            lcout => \tok.n20_adj_845\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_154_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__36457\,
            in1 => \N__25153\,
            in2 => \N__19870\,
            in3 => \N__28993\,
            lcout => OPEN,
            ltout => \tok.n221_adj_753_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i4_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__25499\,
            in1 => \N__18658\,
            in2 => \N__16636\,
            in3 => \N__23209\,
            lcout => \tok.A_low_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38469\,
            ce => \N__25640\,
            sr => \N__29260\
        );

    \tok.i189_1_lut_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36453\,
            lcout => \tok.n127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__16633\,
            in1 => \N__30325\,
            in2 => \N__16615\,
            in3 => \N__36455\,
            lcout => OPEN,
            ltout => \tok.n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_35_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111110"
        )
    port map (
            in0 => \N__16885\,
            in1 => \N__16840\,
            in2 => \N__16867\,
            in3 => \N__22232\,
            lcout => \tok.n26_adj_645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_185_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32190\,
            in1 => \N__30326\,
            in2 => \N__22249\,
            in3 => \N__36456\,
            lcout => \tok.n26_adj_781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.key_rd_15__I_0_401_i14_2_lut_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16855\,
            in2 => \_gnd_net_\,
            in3 => \N__32189\,
            lcout => \tok.n14_adj_644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_2_lut_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18865\,
            in2 => \N__18832\,
            in3 => \N__16834\,
            lcout => \tok.n308\,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \tok.n4782\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_3_lut_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23374\,
            in2 => \N__23547\,
            in3 => \N__16831\,
            lcout => \tok.n307\,
            ltout => OPEN,
            carryin => \tok.n4782\,
            carryout => \tok.n4783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_4_lut_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__31898\,
            in1 => \N__20087\,
            in2 => \N__18874\,
            in3 => \N__16828\,
            lcout => \tok.n6616\,
            ltout => OPEN,
            carryin => \tok.n4783\,
            carryout => \tok.n4784\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_5_lut_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__33022\,
            in1 => \N__23211\,
            in2 => \N__16825\,
            in3 => \N__16816\,
            lcout => \tok.n2613\,
            ltout => OPEN,
            carryin => \tok.n4784\,
            carryout => \tok.n4785\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_6_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17012\,
            in1 => \N__20587\,
            in2 => \N__23852\,
            in3 => \N__16807\,
            lcout => \tok.n6557\,
            ltout => OPEN,
            carryin => \tok.n4785\,
            carryout => \tok.n4786\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_7_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17014\,
            in1 => \N__16804\,
            in2 => \N__22030\,
            in3 => \N__16798\,
            lcout => \tok.n6515\,
            ltout => OPEN,
            carryin => \tok.n4786\,
            carryout => \tok.n4787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_8_lut_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17011\,
            in1 => \N__18637\,
            in2 => \N__25988\,
            in3 => \N__17017\,
            lcout => \tok.n6491\,
            ltout => OPEN,
            carryin => \tok.n4787\,
            carryout => \tok.n4788\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_8_THRU_CRY_0_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__17509\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \tok.n4788\,
            carryout => \tok.n4788_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_9_lut_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17013\,
            in1 => \N__28328\,
            in2 => \N__16981\,
            in3 => \N__16969\,
            lcout => \tok.n6467\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \tok.n4789\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_10_lut_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20500\,
            in2 => \N__17265\,
            in3 => \N__16966\,
            lcout => \tok.n300\,
            ltout => OPEN,
            carryin => \tok.n4789\,
            carryout => \tok.n4790\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_11_lut_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21773\,
            in2 => \N__24019\,
            in3 => \N__16963\,
            lcout => \tok.n299\,
            ltout => OPEN,
            carryin => \tok.n4790\,
            carryout => \tok.n4791\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_12_lut_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20180\,
            in2 => \N__16960\,
            in3 => \N__16948\,
            lcout => \tok.n298\,
            ltout => OPEN,
            carryin => \tok.n4791\,
            carryout => \tok.n4792\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_13_lut_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19504\,
            in2 => \N__20614\,
            in3 => \N__16945\,
            lcout => \tok.n297\,
            ltout => OPEN,
            carryin => \tok.n4792\,
            carryout => \tok.n4793\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_14_lut_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20248\,
            in2 => \N__16942\,
            in3 => \N__16930\,
            lcout => \tok.n296\,
            ltout => OPEN,
            carryin => \tok.n4793\,
            carryout => \tok.n4794\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_15_lut_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17318\,
            in2 => \N__16926\,
            in3 => \N__16888\,
            lcout => \tok.n295\,
            ltout => OPEN,
            carryin => \tok.n4794\,
            carryout => \tok.n4795\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_16_lut_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19321\,
            in2 => \N__32274\,
            in3 => \N__17074\,
            lcout => \tok.n294\,
            ltout => OPEN,
            carryin => \tok.n4795\,
            carryout => \tok.n4796\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_104_add_2_17_lut_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18955\,
            in1 => \N__17053\,
            in2 => \_gnd_net_\,
            in3 => \N__17071\,
            lcout => \tok.n293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6717_4_lut_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011100000"
        )
    port map (
            in0 => \N__17059\,
            in1 => \N__36010\,
            in2 => \N__20406\,
            in3 => \N__23720\,
            lcout => \tok.n6415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i16_1_lut_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24143\,
            lcout => \tok.n310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_adj_246_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__31912\,
            in1 => \N__17047\,
            in2 => \N__34711\,
            in3 => \N__30487\,
            lcout => \tok.n161_adj_825\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i356_4_lut_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101000100"
        )
    port map (
            in0 => \N__17041\,
            in1 => \N__34551\,
            in2 => \N__37747\,
            in3 => \N__31913\,
            lcout => \tok.n208_adj_857\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__31915\,
            in1 => \N__17035\,
            in2 => \N__34712\,
            in3 => \N__27370\,
            lcout => \tok.n161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_adj_305_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010100000"
        )
    port map (
            in0 => \N__17029\,
            in1 => \N__33582\,
            in2 => \N__34713\,
            in3 => \N__31914\,
            lcout => \tok.n161_adj_870\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6746_4_lut_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011100000"
        )
    port map (
            in0 => \N__17023\,
            in1 => \N__36009\,
            in2 => \N__20405\,
            in3 => \N__23719\,
            lcout => \tok.n6460\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i299_4_lut_adj_247_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__17170\,
            in1 => \N__35831\,
            in2 => \N__17164\,
            in3 => \N__33234\,
            lcout => \tok.n197_adj_826\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_103_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36780\,
            in1 => \N__31765\,
            in2 => \_gnd_net_\,
            in3 => \N__34528\,
            lcout => \tok.n4_adj_711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i15_4_lut_adj_285_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17149\,
            in1 => \N__17137\,
            in2 => \N__18886\,
            in3 => \N__17179\,
            lcout => \tok.n31\,
            ltout => \tok.n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6736_4_lut_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__35829\,
            in1 => \N__20400\,
            in2 => \N__17131\,
            in3 => \N__17128\,
            lcout => \tok.n6446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6667_4_lut_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000010000"
        )
    port map (
            in0 => \N__17110\,
            in1 => \N__35830\,
            in2 => \N__20416\,
            in3 => \N__23726\,
            lcout => \tok.n6328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6688_4_lut_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23727\,
            in1 => \N__20404\,
            in2 => \N__36031\,
            in3 => \N__17101\,
            lcout => OPEN,
            ltout => \tok.n6371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i299_4_lut_adj_54_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__17092\,
            in1 => \N__35835\,
            in2 => \N__17086\,
            in3 => \N__33235\,
            lcout => \tok.n197_adj_668\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_172_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__35828\,
            in1 => \_gnd_net_\,
            in2 => \N__36935\,
            in3 => \N__34527\,
            lcout => \tok.n4_adj_680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_45_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__37083\,
            in1 => \N__35206\,
            in2 => \N__17083\,
            in3 => \N__17326\,
            lcout => OPEN,
            ltout => \tok.n200_adj_655_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_48_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__26611\,
            in1 => \N__32188\,
            in2 => \N__17350\,
            in3 => \N__33935\,
            lcout => OPEN,
            ltout => \tok.n6_adj_658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i14_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__25517\,
            in1 => \N__24484\,
            in2 => \N__17347\,
            in3 => \N__17314\,
            lcout => \tok.n44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38489\,
            ce => \N__25650\,
            sr => \N__29269\
        );

    \tok.i2_4_lut_adj_254_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__22189\,
            in1 => \N__33934\,
            in2 => \N__26617\,
            in3 => \N__19396\,
            lcout => OPEN,
            ltout => \tok.n6_adj_832_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i9_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__25518\,
            in1 => \N__20824\,
            in2 => \N__17344\,
            in3 => \N__17251\,
            lcout => \tok.n49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38489\,
            ce => \N__25650\,
            sr => \N__29269\
        );

    \tok.i308_4_lut_adj_44_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__22188\,
            in1 => \N__37082\,
            in2 => \N__26222\,
            in3 => \N__17341\,
            lcout => \tok.n242_adj_654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_106_i14_2_lut_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32169\,
            in2 => \_gnd_net_\,
            in3 => \N__17313\,
            lcout => OPEN,
            ltout => \tok.n14_adj_844_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_282_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__17250\,
            in1 => \N__22167\,
            in2 => \N__17191\,
            in3 => \N__17188\,
            lcout => \tok.n26_adj_851\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6663_3_lut_4_lut_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34558\,
            in1 => \N__36030\,
            in2 => \N__30534\,
            in3 => \N__33100\,
            lcout => OPEN,
            ltout => \tok.n6324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i366_4_lut_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__30859\,
            in1 => \N__33431\,
            in2 => \N__17173\,
            in3 => \N__17414\,
            lcout => OPEN,
            ltout => \tok.n262_adj_858_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6669_4_lut_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__31916\,
            in1 => \N__33432\,
            in2 => \N__17563\,
            in3 => \N__17560\,
            lcout => \tok.n6315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => \CONSTANT_ONE_NET_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_99_add_2_2_lut_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17425\,
            in3 => \N__30858\,
            lcout => \tok.n239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i3_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30524\,
            in1 => \N__20863\,
            in2 => \_gnd_net_\,
            in3 => \N__37540\,
            lcout => sender_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38494\,
            ce => \N__27171\,
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_80_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__29618\,
            in1 => \N__37077\,
            in2 => \N__26227\,
            in3 => \N__17380\,
            lcout => \tok.n242_adj_695\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_79_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__24328\,
            in1 => \N__20344\,
            in2 => \N__18973\,
            in3 => \N__17368\,
            lcout => OPEN,
            ltout => \tok.n248_adj_694_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_81_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__35266\,
            in1 => \N__37078\,
            in2 => \N__17362\,
            in3 => \N__17359\,
            lcout => OPEN,
            ltout => \tok.n200_adj_696_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_84_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__33994\,
            in1 => \N__26609\,
            in2 => \N__17353\,
            in3 => \N__24133\,
            lcout => OPEN,
            ltout => \tok.n6_adj_699_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i16_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__25519\,
            in1 => \N__18972\,
            in2 => \N__17584\,
            in3 => \N__20908\,
            lcout => \tok.n42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38499\,
            ce => \N__25642\,
            sr => \N__29272\
        );

    \tok.i6872_2_lut_3_lut_4_lut_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__37076\,
            in1 => \N__24426\,
            in2 => \N__34080\,
            in3 => \N__29617\,
            lcout => \tok.n6367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6865_2_lut_3_lut_4_lut_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__27362\,
            in1 => \N__33987\,
            in2 => \N__24453\,
            in3 => \N__37075\,
            lcout => \tok.n6456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6869_2_lut_3_lut_4_lut_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__37074\,
            in1 => \N__24425\,
            in2 => \N__34079\,
            in3 => \N__37470\,
            lcout => \tok.n6411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_404_2_lut_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21124\,
            in2 => \_gnd_net_\,
            in3 => \N__17581\,
            lcout => tc_plus_1_0,
            ltout => OPEN,
            carryin => \bfn_6_2_0_\,
            carryout => \tok.n4812\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_404_3_lut_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24955\,
            in2 => \_gnd_net_\,
            in3 => \N__17578\,
            lcout => tc_plus_1_1,
            ltout => OPEN,
            carryin => \tok.n4812\,
            carryout => \tok.n4813\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_404_4_lut_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22456\,
            in2 => \_gnd_net_\,
            in3 => \N__17575\,
            lcout => \tok.tc_plus_1_2\,
            ltout => OPEN,
            carryin => \tok.n4813\,
            carryout => \tok.n4814\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_404_5_lut_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22606\,
            in2 => \_gnd_net_\,
            in3 => \N__17572\,
            lcout => \tok.tc_plus_1_3\,
            ltout => OPEN,
            carryin => \tok.n4814\,
            carryout => \tok.n4815\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_404_6_lut_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21028\,
            in2 => \_gnd_net_\,
            in3 => \N__17569\,
            lcout => \tok.tc_plus_1_4\,
            ltout => OPEN,
            carryin => \tok.n4815\,
            carryout => \tok.n4816\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_404_7_lut_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22306\,
            in2 => \_gnd_net_\,
            in3 => \N__17566\,
            lcout => \tok.tc_plus_1_5\,
            ltout => OPEN,
            carryin => \tok.n4816\,
            carryout => \tok.n4817\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_404_8_lut_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27711\,
            in3 => \N__17635\,
            lcout => \tok.tc_plus_1_6\,
            ltout => OPEN,
            carryin => \tok.n4817\,
            carryout => \tok.n4818\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_404_9_lut_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27977\,
            in2 => \_gnd_net_\,
            in3 => \N__17632\,
            lcout => \tok.tc_plus_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_162_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__31333\,
            in1 => \N__17602\,
            in2 => \N__17593\,
            in3 => \N__35502\,
            lcout => OPEN,
            ltout => \tok.n13_adj_760_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_163_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__29711\,
            in1 => \N__25813\,
            in2 => \N__17629\,
            in3 => \N__22334\,
            lcout => n10_adj_905,
            ltout => \n10_adj_905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_201_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19730\,
            in1 => \_gnd_net_\,
            in2 => \N__17626\,
            in3 => \N__22307\,
            lcout => \tok.tc_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6619_4_lut_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__22931\,
            in1 => \N__22333\,
            in2 => \N__22876\,
            in3 => \N__22287\,
            lcout => OPEN,
            ltout => \tok.ram.n6263_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1492_4_lut_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__22288\,
            in1 => \N__22801\,
            in2 => \N__17605\,
            in3 => \N__31938\,
            lcout => \tok.n1530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_160_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__33101\,
            in1 => \N__22286\,
            in2 => \N__19906\,
            in3 => \N__31332\,
            lcout => OPEN,
            ltout => \tok.n83_adj_759_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6973_2_lut_3_lut_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36324\,
            in2 => \N__17596\,
            in3 => \N__31937\,
            lcout => \tok.n6660\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i5_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22308\,
            in1 => \N__17695\,
            in2 => \_gnd_net_\,
            in3 => \N__19731\,
            lcout => tc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38452\,
            ce => 'H',
            sr => \N__29230\
        );

    \tok.i125_4_lut_adj_195_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__27854\,
            in1 => \N__33162\,
            in2 => \N__21681\,
            in3 => \N__31324\,
            lcout => OPEN,
            ltout => \tok.n83_adj_764_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6978_2_lut_3_lut_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36184\,
            in2 => \N__17689\,
            in3 => \N__32023\,
            lcout => \tok.n6662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6596_4_lut_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__28363\,
            in1 => \N__22944\,
            in2 => \N__27859\,
            in3 => \N__22863\,
            lcout => OPEN,
            ltout => \tok.ram.n6277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1600_4_lut_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__22802\,
            in1 => \N__27858\,
            in2 => \N__17686\,
            in3 => \N__32024\,
            lcout => \tok.n1635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_197_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__17647\,
            in1 => \N__29719\,
            in2 => \N__28373\,
            in3 => \N__25806\,
            lcout => n10,
            ltout => \n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27970\,
            in2 => \N__17683\,
            in3 => \N__19728\,
            lcout => \tok.tc_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_196_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__17662\,
            in1 => \N__35443\,
            in2 => \N__17656\,
            in3 => \N__31325\,
            lcout => \tok.n13_adj_790\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i7_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27979\,
            in1 => \N__17641\,
            in2 => \_gnd_net_\,
            in3 => \N__19729\,
            lcout => tc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38458\,
            ce => 'H',
            sr => \N__29180\
        );

    \tok.i1_2_lut_adj_236_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35394\,
            in2 => \_gnd_net_\,
            in3 => \N__37003\,
            lcout => \tok.n5_adj_715\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_78_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__37002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36179\,
            lcout => \tok.n5_adj_675\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6962_4_lut_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__33609\,
            in1 => \N__35395\,
            in2 => \N__36294\,
            in3 => \N__34704\,
            lcout => \tok.n6632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_98_i7_3_lut_4_lut_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000111"
        )
    port map (
            in0 => \N__37001\,
            in1 => \N__36178\,
            in2 => \N__35495\,
            in3 => \N__33608\,
            lcout => \tok.n206_adj_794\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6121_2_lut_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__29413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31110\,
            lcout => OPEN,
            ltout => \tok.n6205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_127_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__27133\,
            in1 => \N__18606\,
            in2 => \N__18592\,
            in3 => \N__26260\,
            lcout => \tok.n270\,
            ltout => \tok.n270_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i2_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__33610\,
            in1 => \_gnd_net_\,
            in2 => \N__18481\,
            in3 => \N__17967\,
            lcout => \tok.S_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38464\,
            ce => \N__17956\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i2_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18478\,
            in1 => \N__18254\,
            in2 => \_gnd_net_\,
            in3 => \N__20076\,
            lcout => \tok.A_stk.tail_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38464\,
            ce => \N__17956\,
            sr => \_gnd_net_\
        );

    \tok.i339_4_lut_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__22984\,
            in1 => \N__21310\,
            in2 => \N__23458\,
            in3 => \N__36950\,
            lcout => OPEN,
            ltout => \tok.n283_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i347_4_lut_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__21394\,
            in1 => \N__26317\,
            in2 => \N__18664\,
            in3 => \N__35479\,
            lcout => OPEN,
            ltout => \tok.n223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_153_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__34083\,
            in1 => \N__36951\,
            in2 => \N__18661\,
            in3 => \N__18649\,
            lcout => \tok.n4_adj_752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6826_4_lut_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__20695\,
            in1 => \N__34082\,
            in2 => \N__36534\,
            in3 => \N__19951\,
            lcout => OPEN,
            ltout => \tok.n6586_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i340_4_lut_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011101"
        )
    port map (
            in0 => \N__23035\,
            in1 => \N__18643\,
            in2 => \N__18652\,
            in3 => \N__36185\,
            lcout => \tok.n226_adj_744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_146_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__21415\,
            in1 => \N__34081\,
            in2 => \N__19975\,
            in3 => \N__35478\,
            lcout => \tok.n254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i7_1_lut_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29931\,
            lcout => \tok.n319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6811_2_lut_3_lut_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__36948\,
            in1 => \N__30393\,
            in2 => \_gnd_net_\,
            in3 => \N__33945\,
            lcout => \tok.n6567\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i364_4_lut_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__35474\,
            in1 => \N__18628\,
            in2 => \N__19141\,
            in3 => \N__31222\,
            lcout => OPEN,
            ltout => \tok.n387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_296_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110010"
        )
    port map (
            in0 => \N__23020\,
            in1 => \N__18833\,
            in2 => \N__18616\,
            in3 => \N__33946\,
            lcout => OPEN,
            ltout => \tok.n254_adj_860_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_297_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__21916\,
            in1 => \N__34705\,
            in2 => \N__18613\,
            in3 => \N__31223\,
            lcout => \tok.n256_adj_862\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i178_1_lut_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30391\,
            lcout => \tok.n163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_303_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__30394\,
            in1 => \N__36949\,
            in2 => \N__19846\,
            in3 => \N__18859\,
            lcout => OPEN,
            ltout => \tok.n6_adj_868_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011011100000100"
        )
    port map (
            in0 => \N__18853\,
            in1 => \N__25482\,
            in2 => \N__18838\,
            in3 => \N__18834\,
            lcout => \tok.A_low_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38473\,
            ce => \N__25639\,
            sr => \N__29237\
        );

    \tok.i6804_2_lut_3_lut_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__30392\,
            in1 => \N__36947\,
            in2 => \_gnd_net_\,
            in3 => \N__31221\,
            lcout => \tok.n6532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i12_4_lut_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18705\,
            in1 => \N__18688\,
            in2 => \N__18733\,
            in3 => \N__18753\,
            lcout => \tok.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__23966\,
            in1 => \N__32356\,
            in2 => \N__18754\,
            in3 => \N__18729\,
            lcout => \tok.n23_adj_638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_4_lut_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__26773\,
            in1 => \N__24185\,
            in2 => \N__18706\,
            in3 => \N__18687\,
            lcout => \tok.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i12_4_lut_adj_182_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23967\,
            in1 => \N__24186\,
            in2 => \N__32373\,
            in3 => \N__26774\,
            lcout => OPEN,
            ltout => \tok.n28_adj_778_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i15_4_lut_adj_192_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18988\,
            in1 => \N__19063\,
            in2 => \N__18982\,
            in3 => \N__18979\,
            lcout => \tok.tc__7__N_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_191_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27358\,
            in1 => \N__27510\,
            in2 => \N__30053\,
            in3 => \N__30410\,
            lcout => \tok.n25_adj_788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_279_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__32355\,
            in1 => \N__19320\,
            in2 => \N__19487\,
            in3 => \N__23965\,
            lcout => \tok.n23_adj_848\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_4_lut_adj_277_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24184\,
            in1 => \N__26772\,
            in2 => \N__21777\,
            in3 => \N__18950\,
            lcout => \tok.n24_adj_846\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i3_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__25500\,
            in1 => \N__18907\,
            in2 => \N__20090\,
            in3 => \N__23413\,
            lcout => \tok.A_low_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38483\,
            ce => \N__25641\,
            sr => \N__29117\
        );

    \tok.i6983_4_lut_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__33564\,
            in1 => \N__36375\,
            in2 => \N__19627\,
            in3 => \N__19591\,
            lcout => \tok.n6634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_280_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__20249\,
            in1 => \N__20179\,
            in2 => \N__29562\,
            in3 => \N__26987\,
            lcout => OPEN,
            ltout => \tok.n21_adj_849_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i14_4_lut_adj_283_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18901\,
            in1 => \N__19069\,
            in2 => \N__18895\,
            in3 => \N__18892\,
            lcout => \tok.n30_adj_852\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i3_1_lut_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33561\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_278_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__28298\,
            in1 => \N__20077\,
            in2 => \N__37400\,
            in3 => \N__33562\,
            lcout => \tok.n22_adj_847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i11_4_lut_adj_186_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33563\,
            in1 => \N__37359\,
            in2 => \N__27012\,
            in3 => \N__29529\,
            lcout => \tok.n27_adj_782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6728_4_lut_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23728\,
            in1 => \N__20426\,
            in2 => \N__36213\,
            in3 => \N__19057\,
            lcout => OPEN,
            ltout => \tok.n6429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i299_4_lut_adj_307_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__19051\,
            in1 => \N__36015\,
            in2 => \N__19045\,
            in3 => \N__32960\,
            lcout => OPEN,
            ltout => \tok.n197_adj_872_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_308_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__20322\,
            in1 => \N__24333\,
            in2 => \N__19042\,
            in3 => \N__20190\,
            lcout => \tok.n248_adj_873\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6708_4_lut_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011100000"
        )
    port map (
            in0 => \N__19024\,
            in1 => \N__36014\,
            in2 => \N__20433\,
            in3 => \N__23729\,
            lcout => OPEN,
            ltout => \tok.n6400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i299_4_lut_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__36016\,
            in1 => \N__32958\,
            in2 => \N__19018\,
            in3 => \N__19015\,
            lcout => \tok.n197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_adj_323_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__34535\,
            in1 => \N__36509\,
            in2 => \N__19009\,
            in3 => \N__32020\,
            lcout => OPEN,
            ltout => \tok.n161_adj_882_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i299_4_lut_adj_324_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__36018\,
            in1 => \N__18997\,
            in2 => \N__18991\,
            in3 => \N__32959\,
            lcout => \tok.n197_adj_883\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i363_4_lut_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__19159\,
            in1 => \N__36017\,
            in2 => \N__19150\,
            in3 => \N__32961\,
            lcout => \tok.n250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_adj_237_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001001000"
        )
    port map (
            in0 => \N__36747\,
            in1 => \N__32018\,
            in2 => \N__30499\,
            in3 => \N__31049\,
            lcout => \tok.n190_adj_774\,
            ltout => \tok.n190_adj_774_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_adj_176_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__26383\,
            in1 => \N__19935\,
            in2 => \N__19129\,
            in3 => \N__36748\,
            lcout => \tok.n255_adj_775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_206_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36746\,
            in1 => \N__35723\,
            in2 => \_gnd_net_\,
            in3 => \N__31048\,
            lcout => \tok.n833\,
            ltout => \tok.n833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6800_4_lut_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__32019\,
            in1 => \N__19126\,
            in2 => \N__19114\,
            in3 => \N__19111\,
            lcout => OPEN,
            ltout => \tok.n6534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i303_4_lut_adj_187_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__25893\,
            in1 => \N__19075\,
            in2 => \N__19102\,
            in3 => \N__35300\,
            lcout => OPEN,
            ltout => \tok.n252_adj_783_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_189_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__35301\,
            in1 => \N__19081\,
            in2 => \N__19099\,
            in3 => \N__34536\,
            lcout => \tok.n4_adj_786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_184_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__26316\,
            in1 => \N__19096\,
            in2 => \N__19090\,
            in3 => \N__35724\,
            lcout => \tok.n258_adj_780\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i317_4_lut_adj_183_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000001010"
        )
    port map (
            in0 => \N__31050\,
            in1 => \N__22014\,
            in2 => \N__30312\,
            in3 => \N__36749\,
            lcout => \tok.n177_adj_779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_56_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__36978\,
            in1 => \N__26780\,
            in2 => \N__26217\,
            in3 => \N__19363\,
            lcout => \tok.n242_adj_670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_55_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__19354\,
            in1 => \N__20340\,
            in2 => \N__24317\,
            in3 => \N__19334\,
            lcout => OPEN,
            ltout => \tok.n248_adj_669_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_57_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__36979\,
            in1 => \N__35198\,
            in2 => \N__19348\,
            in3 => \N__19345\,
            lcout => OPEN,
            ltout => \tok.n200_adj_671_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_60_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__26587\,
            in1 => \N__33995\,
            in2 => \N__19339\,
            in3 => \N__32330\,
            lcout => OPEN,
            ltout => \tok.n6_adj_674_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i15_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__19335\,
            in1 => \N__25515\,
            in2 => \N__19270\,
            in3 => \N__20896\,
            lcout => \tok.n43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38495\,
            ce => \N__25644\,
            sr => \N__29262\
        );

    \tok.i312_4_lut_adj_244_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__32965\,
            in1 => \N__30907\,
            in2 => \N__19267\,
            in3 => \N__19389\,
            lcout => OPEN,
            ltout => \tok.n203_adj_822_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_319_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__19390\,
            in1 => \N__19245\,
            in2 => \N__19168\,
            in3 => \N__32064\,
            lcout => OPEN,
            ltout => \tok.n212_adj_824_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6928_4_lut_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__32065\,
            in1 => \N__33471\,
            in2 => \N__19165\,
            in3 => \N__20620\,
            lcout => OPEN,
            ltout => \tok.n6457_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_249_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__26207\,
            in1 => \N__36957\,
            in2 => \N__19162\,
            in3 => \N__36535\,
            lcout => OPEN,
            ltout => \tok.n242_adj_828_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_250_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__36958\,
            in1 => \N__19411\,
            in2 => \N__19399\,
            in3 => \N__35329\,
            lcout => \tok.n200_adj_829\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_32_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35264\,
            in2 => \_gnd_net_\,
            in3 => \N__36029\,
            lcout => \tok.n4_adj_640\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_100_i9_2_lut_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27374\,
            in2 => \_gnd_net_\,
            in3 => \N__20793\,
            lcout => \tok.n231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_2_lut_3_lut_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__30906\,
            in1 => \N__36956\,
            in2 => \_gnd_net_\,
            in3 => \N__32063\,
            lcout => \tok.n838\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_328_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__35465\,
            in1 => \N__36955\,
            in2 => \N__19423\,
            in3 => \N__19381\,
            lcout => OPEN,
            ltout => \tok.n200_adj_886_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_331_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__26610\,
            in1 => \N__33952\,
            in2 => \N__19372\,
            in3 => \N__23953\,
            lcout => OPEN,
            ltout => \tok.n6_adj_889_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i12_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__25516\,
            in1 => \N__22390\,
            in2 => \N__19369\,
            in3 => \N__19522\,
            lcout => \tok.n46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38502\,
            ce => \N__25643\,
            sr => \N__29271\
        );

    \tok.i289_2_lut_3_lut_4_lut_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__36032\,
            in1 => \N__35265\,
            in2 => \N__34060\,
            in3 => \N__36952\,
            lcout => \tok.n8\,
            ltout => \tok.n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6868_2_lut_3_lut_4_lut_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__36953\,
            in1 => \N__30063\,
            in2 => \N__19366\,
            in3 => \N__33950\,
            lcout => \tok.n6425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_325_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__20339\,
            in1 => \N__24329\,
            in2 => \N__19521\,
            in3 => \N__19435\,
            lcout => \tok.n248_adj_884\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6875_2_lut_3_lut_4_lut_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000010"
        )
    port map (
            in0 => \N__36954\,
            in1 => \N__33951\,
            in2 => \N__24433\,
            in3 => \N__23952\,
            lcout => \tok.n6346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i3_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19753\,
            in1 => \N__21264\,
            in2 => \_gnd_net_\,
            in3 => \N__22610\,
            lcout => tc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38453\,
            ce => 'H',
            sr => \N__29169\
        );

    \tok.tc_i2_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21199\,
            in1 => \N__19752\,
            in2 => \_gnd_net_\,
            in3 => \N__22460\,
            lcout => tc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38453\,
            ce => 'H',
            sr => \N__29169\
        );

    \tok.tc_i1_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19751\,
            in1 => \_gnd_net_\,
            in2 => \N__22723\,
            in3 => \N__24959\,
            lcout => tc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38453\,
            ce => 'H',
            sr => \N__29169\
        );

    \tok.tc_i0_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19794\,
            in1 => \N__19750\,
            in2 => \_gnd_net_\,
            in3 => \N__21128\,
            lcout => tc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38453\,
            ce => 'H',
            sr => \N__29169\
        );

    \tok.i2534_2_lut_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__35500\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33267\,
            lcout => \tok.n2557\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_157_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__21004\,
            in1 => \N__33268\,
            in2 => \N__21646\,
            in3 => \N__31230\,
            lcout => OPEN,
            ltout => \tok.n83_adj_756_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6644_2_lut_3_lut_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36316\,
            in2 => \N__19414\,
            in3 => \N__31935\,
            lcout => \tok.n6295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6609_4_lut_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__21055\,
            in1 => \N__22932\,
            in2 => \N__21010\,
            in3 => \N__22874\,
            lcout => OPEN,
            ltout => \tok.ram.n6260_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1528_4_lut_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__21008\,
            in1 => \N__22790\,
            in2 => \N__19573\,
            in3 => \N__31936\,
            lcout => OPEN,
            ltout => \tok.n1565_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_158_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__19570\,
            in1 => \N__35501\,
            in2 => \N__19564\,
            in3 => \N__31231\,
            lcout => OPEN,
            ltout => \tok.n13_adj_757_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_159_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__29710\,
            in1 => \N__25804\,
            in2 => \N__19561\,
            in3 => \N__21056\,
            lcout => n10_adj_906,
            ltout => \n10_adj_906_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_205_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21029\,
            in2 => \N__19558\,
            in3 => \N__19748\,
            lcout => \tok.tc_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i4_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__19749\,
            in1 => \_gnd_net_\,
            in2 => \N__21034\,
            in3 => \N__19537\,
            lcout => tc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38459\,
            ce => 'H',
            sr => \N__29179\
        );

    \tok.i6857_4_lut_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__36251\,
            in1 => \N__19528\,
            in2 => \N__37138\,
            in3 => \N__31319\,
            lcout => \tok.n6622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i303_4_lut_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000110001001"
        )
    port map (
            in0 => \N__36250\,
            in1 => \N__32096\,
            in2 => \N__35523\,
            in3 => \N__31318\,
            lcout => OPEN,
            ltout => \tok.n324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i307_4_lut_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110011"
        )
    port map (
            in0 => \N__19642\,
            in1 => \N__37130\,
            in2 => \N__19531\,
            in3 => \N__33265\,
            lcout => \tok.n239_adj_679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_63_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__35496\,
            in1 => \N__32095\,
            in2 => \_gnd_net_\,
            in3 => \N__31316\,
            lcout => \tok.n225_adj_678\,
            ltout => \tok.n225_adj_678_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6686_3_lut_4_lut_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__31317\,
            in1 => \N__37129\,
            in2 => \N__19645\,
            in3 => \N__36249\,
            lcout => \tok.n6351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2596_rep_330_2_lut_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__34059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32097\,
            lcout => OPEN,
            ltout => \tok.n7456_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i283_4_lut_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001100"
        )
    port map (
            in0 => \N__19636\,
            in1 => \N__25727\,
            in2 => \N__19630\,
            in3 => \N__33266\,
            lcout => \tok.n176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_4_lut_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36232\,
            in1 => \N__34751\,
            in2 => \N__37099\,
            in3 => \N__32043\,
            lcout => \tok.n8_adj_686\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_adj_175_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111100"
        )
    port map (
            in0 => \N__32045\,
            in1 => \N__20560\,
            in2 => \N__34104\,
            in3 => \N__33270\,
            lcout => \tok.n877\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_62_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000101"
        )
    port map (
            in0 => \N__37134\,
            in1 => \N__19651\,
            in2 => \N__35505\,
            in3 => \N__34055\,
            lcout => \tok.n900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_121_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__34752\,
            in1 => \N__19600\,
            in2 => \N__21325\,
            in3 => \N__33269\,
            lcout => OPEN,
            ltout => \tok.n237_adj_724_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_129_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__19579\,
            in1 => \N__20514\,
            in2 => \N__19594\,
            in3 => \N__31235\,
            lcout => \tok.n4893\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_273_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__32044\,
            in1 => \N__20559\,
            in2 => \_gnd_net_\,
            in3 => \N__35423\,
            lcout => \tok.n286\,
            ltout => \tok.n286_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i371_4_lut_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33271\,
            in1 => \N__21316\,
            in2 => \N__19873\,
            in3 => \N__31236\,
            lcout => OPEN,
            ltout => \tok.n394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_298_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19860\,
            in2 => \N__19849\,
            in3 => \N__25120\,
            lcout => \tok.n6143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i7_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25449\,
            in1 => \N__25964\,
            in2 => \_gnd_net_\,
            in3 => \N__26527\,
            lcout => \tok.A_low_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38474\,
            ce => \N__25635\,
            sr => \N__29255\
        );

    \tok.i129_3_lut_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19716\,
            in1 => \N__21265\,
            in2 => \_gnd_net_\,
            in3 => \N__22620\,
            lcout => \tok.tc_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i129_3_lut_adj_209_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24963\,
            in1 => \N__22719\,
            in2 => \_gnd_net_\,
            in3 => \N__19717\,
            lcout => \tok.tc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i129_3_lut_adj_211_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19718\,
            in1 => \_gnd_net_\,
            in2 => \N__19795\,
            in3 => \N__21130\,
            lcout => \tok.tc_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_207_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__22464\,
            in1 => \_gnd_net_\,
            in2 => \N__21198\,
            in3 => \N__19719\,
            lcout => \tok.tc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__25106\,
            in1 => \N__19942\,
            in2 => \_gnd_net_\,
            in3 => \N__36252\,
            lcout => \tok.n6140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6668_3_lut_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__35419\,
            in1 => \N__34753\,
            in2 => \_gnd_net_\,
            in3 => \N__33183\,
            lcout => \tok.n6331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6954_2_lut_3_lut_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__34754\,
            in1 => \N__32059\,
            in2 => \_gnd_net_\,
            in3 => \N__31224\,
            lcout => \tok.n6582\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1500_3_lut_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28483\,
            in1 => \N__22347\,
            in2 => \_gnd_net_\,
            in3 => \N__21991\,
            lcout => \tok.table_wr_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i127_4_lut_4_lut_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001111001111"
        )
    port map (
            in0 => \N__33167\,
            in1 => \N__35396\,
            in2 => \N__31311\,
            in3 => \N__31979\,
            lcout => \tok.n127_adj_772\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i336_4_lut_adj_141_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__23355\,
            in1 => \N__20017\,
            in2 => \N__23746\,
            in3 => \N__31220\,
            lcout => OPEN,
            ltout => \tok.n199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_142_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34612\,
            in2 => \N__19954\,
            in3 => \N__31981\,
            lcout => \tok.n262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2588_3_lut_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__31980\,
            in1 => \N__23993\,
            in2 => \_gnd_net_\,
            in3 => \N__33168\,
            lcout => \tok.n2611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i291_4_lut_4_lut_4_lut_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100100010"
        )
    port map (
            in0 => \N__36215\,
            in1 => \N__34611\,
            in2 => \N__32112\,
            in3 => \N__35397\,
            lcout => \tok.n311_adj_721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_38_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31216\,
            in2 => \_gnd_net_\,
            in3 => \N__33166\,
            lcout => \tok.n4_adj_648\,
            ltout => \tok.n4_adj_648_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i305_4_lut_4_lut_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011001100"
        )
    port map (
            in0 => \N__36214\,
            in1 => \N__34610\,
            in2 => \N__19945\,
            in3 => \N__31978\,
            lcout => \tok.n326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i304_4_lut_4_lut_adj_333_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__31239\,
            in1 => \N__19936\,
            in2 => \N__19905\,
            in3 => \N__31905\,
            lcout => \tok.n210_adj_784\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_4_lut_adj_332_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__31906\,
            in1 => \N__31240\,
            in2 => \N__23113\,
            in3 => \N__37112\,
            lcout => OPEN,
            ltout => \tok.n4842_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_122_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__20437\,
            in1 => \N__20026\,
            in2 => \N__20110\,
            in3 => \N__22943\,
            lcout => \tok.n239_adj_727\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_rep_325_2_lut_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37111\,
            in2 => \_gnd_net_\,
            in3 => \N__31237\,
            lcout => OPEN,
            ltout => \tok.n7451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6956_4_lut_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__34722\,
            in1 => \N__20088\,
            in2 => \N__20107\,
            in3 => \N__20104\,
            lcout => \tok.n6624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i297_4_lut_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000101100"
        )
    port map (
            in0 => \N__20089\,
            in1 => \N__31238\,
            in2 => \N__37135\,
            in3 => \N__33581\,
            lcout => \tok.n164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6833_4_lut_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__34723\,
            in1 => \N__23216\,
            in2 => \N__35503\,
            in3 => \N__33031\,
            lcout => \tok.n6597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i335_4_lut_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001010"
        )
    port map (
            in0 => \N__20011\,
            in1 => \N__20488\,
            in2 => \N__19999\,
            in3 => \N__35415\,
            lcout => \tok.n247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__37124\,
            in1 => \N__37386\,
            in2 => \N__26221\,
            in3 => \N__19987\,
            lcout => OPEN,
            ltout => \tok.n242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_27_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__35377\,
            in1 => \N__37125\,
            in2 => \N__19978\,
            in3 => \N__20278\,
            lcout => \tok.n200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_26_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__20284\,
            in1 => \N__20321\,
            in2 => \N__24337\,
            in3 => \N__20259\,
            lcout => \tok.n248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6630_4_lut_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__37387\,
            in1 => \N__34129\,
            in2 => \N__26615\,
            in3 => \N__21796\,
            lcout => OPEN,
            ltout => \tok.n6606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i8_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25467\,
            in1 => \_gnd_net_\,
            in2 => \N__20272\,
            in3 => \N__28329\,
            lcout => \A_low_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38486\,
            ce => \N__25651\,
            sr => \N__29241\
        );

    \tok.i2_4_lut_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__34005\,
            in1 => \N__27011\,
            in2 => \N__26616\,
            in3 => \N__20269\,
            lcout => OPEN,
            ltout => \tok.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i13_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__25466\,
            in1 => \N__21688\,
            in2 => \N__20263\,
            in3 => \N__20260\,
            lcout => \tok.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38486\,
            ce => \N__25651\,
            sr => \N__29241\
        );

    \tok.i6591_2_lut_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34030\,
            in2 => \_gnd_net_\,
            in3 => \N__29547\,
            lcout => \tok.n6344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_314_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__29549\,
            in1 => \N__26586\,
            in2 => \N__34100\,
            in3 => \N__20203\,
            lcout => OPEN,
            ltout => \tok.n6_adj_878_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i11_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__25479\,
            in1 => \N__20926\,
            in2 => \N__20194\,
            in3 => \N__20191\,
            lcout => \tok.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38490\,
            ce => \N__25649\,
            sr => \N__29270\
        );

    \tok.i2577_2_lut_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__34031\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30258\,
            lcout => OPEN,
            ltout => \tok.n2600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i310_4_lut_adj_311_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__31072\,
            in1 => \N__33417\,
            in2 => \N__20473\,
            in3 => \N__29548\,
            lcout => \tok.n215_adj_876\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6777_4_lut_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__26583\,
            in1 => \N__30259\,
            in2 => \N__30547\,
            in3 => \N__20446\,
            lcout => OPEN,
            ltout => \tok.n6610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i6_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25480\,
            in1 => \_gnd_net_\,
            in2 => \N__20470\,
            in3 => \N__22029\,
            lcout => \tok.A_low_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38490\,
            ce => \N__25649\,
            sr => \N__29270\
        );

    \tok.i310_4_lut_adj_82_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__33416\,
            in1 => \N__24179\,
            in2 => \N__20467\,
            in3 => \N__31071\,
            lcout => \tok.n215_adj_697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001000000000"
        )
    port map (
            in0 => \N__32956\,
            in1 => \N__35279\,
            in2 => \N__36138\,
            in3 => \N__34843\,
            lcout => OPEN,
            ltout => \tok.n269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_110_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111101"
        )
    port map (
            in0 => \N__31069\,
            in1 => \N__26013\,
            in2 => \N__20458\,
            in3 => \N__20575\,
            lcout => \tok.n229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_193_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__32957\,
            in1 => \N__33986\,
            in2 => \N__20455\,
            in3 => \N__21922\,
            lcout => \tok.n205_adj_789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6683_3_lut_4_lut_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35278\,
            in1 => \N__35918\,
            in2 => \N__20425\,
            in3 => \N__32955\,
            lcout => OPEN,
            ltout => \tok.n6341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i311_4_lut_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__20573\,
            in1 => \N__27122\,
            in2 => \N__20347\,
            in3 => \N__31068\,
            lcout => \tok.n170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i5_1_lut_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27262\,
            lcout => \tok.n321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_64_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110100"
        )
    port map (
            in0 => \N__20574\,
            in1 => \N__31956\,
            in2 => \N__20558\,
            in3 => \N__31070\,
            lcout => OPEN,
            ltout => \tok.n238_adj_681_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_65_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__34844\,
            in1 => \N__20530\,
            in2 => \N__20518\,
            in3 => \N__20515\,
            lcout => \tok.n194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6870_2_lut_3_lut_4_lut_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__22191\,
            in1 => \N__33872\,
            in2 => \N__24463\,
            in3 => \N__37046\,
            lcout => \tok.n6396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i9_1_lut_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22190\,
            lcout => \tok.n317_adj_659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2639_3_lut_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__37045\,
            in1 => \N__26831\,
            in2 => \_gnd_net_\,
            in3 => \N__34514\,
            lcout => \tok.n2663\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6100_2_lut_3_lut_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__25376\,
            in1 => \N__33871\,
            in2 => \_gnd_net_\,
            in3 => \N__35127\,
            lcout => \tok.n6183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i6_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27205\,
            in1 => \N__37565\,
            in2 => \_gnd_net_\,
            in3 => \N__36555\,
            lcout => \tok.uart.sender_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38500\,
            ce => \N__27170\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i5_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__33632\,
            in1 => \_gnd_net_\,
            in2 => \N__37567\,
            in3 => \N__20479\,
            lcout => \tok.uart.sender_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38500\,
            ce => \N__27170\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i4_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20869\,
            in1 => \N__37561\,
            in2 => \_gnd_net_\,
            in3 => \N__27544\,
            lcout => \tok.uart.sender_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38500\,
            ce => \N__27170\,
            sr => \_gnd_net_\
        );

    \tok.i6935_3_lut_4_lut_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__27378\,
            in1 => \N__34054\,
            in2 => \N__24437\,
            in3 => \N__36148\,
            lcout => \tok.n6450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i310_4_lut_adj_251_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100100010"
        )
    port map (
            in0 => \N__22245\,
            in1 => \N__33479\,
            in2 => \N__20851\,
            in3 => \N__31090\,
            lcout => OPEN,
            ltout => \tok.n215_adj_830_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6792_4_lut_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__26938\,
            in1 => \N__20836\,
            in2 => \N__20830\,
            in3 => \N__35389\,
            lcout => OPEN,
            ltout => \tok.n6605_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7003_4_lut_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__34483\,
            in1 => \N__35390\,
            in2 => \N__20827\,
            in3 => \N__20800\,
            lcout => \tok.n6604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i309_4_lut_adj_253_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__20812\,
            in1 => \N__22244\,
            in2 => \N__24551\,
            in3 => \N__36149\,
            lcout => \tok.n179_adj_831\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6747_3_lut_4_lut_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__34482\,
            in1 => \N__31089\,
            in2 => \N__27392\,
            in3 => \N__20794\,
            lcout => OPEN,
            ltout => \tok.n6462_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i300_4_lut_adj_245_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__36281\,
            in1 => \N__22243\,
            in2 => \N__20698\,
            in3 => \N__20691\,
            lcout => \tok.n206_adj_823\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i12_1_lut_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23968\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.n314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i309_4_lut_adj_313_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__36150\,
            in1 => \N__20956\,
            in2 => \N__29596\,
            in3 => \N__24540\,
            lcout => \tok.n179_adj_877\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i309_4_lut_adj_83_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__24541\,
            in1 => \N__36152\,
            in2 => \N__24180\,
            in3 => \N__20950\,
            lcout => \tok.n179_adj_698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6844_4_lut_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__35384\,
            in1 => \N__26931\,
            in2 => \N__22381\,
            in3 => \N__20944\,
            lcout => OPEN,
            ltout => \tok.n6553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6995_4_lut_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__34792\,
            in1 => \N__20935\,
            in2 => \N__20929\,
            in3 => \N__35386\,
            lcout => \tok.n6552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6948_4_lut_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__35388\,
            in1 => \N__20914\,
            in2 => \N__22357\,
            in3 => \N__34794\,
            lcout => \tok.n6537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6772_4_lut_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__24073\,
            in1 => \N__21892\,
            in2 => \N__26937\,
            in3 => \N__35385\,
            lcout => OPEN,
            ltout => \tok.n6541_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6847_4_lut_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__35387\,
            in1 => \N__20875\,
            in2 => \N__20899\,
            in3 => \N__34793\,
            lcout => \tok.n6540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i309_4_lut_adj_59_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__20884\,
            in1 => \N__36151\,
            in2 => \N__24554\,
            in3 => \N__32354\,
            lcout => \tok.n179_adj_673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i0_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24696\,
            in1 => \N__28733\,
            in2 => \_gnd_net_\,
            in3 => \N__21089\,
            lcout => \tok.C_stk.tail_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38454\,
            ce => \N__28909\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i6146_3_lut_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21069\,
            in1 => \N__28116\,
            in2 => \_gnd_net_\,
            in3 => \N__21171\,
            lcout => OPEN,
            ltout => \tok.C_stk.n6230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i0_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__28054\,
            in1 => \N__27929\,
            in2 => \N__21133\,
            in3 => \N__21129\,
            lcout => c_stk_r_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38454\,
            ce => \N__28909\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i8_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__28734\,
            in1 => \_gnd_net_\,
            in2 => \N__21073\,
            in3 => \N__24670\,
            lcout => tail_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38454\,
            ce => \N__28909\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i4_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28747\,
            in1 => \N__20977\,
            in2 => \_gnd_net_\,
            in3 => \N__21009\,
            lcout => \tok.C_stk.tail_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38460\,
            ce => \N__28918\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i6155_3_lut_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20985\,
            in1 => \N__28098\,
            in2 => \_gnd_net_\,
            in3 => \N__21061\,
            lcout => OPEN,
            ltout => \tok.C_stk.n6239_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i4_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27924\,
            in1 => \N__28047\,
            in2 => \N__21037\,
            in3 => \N__21033\,
            lcout => \tok.c_stk_r_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38460\,
            ce => \N__28918\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i12_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__20986\,
            in1 => \_gnd_net_\,
            in2 => \N__20968\,
            in3 => \N__28742\,
            lcout => \tok.tail_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38460\,
            ce => \N__28918\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i20_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28743\,
            in1 => \N__21220\,
            in2 => \_gnd_net_\,
            in3 => \N__20976\,
            lcout => \tok.C_stk.tail_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38460\,
            ce => \N__28918\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i28_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20964\,
            in1 => \N__21211\,
            in2 => \_gnd_net_\,
            in3 => \N__28744\,
            lcout => \tok.tail_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38460\,
            ce => \N__28918\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i36_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28745\,
            in1 => \N__24870\,
            in2 => \_gnd_net_\,
            in3 => \N__21219\,
            lcout => \tok.C_stk.tail_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38460\,
            ce => \N__28918\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i44_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24751\,
            in1 => \N__21210\,
            in2 => \_gnd_net_\,
            in3 => \N__28746\,
            lcout => \tok.tail_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38460\,
            ce => \N__28918\,
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_140_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__21562\,
            in1 => \N__33274\,
            in2 => \N__22435\,
            in3 => \N__31297\,
            lcout => OPEN,
            ltout => \tok.n83_adj_723_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6979_2_lut_3_lut_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__36315\,
            in1 => \_gnd_net_\,
            in2 => \N__21202\,
            in3 => \N__31879\,
            lcout => \tok.n6664\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_148_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__21292\,
            in1 => \N__29706\,
            in2 => \N__22501\,
            in3 => \N__25808\,
            lcout => n10_adj_908,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_181_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__33273\,
            in1 => \_gnd_net_\,
            in2 => \N__36325\,
            in3 => \_gnd_net_\,
            lcout => \tok.n2573\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_194_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36311\,
            in2 => \_gnd_net_\,
            in3 => \N__33272\,
            lcout => \tok.n4_adj_726\,
            ltout => \tok.n4_adj_726_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6600_4_lut_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__22432\,
            in1 => \N__22497\,
            in2 => \N__21178\,
            in3 => \N__22870\,
            lcout => OPEN,
            ltout => \tok.ram.n6257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1564_4_lut_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__31880\,
            in1 => \N__22775\,
            in2 => \N__21175\,
            in3 => \N__22433\,
            lcout => OPEN,
            ltout => \tok.n1600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__31298\,
            in1 => \N__21301\,
            in2 => \N__21295\,
            in3 => \N__35331\,
            lcout => \tok.n13_adj_742\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6675_4_lut_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__22914\,
            in1 => \N__22583\,
            in2 => \N__22660\,
            in3 => \N__22868\,
            lcout => OPEN,
            ltout => \tok.n6301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i124_4_lut_adj_152_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__22584\,
            in1 => \N__32122\,
            in2 => \N__21286\,
            in3 => \N__22791\,
            lcout => OPEN,
            ltout => \tok.n80_adj_751_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i126_4_lut_adj_155_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__31323\,
            in1 => \N__21277\,
            in2 => \N__21283\,
            in3 => \N__35330\,
            lcout => \tok.n89_adj_754\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_149_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__22582\,
            in1 => \N__33275\,
            in2 => \N__21244\,
            in3 => \N__31320\,
            lcout => OPEN,
            ltout => \tok.n83_adj_746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6647_2_lut_3_lut_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36253\,
            in2 => \N__21280\,
            in3 => \N__32121\,
            lcout => \tok.n6297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_156_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__21271\,
            in1 => \N__25807\,
            in2 => \N__29724\,
            in3 => \N__22659\,
            lcout => n92_adj_898,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i335_4_lut_adj_135_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111001010100"
        )
    port map (
            in0 => \N__31321\,
            in1 => \N__21243\,
            in2 => \N__33300\,
            in3 => \N__21487\,
            lcout => \tok.n2700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_3_lut_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21486\,
            in1 => \N__33279\,
            in2 => \_gnd_net_\,
            in3 => \N__31322\,
            lcout => \tok.n236_adj_737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_4_lut_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__35490\,
            in1 => \N__37091\,
            in2 => \N__34113\,
            in3 => \N__36233\,
            lcout => \tok.n14_adj_683\,
            ltout => \tok.n14_adj_683_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_adj_67_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21370\,
            in3 => \N__21381\,
            lcout => \tok.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.stall_I_0_400_i15_2_lut_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__35492\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37093\,
            lcout => OPEN,
            ltout => \tok.n15_adj_807_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_222_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23119\,
            in1 => \N__21367\,
            in2 => \N__21352\,
            in3 => \N__33485\,
            lcout => \tok.n903\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.i406_4_lut_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__21382\,
            in1 => \N__23002\,
            in2 => \N__21337\,
            in3 => \N__28004\,
            lcout => \tok.C_stk.n449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_111_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111011"
        )
    port map (
            in0 => \N__36235\,
            in1 => \N__35493\,
            in2 => \N__26131\,
            in3 => \N__37097\,
            lcout => \tok.n278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6855_4_lut_4_lut_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000111111111"
        )
    port map (
            in0 => \N__35491\,
            in1 => \N__36234\,
            in2 => \N__32126\,
            in3 => \N__37092\,
            lcout => \tok.n6621\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i362_4_lut_4_lut_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000100010"
        )
    port map (
            in0 => \N__32106\,
            in1 => \N__34790\,
            in2 => \N__36310\,
            in3 => \N__37098\,
            lcout => \tok.n241_adj_747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6829_4_lut_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010001010"
        )
    port map (
            in0 => \N__31877\,
            in1 => \N__22039\,
            in2 => \N__34759\,
            in3 => \N__21451\,
            lcout => \tok.n6593\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_137_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__31161\,
            in1 => \N__21480\,
            in2 => \_gnd_net_\,
            in3 => \N__36254\,
            lcout => \tok.n4925\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6726_2_lut_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21445\,
            in2 => \_gnd_net_\,
            in3 => \N__33165\,
            lcout => OPEN,
            ltout => \tok.n6578_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6840_4_lut_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010100000"
        )
    port map (
            in0 => \N__21406\,
            in1 => \N__21433\,
            in2 => \N__21418\,
            in3 => \N__31876\,
            lcout => \tok.n6581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_219_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31160\,
            lcout => \tok.n4_adj_739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6953_4_lut_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110001"
        )
    port map (
            in0 => \N__31163\,
            in1 => \N__21400\,
            in2 => \N__23143\,
            in3 => \N__36255\,
            lcout => \tok.n6580\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_4_lut_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__31875\,
            in1 => \N__33164\,
            in2 => \N__34758\,
            in3 => \N__31159\,
            lcout => \tok.n4_adj_684\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_228_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__31162\,
            in1 => \N__25238\,
            in2 => \N__22081\,
            in3 => \N__31878\,
            lcout => \tok.n273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_107_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001000100"
        )
    port map (
            in0 => \N__23302\,
            in1 => \N__31174\,
            in2 => \N__36303\,
            in3 => \N__23742\,
            lcout => \tok.n251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6854_2_lut_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__34614\,
            in1 => \N__28207\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \tok.n6620_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i296_4_lut_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__36206\,
            in1 => \N__23741\,
            in2 => \N__21373\,
            in3 => \N__33185\,
            lcout => OPEN,
            ltout => \tok.n167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_124_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21580\,
            in2 => \N__21574\,
            in3 => \N__24318\,
            lcout => \tok.n179_adj_730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_165_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__21520\,
            in1 => \N__21571\,
            in2 => \N__36304\,
            in3 => \N__33186\,
            lcout => \tok.n186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i288_4_lut_4_lut_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__31173\,
            in1 => \N__23259\,
            in2 => \N__21561\,
            in3 => \N__32071\,
            lcout => OPEN,
            ltout => \tok.n209_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6959_3_lut_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010000"
        )
    port map (
            in0 => \N__37113\,
            in1 => \N__34613\,
            in2 => \N__21535\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \tok.n6625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_120_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__33184\,
            in1 => \N__35494\,
            in2 => \N__21532\,
            in3 => \N__21529\,
            lcout => \tok.n162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i320_4_lut_4_lut_4_lut_adj_85_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010110000000"
        )
    port map (
            in0 => \N__31165\,
            in1 => \N__28225\,
            in2 => \N__32116\,
            in3 => \N__27022\,
            lcout => OPEN,
            ltout => \tok.n168_adj_700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6621_4_lut_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__32460\,
            in1 => \N__36341\,
            in2 => \N__21523\,
            in3 => \N__27346\,
            lcout => \tok.n6569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2525_2_lut_4_lut_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32034\,
            in1 => \N__34750\,
            in2 => \N__36256\,
            in3 => \N__33287\,
            lcout => \tok.n2548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i309_4_lut_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__27023\,
            in1 => \N__36102\,
            in2 => \N__21502\,
            in3 => \N__24556\,
            lcout => OPEN,
            ltout => \tok.n179_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6997_4_lut_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__26875\,
            in1 => \N__35442\,
            in2 => \N__21691\,
            in3 => \N__34846\,
            lcout => \tok.n6546\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i304_4_lut_4_lut_adj_315_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__21607\,
            in1 => \N__32041\,
            in2 => \N__21682\,
            in3 => \N__31167\,
            lcout => \tok.n210_adj_816\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i304_4_lut_4_lut_adj_317_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__31166\,
            in1 => \N__21642\,
            in2 => \N__32117\,
            in3 => \N__21859\,
            lcout => \tok.n210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_66_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32033\,
            in2 => \_gnd_net_\,
            in3 => \N__31164\,
            lcout => \tok.n5_adj_682\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_234_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__26305\,
            in1 => \N__21586\,
            in2 => \N__32251\,
            in3 => \N__36098\,
            lcout => \tok.n258_adj_814\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i303_4_lut_adj_235_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__35374\,
            in1 => \N__26410\,
            in2 => \N__23629\,
            in3 => \N__25894\,
            lcout => OPEN,
            ltout => \tok.n252_adj_815_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_240_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__35376\,
            in1 => \N__21616\,
            in2 => \N__21610\,
            in3 => \N__34845\,
            lcout => \tok.n4_adj_818\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_adj_226_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__32247\,
            in1 => \N__21606\,
            in2 => \N__26392\,
            in3 => \N__37122\,
            lcout => \tok.n255_adj_808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_218_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__34821\,
            in1 => \N__36097\,
            in2 => \_gnd_net_\,
            in3 => \N__35373\,
            lcout => \tok.n872\,
            ltout => \tok.n872_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i306_4_lut_adj_239_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__21814\,
            in1 => \N__37123\,
            in2 => \N__21808\,
            in3 => \N__23878\,
            lcout => OPEN,
            ltout => \tok.n174_adj_817_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_242_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010000"
        )
    port map (
            in0 => \N__33217\,
            in1 => \N__34040\,
            in2 => \N__21805\,
            in3 => \N__21802\,
            lcout => \tok.n205_adj_820\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6888_2_lut_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34035\,
            in2 => \_gnd_net_\,
            in3 => \N__26736\,
            lcout => \tok.n6365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_274_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__26585\,
            in1 => \N__26738\,
            in2 => \N__34101\,
            in3 => \N__21790\,
            lcout => OPEN,
            ltout => \tok.n6_adj_843_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i10_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__24574\,
            in1 => \N__25477\,
            in2 => \N__21781\,
            in3 => \N__21778\,
            lcout => \tok.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38496\,
            ce => \N__25645\,
            sr => \N__29261\
        );

    \tok.i6920_2_lut_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__34036\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27293\,
            lcout => OPEN,
            ltout => \tok.n6440_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i310_4_lut_adj_271_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__33429\,
            in1 => \N__26737\,
            in2 => \N__21697\,
            in3 => \N__31213\,
            lcout => \tok.n215_adj_841\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6794_4_lut_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__26584\,
            in1 => \N__27294\,
            in2 => \N__23062\,
            in3 => \N__21865\,
            lcout => OPEN,
            ltout => \tok.n6612_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i5_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25478\,
            in2 => \N__21694\,
            in3 => \N__23856\,
            lcout => \tok.A_low_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38496\,
            ce => \N__25645\,
            sr => \N__29261\
        );

    \tok.i310_4_lut_adj_58_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__31212\,
            in1 => \N__33428\,
            in2 => \N__21901\,
            in3 => \N__32372\,
            lcout => \tok.n215_adj_672\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_170_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__21823\,
            in1 => \N__35372\,
            in2 => \N__34791\,
            in3 => \N__21880\,
            lcout => OPEN,
            ltout => \tok.n4_adj_769_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_171_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__33980\,
            in2 => \N__21868\,
            in3 => \N__23752\,
            lcout => \tok.n205_adj_770\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_231_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__35764\,
            in1 => \N__31955\,
            in2 => \_gnd_net_\,
            in3 => \N__31211\,
            lcout => \tok.n190\,
            ltout => \tok.n190_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_adj_161_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__26384\,
            in1 => \N__21858\,
            in2 => \N__21835\,
            in3 => \N__36797\,
            lcout => OPEN,
            ltout => \tok.n255_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_166_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__35766\,
            in1 => \N__21832\,
            in2 => \N__21826\,
            in3 => \N__26315\,
            lcout => \tok.n258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6939_3_lut_4_lut_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__22240\,
            in1 => \N__33979\,
            in2 => \N__24460\,
            in3 => \N__35765\,
            lcout => \tok.n6390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6787_2_lut_3_lut_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__27541\,
            in1 => \N__35370\,
            in2 => \_gnd_net_\,
            in3 => \N__31210\,
            lcout => OPEN,
            ltout => \tok.n6508_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i305_4_lut_adj_202_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__35371\,
            in1 => \N__23400\,
            in2 => \N__21817\,
            in3 => \N__35763\,
            lcout => \tok.n213_adj_795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_98_i6_3_lut_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111111010"
        )
    port map (
            in0 => \N__27543\,
            in1 => \_gnd_net_\,
            in2 => \N__36322\,
            in3 => \N__37063\,
            lcout => OPEN,
            ltout => \tok.n207_adj_771_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i305_4_lut_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__22057\,
            in1 => \N__36279\,
            in2 => \N__22042\,
            in3 => \N__35375\,
            lcout => \tok.n213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6836_3_lut_4_lut_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36554\,
            in1 => \N__33064\,
            in2 => \N__36320\,
            in3 => \N__30954\,
            lcout => \tok.n6583\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i318_4_lut_adj_179_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__22028\,
            in1 => \N__34523\,
            in2 => \N__23677\,
            in3 => \N__36280\,
            lcout => OPEN,
            ltout => \tok.n207_adj_776_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6823_4_lut_4_lut_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__31897\,
            in1 => \N__21946\,
            in2 => \N__21940\,
            in3 => \N__24287\,
            lcout => OPEN,
            ltout => \tok.n6529_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i306_4_lut_adj_188_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__37064\,
            in1 => \N__24223\,
            in2 => \N__21937\,
            in3 => \N__21934\,
            lcout => \tok.n174_adj_785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2641_2_lut_3_lut_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__27542\,
            in1 => \_gnd_net_\,
            in2 => \N__36321\,
            in3 => \N__33065\,
            lcout => \tok.n2665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_261_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__30955\,
            in1 => \_gnd_net_\,
            in2 => \N__33223\,
            in3 => \N__31896\,
            lcout => \tok.n847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i369_4_lut_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010001"
        )
    port map (
            in0 => \N__26504\,
            in1 => \N__30533\,
            in2 => \N__22264\,
            in3 => \N__36147\,
            lcout => \tok.n229_adj_861\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6662_3_lut_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__35379\,
            in1 => \_gnd_net_\,
            in2 => \N__34102\,
            in3 => \N__31086\,
            lcout => \tok.n6320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6895_2_lut_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__22228\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34045\,
            lcout => OPEN,
            ltout => \tok.n6380_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i310_4_lut_adj_46_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__33475\,
            in1 => \N__32220\,
            in2 => \N__22108\,
            in3 => \N__31087\,
            lcout => OPEN,
            ltout => \tok.n215_adj_656_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6745_4_lut_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__26932\,
            in1 => \N__24565\,
            in2 => \N__22105\,
            in3 => \N__35380\,
            lcout => \tok.n6544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i338_4_lut_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110011"
        )
    port map (
            in0 => \N__33219\,
            in1 => \N__34842\,
            in2 => \N__22093\,
            in3 => \N__22102\,
            lcout => \tok.n256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_225_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34041\,
            in2 => \_gnd_net_\,
            in3 => \N__35378\,
            lcout => \tok.n4_adj_719\,
            ltout => \tok.n4_adj_719_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_227_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33218\,
            in1 => \N__34841\,
            in2 => \N__22084\,
            in3 => \N__36571\,
            lcout => \tok.n10_adj_809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i309_4_lut_adj_330_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__22066\,
            in1 => \N__36145\,
            in2 => \N__24555\,
            in3 => \N__23988\,
            lcout => \tok.n179_adj_888\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6938_3_lut_4_lut_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__36146\,
            in1 => \N__24452\,
            in2 => \N__34103\,
            in3 => \N__37465\,
            lcout => OPEN,
            ltout => \tok.n6404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6821_4_lut_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__35382\,
            in1 => \N__26927\,
            in2 => \N__22402\,
            in3 => \N__23890\,
            lcout => OPEN,
            ltout => \tok.n6550_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6999_4_lut_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__22399\,
            in1 => \N__35383\,
            in2 => \N__22393\,
            in3 => \N__34795\,
            lcout => \tok.n6549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6863_2_lut_3_lut_4_lut_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__34046\,
            in1 => \N__37065\,
            in2 => \N__24461\,
            in3 => \N__30323\,
            lcout => \tok.n6442\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6937_3_lut_4_lut_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100010"
        )
    port map (
            in0 => \N__36143\,
            in1 => \N__24448\,
            in2 => \N__30074\,
            in3 => \N__34047\,
            lcout => \tok.n6419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6674_3_lut_4_lut_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__34048\,
            in1 => \N__36144\,
            in2 => \N__24462\,
            in3 => \N__23987\,
            lcout => OPEN,
            ltout => \tok.n6337_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6771_4_lut_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__26926\,
            in1 => \N__22372\,
            in2 => \N__22360\,
            in3 => \N__35381\,
            lcout => \tok.n6538\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i5_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28753\,
            in1 => \N__22540\,
            in2 => \_gnd_net_\,
            in3 => \N__22278\,
            lcout => \tok.C_stk.tail_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38461\,
            ce => \N__28919\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i6152_3_lut_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22548\,
            in1 => \N__28122\,
            in2 => \_gnd_net_\,
            in3 => \N__22348\,
            lcout => OPEN,
            ltout => \tok.C_stk.n6236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i5_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__28051\,
            in1 => \N__27940\,
            in2 => \N__22318\,
            in3 => \N__22315\,
            lcout => \tok.c_stk_r_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38461\,
            ce => \N__28919\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i13_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22549\,
            in1 => \_gnd_net_\,
            in2 => \N__22531\,
            in3 => \N__28748\,
            lcout => \tok.tail_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38461\,
            ce => \N__28919\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i21_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28749\,
            in1 => \N__22519\,
            in2 => \_gnd_net_\,
            in3 => \N__22539\,
            lcout => \tok.C_stk.tail_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38461\,
            ce => \N__28919\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i29_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22527\,
            in1 => \N__22510\,
            in2 => \_gnd_net_\,
            in3 => \N__28750\,
            lcout => \tok.tail_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38461\,
            ce => \N__28919\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i37_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28751\,
            in1 => \N__24618\,
            in2 => \_gnd_net_\,
            in3 => \N__22518\,
            lcout => \tok.C_stk.tail_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38461\,
            ce => \N__28919\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i45_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25033\,
            in1 => \N__22509\,
            in2 => \_gnd_net_\,
            in3 => \N__28752\,
            lcout => \tok.tail_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38461\,
            ce => \N__28919\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i2_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28739\,
            in1 => \N__22699\,
            in2 => \_gnd_net_\,
            in3 => \N__22434\,
            lcout => \tok.C_stk.tail_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38465\,
            ce => \N__28905\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i6161_3_lut_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22410\,
            in1 => \N__28103\,
            in2 => \_gnd_net_\,
            in3 => \N__22496\,
            lcout => OPEN,
            ltout => \tok.C_stk.n6245_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i2_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__28050\,
            in1 => \N__27933\,
            in2 => \N__22468\,
            in3 => \N__22465\,
            lcout => \tok.c_stk_r_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38465\,
            ce => \N__28905\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i10_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22411\,
            in1 => \_gnd_net_\,
            in2 => \N__22690\,
            in3 => \N__28736\,
            lcout => \tok.tail_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38465\,
            ce => \N__28905\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i18_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28737\,
            in1 => \N__22678\,
            in2 => \_gnd_net_\,
            in3 => \N__22698\,
            lcout => \tok.C_stk.tail_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38465\,
            ce => \N__28905\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i26_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22686\,
            in1 => \N__22669\,
            in2 => \_gnd_net_\,
            in3 => \N__28738\,
            lcout => \tok.tail_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38465\,
            ce => \N__28905\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i34_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28740\,
            in1 => \N__24856\,
            in2 => \_gnd_net_\,
            in3 => \N__22677\,
            lcout => \tok.C_stk.tail_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38465\,
            ce => \N__28905\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i42_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27781\,
            in1 => \N__22668\,
            in2 => \_gnd_net_\,
            in3 => \N__28741\,
            lcout => \tok.tail_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38465\,
            ce => \N__28905\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i3_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28679\,
            in1 => \N__22558\,
            in2 => \_gnd_net_\,
            in3 => \N__22585\,
            lcout => \tok.C_stk.tail_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38470\,
            ce => \N__28921\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i6158_3_lut_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28102\,
            in1 => \N__22566\,
            in2 => \_gnd_net_\,
            in3 => \N__22655\,
            lcout => OPEN,
            ltout => \tok.C_stk.n6242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i3_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__28049\,
            in1 => \N__27925\,
            in2 => \N__22624\,
            in3 => \N__22621\,
            lcout => \tok.c_stk_r_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38470\,
            ce => \N__28921\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i11_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22972\,
            in1 => \N__22567\,
            in2 => \_gnd_net_\,
            in3 => \N__28675\,
            lcout => \tok.C_stk.tail_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38470\,
            ce => \N__28921\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i19_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28676\,
            in1 => \N__22963\,
            in2 => \_gnd_net_\,
            in3 => \N__22557\,
            lcout => \tok.C_stk.tail_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38470\,
            ce => \N__28921\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i27_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22971\,
            in1 => \N__22954\,
            in2 => \_gnd_net_\,
            in3 => \N__28677\,
            lcout => \tok.C_stk.tail_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38470\,
            ce => \N__28921\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i35_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28678\,
            in1 => \N__22962\,
            in2 => \_gnd_net_\,
            in3 => \N__24636\,
            lcout => \tok.C_stk.tail_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38470\,
            ce => \N__28921\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i43_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24840\,
            in1 => \N__22953\,
            in2 => \_gnd_net_\,
            in3 => \N__28680\,
            lcout => \tok.C_stk.tail_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38470\,
            ce => \N__28921\,
            sr => \_gnd_net_\
        );

    \tok.i6605_4_lut_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__22915\,
            in1 => \N__24995\,
            in2 => \N__24934\,
            in3 => \N__22869\,
            lcout => OPEN,
            ltout => \tok.n6291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i124_4_lut_adj_133_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__32120\,
            in1 => \N__22779\,
            in2 => \N__22744\,
            in3 => \N__24933\,
            lcout => OPEN,
            ltout => \tok.n80_adj_735_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i126_4_lut_adj_136_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__35517\,
            in1 => \N__22735\,
            in2 => \N__22741\,
            in3 => \N__31328\,
            lcout => \tok.n89_adj_736\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_132_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010001000"
        )
    port map (
            in0 => \N__31327\,
            in1 => \N__24929\,
            in2 => \N__23296\,
            in3 => \N__33264\,
            lcout => OPEN,
            ltout => \tok.n83_adj_725_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6641_2_lut_3_lut_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36299\,
            in2 => \N__22738\,
            in3 => \N__32119\,
            lcout => \tok.n6287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_139_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__24996\,
            in1 => \N__25797\,
            in2 => \N__29723\,
            in3 => \N__22729\,
            lcout => n92,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i307_3_lut_3_lut_3_lut_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111101110"
        )
    port map (
            in0 => \N__33263\,
            in1 => \N__32118\,
            in2 => \_gnd_net_\,
            in3 => \N__31326\,
            lcout => \tok.n180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_147_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31329\,
            in1 => \N__34820\,
            in2 => \N__26511\,
            in3 => \N__36533\,
            lcout => \tok.n4926\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2664_4_lut_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33283\,
            in1 => \N__36296\,
            in2 => \N__34839\,
            in3 => \N__35516\,
            lcout => OPEN,
            ltout => \tok.n2692_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i359_4_lut_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001000"
        )
    port map (
            in0 => \N__23008\,
            in1 => \N__25875\,
            in2 => \N__23023\,
            in3 => \N__31303\,
            lcout => \tok.n217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_rep_28_2_lut_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35515\,
            in2 => \_gnd_net_\,
            in3 => \N__34785\,
            lcout => \tok.n7154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36295\,
            in1 => \N__32098\,
            in2 => \_gnd_net_\,
            in3 => \N__33282\,
            lcout => \tok.n815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_rep_332_2_lut_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37110\,
            lcout => \tok.n7458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_3_lut_4_lut_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__31302\,
            in1 => \N__34786\,
            in2 => \N__33301\,
            in3 => \N__32107\,
            lcout => \tok.n6_adj_701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_138_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001101"
        )
    port map (
            in0 => \N__22996\,
            in1 => \N__22990\,
            in2 => \N__33489\,
            in3 => \N__32100\,
            lcout => \tok.n239_adj_738\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_4_lut_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34106\,
            in2 => \_gnd_net_\,
            in3 => \N__36298\,
            lcout => \tok.n864\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2679_3_lut_3_lut_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101110111"
        )
    port map (
            in0 => \N__32123\,
            in1 => \N__33288\,
            in2 => \_gnd_net_\,
            in3 => \N__31249\,
            lcout => \tok.n2679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_336_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36297\,
            in2 => \_gnd_net_\,
            in3 => \N__34797\,
            lcout => \tok.n5_adj_821\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_334_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__34105\,
            in1 => \N__25368\,
            in2 => \_gnd_net_\,
            in3 => \N__29408\,
            lcout => \tok.n17\,
            ltout => \tok.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_243_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__23106\,
            in1 => \N__23092\,
            in2 => \N__23086\,
            in3 => \N__25737\,
            lcout => \tok.n2559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6809_4_lut_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__32551\,
            in1 => \N__32601\,
            in2 => \N__23083\,
            in3 => \N__27393\,
            lcout => OPEN,
            ltout => \tok.n6562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i315_4_lut_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__35520\,
            in1 => \N__23074\,
            in2 => \N__23065\,
            in3 => \N__34799\,
            lcout => \tok.n338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6867_4_lut_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34798\,
            in1 => \N__23470\,
            in2 => \N__25110\,
            in3 => \N__35521\,
            lcout => \tok.n6637\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_123_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__23047\,
            in1 => \N__29458\,
            in2 => \N__23227\,
            in3 => \N__35468\,
            lcout => OPEN,
            ltout => \tok.n197_adj_729_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_125_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__36219\,
            in1 => \N__23041\,
            in2 => \N__23314\,
            in3 => \N__23311\,
            lcout => \tok.n203_adj_731\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2521_2_lut_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23549\,
            in2 => \_gnd_net_\,
            in3 => \N__34800\,
            lcout => \tok.n2544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_3_lut_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110100000"
        )
    port map (
            in0 => \N__35467\,
            in1 => \_gnd_net_\,
            in2 => \N__36305\,
            in3 => \N__33290\,
            lcout => \tok.n256_adj_749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2598_rep_349_2_lut_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37137\,
            in2 => \_gnd_net_\,
            in3 => \N__34802\,
            lcout => OPEN,
            ltout => \tok.n7475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6981_4_lut_4_lut_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__35466\,
            in1 => \N__23295\,
            in2 => \N__23263\,
            in3 => \N__32125\,
            lcout => \tok.n6645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6984_4_lut_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__23260\,
            in1 => \N__37136\,
            in2 => \N__23239\,
            in3 => \N__34801\,
            lcout => \tok.n6628\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i337_4_lut_adj_145_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001010101"
        )
    port map (
            in0 => \N__23217\,
            in1 => \N__32124\,
            in2 => \N__37891\,
            in3 => \N__33289\,
            lcout => \tok.n241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_112_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__36287\,
            in1 => \N__27129\,
            in2 => \N__37126\,
            in3 => \N__23329\,
            lcout => OPEN,
            ltout => \tok.n284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_113_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__36230\,
            in1 => \N__23131\,
            in2 => \N__23122\,
            in3 => \N__26023\,
            lcout => OPEN,
            ltout => \tok.n244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_116_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110010"
        )
    port map (
            in0 => \N__25672\,
            in1 => \N__27461\,
            in2 => \N__23380\,
            in3 => \N__34076\,
            lcout => OPEN,
            ltout => \tok.n4_adj_720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i2_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__25481\,
            in1 => \N__23553\,
            in2 => \N__23377\,
            in3 => \N__27577\,
            lcout => \tok.A_low_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38491\,
            ce => \N__25607\,
            sr => \N__29204\
        );

    \tok.inv_105_i2_1_lut_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27457\,
            lcout => \tok.n145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_108_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001101"
        )
    port map (
            in0 => \N__27090\,
            in1 => \N__36285\,
            in2 => \N__34813\,
            in3 => \N__23365\,
            lcout => OPEN,
            ltout => \tok.n4_adj_714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_4_lut_adj_316_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110010"
        )
    port map (
            in0 => \N__36286\,
            in1 => \N__23359\,
            in2 => \N__23332\,
            in3 => \N__32042\,
            lcout => \tok.n218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6795_2_lut_4_lut_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__34075\,
            in1 => \N__37069\,
            in2 => \N__27509\,
            in3 => \N__36284\,
            lcout => \tok.n6525\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i57_4_lut_3_lut_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100000"
        )
    port map (
            in0 => \N__31206\,
            in1 => \_gnd_net_\,
            in2 => \N__33281\,
            in3 => \N__31973\,
            lcout => \tok.n39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6628_4_lut_4_lut_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000100000000"
        )
    port map (
            in0 => \N__31974\,
            in1 => \N__33196\,
            in2 => \N__36323\,
            in3 => \N__31207\,
            lcout => OPEN,
            ltout => \tok.n6269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i58_4_lut_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__23323\,
            in1 => \N__35455\,
            in2 => \N__23317\,
            in3 => \N__36293\,
            lcout => \tok.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_104_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31958\,
            in2 => \_gnd_net_\,
            in3 => \N__33192\,
            lcout => \tok.n6_adj_676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6765_4_lut_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__31960\,
            in1 => \N__23653\,
            in2 => \N__23617\,
            in3 => \N__23638\,
            lcout => \tok.n6486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6783_4_lut_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__23612\,
            in1 => \N__23581\,
            in2 => \N__23569\,
            in3 => \N__31959\,
            lcout => \tok.n6510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i336_4_lut_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110001000"
        )
    port map (
            in0 => \N__31208\,
            in1 => \N__27471\,
            in2 => \N__23554\,
            in3 => \N__37073\,
            lcout => \tok.n208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6824_4_lut_4_lut_4_lut_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__34697\,
            in1 => \N__33197\,
            in2 => \N__32094\,
            in3 => \N__31209\,
            lcout => \tok.n6589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i17_4_lut_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__34062\,
            in1 => \N__33635\,
            in2 => \N__32605\,
            in3 => \N__32077\,
            lcout => OPEN,
            ltout => \tok.n6_adj_728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_128_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__23440\,
            in1 => \N__32550\,
            in2 => \N__23428\,
            in3 => \N__34063\,
            lcout => OPEN,
            ltout => \tok.n200_adj_732_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_130_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__35519\,
            in1 => \N__34107\,
            in2 => \N__23425\,
            in3 => \N__23422\,
            lcout => \tok.n6_adj_733\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6778_2_lut_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32469\,
            in2 => \_gnd_net_\,
            in3 => \N__23401\,
            lcout => \tok.n6501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6769_3_lut_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__34061\,
            in1 => \N__33634\,
            in2 => \_gnd_net_\,
            in3 => \N__31130\,
            lcout => \tok.n6484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i318_4_lut_adj_230_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000000010"
        )
    port map (
            in0 => \N__28334\,
            in1 => \N__36292\,
            in2 => \N__34803\,
            in3 => \N__23675\,
            lcout => OPEN,
            ltout => \tok.n207_adj_811_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6834_4_lut_4_lut_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__24324\,
            in1 => \N__23863\,
            in2 => \N__23881\,
            in3 => \N__32076\,
            lcout => \tok.n6481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i305_4_lut_adj_229_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__32407\,
            in1 => \N__35518\,
            in2 => \N__23872\,
            in3 => \N__36291\,
            lcout => \tok.n213_adj_810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i318_4_lut_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__35779\,
            in1 => \N__34682\,
            in2 => \N__23857\,
            in3 => \N__23676\,
            lcout => OPEN,
            ltout => \tok.n207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6822_4_lut_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__24323\,
            in1 => \N__27058\,
            in2 => \N__23767\,
            in3 => \N__24472\,
            lcout => OPEN,
            ltout => \tok.n6572_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i306_4_lut_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__24219\,
            in1 => \N__23764\,
            in2 => \N__23755\,
            in3 => \N__36796\,
            lcout => \tok.n174_adj_768\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_3_lut_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__34680\,
            in1 => \N__23732\,
            in2 => \_gnd_net_\,
            in3 => \N__31943\,
            lcout => \tok.n26_adj_763\,
            ltout => \tok.n26_adj_763_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i318_4_lut_adj_203_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__25993\,
            in1 => \N__35767\,
            in2 => \N__23656\,
            in3 => \N__34681\,
            lcout => OPEN,
            ltout => \tok.n207_adj_796_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6816_4_lut_4_lut_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__24322\,
            in1 => \N__24232\,
            in2 => \N__24226\,
            in3 => \N__31944\,
            lcout => OPEN,
            ltout => \tok.n6505_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i306_4_lut_adj_214_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__24218\,
            in1 => \N__24028\,
            in2 => \N__24202\,
            in3 => \N__36795\,
            lcout => \tok.n174_adj_803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_4_lut_4_lut_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000110"
        )
    port map (
            in0 => \N__31112\,
            in1 => \N__31942\,
            in2 => \N__34796\,
            in3 => \N__33198\,
            lcout => \tok.n867\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i320_4_lut_4_lut_4_lut_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000100010"
        )
    port map (
            in0 => \N__24169\,
            in1 => \N__31885\,
            in2 => \N__37645\,
            in3 => \N__30787\,
            lcout => \tok.n168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6943_3_lut_4_lut_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__36229\,
            in1 => \N__24454\,
            in2 => \N__34096\,
            in3 => \N__29619\,
            lcout => \tok.n6360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i304_4_lut_4_lut_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__26349\,
            in1 => \N__31884\,
            in2 => \N__24061\,
            in3 => \N__30786\,
            lcout => \tok.n210_adj_802\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i10_1_lut_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26758\,
            lcout => \tok.n316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6909_2_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30058\,
            in2 => \_gnd_net_\,
            in3 => \N__34026\,
            lcout => OPEN,
            ltout => \tok.n6409_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i310_4_lut_adj_329_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__30788\,
            in1 => \N__33484\,
            in2 => \N__24004\,
            in3 => \N__23999\,
            lcout => \tok.n215_adj_887\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i309_4_lut_adj_272_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__24604\,
            in1 => \N__36154\,
            in2 => \N__24552\,
            in3 => \N__26768\,
            lcout => \tok.n179_adj_842\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6936_3_lut_4_lut_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__36155\,
            in1 => \N__34070\,
            in2 => \N__30345\,
            in3 => \N__24441\,
            lcout => OPEN,
            ltout => \tok.n6433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6655_4_lut_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__35457\,
            in1 => \N__26933\,
            in2 => \N__24598\,
            in3 => \N__24595\,
            lcout => OPEN,
            ltout => \tok.n6602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6987_4_lut_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__34675\,
            in1 => \N__24583\,
            in2 => \N__24577\,
            in3 => \N__35459\,
            lcout => \tok.n6601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6940_3_lut_4_lut_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__34069\,
            in1 => \N__36153\,
            in2 => \N__24459\,
            in3 => \N__26767\,
            lcout => \tok.n6375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i309_4_lut_adj_47_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__36156\,
            in1 => \N__24343\,
            in2 => \N__24553\,
            in3 => \N__32231\,
            lcout => OPEN,
            ltout => \tok.n179_adj_657_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6980_4_lut_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__35458\,
            in1 => \N__24493\,
            in2 => \N__24487\,
            in3 => \N__34676\,
            lcout => \tok.n6543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i305_3_lut_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30532\,
            in1 => \N__35456\,
            in2 => \_gnd_net_\,
            in3 => \N__31088\,
            lcout => \tok.n464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6874_2_lut_3_lut_4_lut_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__34071\,
            in1 => \N__37127\,
            in2 => \N__24458\,
            in3 => \N__26792\,
            lcout => \tok.n6382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i40_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24801\,
            in1 => \N__24681\,
            in2 => \_gnd_net_\,
            in3 => \N__28692\,
            lcout => tail_40,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38466\,
            ce => \N__28920\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i32_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24706\,
            in1 => \N__24651\,
            in2 => \_gnd_net_\,
            in3 => \N__28691\,
            lcout => \tok.C_stk.tail_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38466\,
            ce => \N__28920\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i48_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28693\,
            in1 => \N__24784\,
            in2 => \_gnd_net_\,
            in3 => \N__24705\,
            lcout => tail_48_adj_900,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38466\,
            ce => \N__28920\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i16_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24652\,
            in1 => \N__24697\,
            in2 => \_gnd_net_\,
            in3 => \N__28689\,
            lcout => \tok.C_stk.tail_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38466\,
            ce => \N__28920\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i24_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24682\,
            in1 => \N__24663\,
            in2 => \_gnd_net_\,
            in3 => \N__28690\,
            lcout => tail_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38466\,
            ce => \N__28920\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i49_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24766\,
            in1 => \N__25186\,
            in2 => \_gnd_net_\,
            in3 => \N__28623\,
            lcout => tail_49_adj_899,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38471\,
            ce => \N__28889\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i51_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24817\,
            in1 => \N__24640\,
            in2 => \_gnd_net_\,
            in3 => \N__28625\,
            lcout => tail_51,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38471\,
            ce => \N__28889\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i54_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28628\,
            in1 => \N__24721\,
            in2 => \_gnd_net_\,
            in3 => \N__28134\,
            lcout => \tok.tail_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38471\,
            ce => \N__28889\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i53_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25012\,
            in1 => \N__24622\,
            in2 => \_gnd_net_\,
            in3 => \N__28627\,
            lcout => \tok.tail_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38471\,
            ce => \N__28889\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i52_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28626\,
            in1 => \N__24733\,
            in2 => \_gnd_net_\,
            in3 => \N__24871\,
            lcout => \tok.tail_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38471\,
            ce => \N__28889\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i50_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24855\,
            in1 => \N__27760\,
            in2 => \_gnd_net_\,
            in3 => \N__28624\,
            lcout => \tok.tail_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38471\,
            ce => \N__28889\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i55_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28629\,
            in1 => \N__28501\,
            in2 => \_gnd_net_\,
            in3 => \N__28939\,
            lcout => \tok.tail_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38471\,
            ce => \N__28889\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i59_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__28607\,
            in1 => \N__24816\,
            in2 => \N__24841\,
            in3 => \N__28834\,
            lcout => tail_59,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i56_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__28832\,
            in1 => \N__24780\,
            in2 => \N__24805\,
            in3 => \N__28606\,
            lcout => tail_56,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2545_2_lut_4_lut_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__25068\,
            in1 => \N__25050\,
            in2 => \N__29838\,
            in3 => \N__25247\,
            lcout => \C_stk_delta_1\,
            ltout => \C_stk_delta_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i57_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__28833\,
            in1 => \N__25209\,
            in2 => \N__24769\,
            in3 => \N__24762\,
            lcout => tail_57,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i60_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__28608\,
            in1 => \N__24732\,
            in2 => \N__24750\,
            in3 => \N__28830\,
            lcout => \tok.tail_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i62_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__28831\,
            in1 => \N__24717\,
            in2 => \N__28159\,
            in3 => \N__28610\,
            lcout => \tok.tail_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i427_2_lut_4_lut_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110110011"
        )
    port map (
            in0 => \N__25069\,
            in1 => \N__25051\,
            in2 => \N__29839\,
            in3 => \N__25248\,
            lcout => \rd_7__N_373\,
            ltout => \rd_7__N_373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i61_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__25029\,
            in1 => \N__25011\,
            in2 => \N__25015\,
            in3 => \N__28609\,
            lcout => \tok.tail_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i1_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28618\,
            in1 => \N__24901\,
            in2 => \_gnd_net_\,
            in3 => \N__24928\,
            lcout => \tok.C_stk.tail_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38480\,
            ce => \N__28873\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i6164_3_lut_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24909\,
            in1 => \N__28117\,
            in2 => \_gnd_net_\,
            in3 => \N__25000\,
            lcout => OPEN,
            ltout => \tok.C_stk.n6248_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i1_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__28053\,
            in1 => \N__27941\,
            in2 => \N__24970\,
            in3 => \N__24967\,
            lcout => c_stk_r_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38480\,
            ce => \N__28873\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i9_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24910\,
            in1 => \_gnd_net_\,
            in2 => \N__24892\,
            in3 => \N__28622\,
            lcout => tail_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38480\,
            ce => \N__28873\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i17_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28617\,
            in1 => \N__24880\,
            in2 => \_gnd_net_\,
            in3 => \N__24900\,
            lcout => \tok.C_stk.tail_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38480\,
            ce => \N__28873\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i25_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24888\,
            in1 => \N__25195\,
            in2 => \_gnd_net_\,
            in3 => \N__28619\,
            lcout => tail_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38480\,
            ce => \N__28873\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i33_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28620\,
            in1 => \N__24879\,
            in2 => \_gnd_net_\,
            in3 => \N__25185\,
            lcout => \tok.C_stk.tail_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38480\,
            ce => \N__28873\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i41_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25210\,
            in1 => \N__25194\,
            in2 => \_gnd_net_\,
            in3 => \N__28621\,
            lcout => tail_41,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38480\,
            ce => \N__28873\,
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_144_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011111100"
        )
    port map (
            in0 => \N__25171\,
            in1 => \N__36318\,
            in2 => \N__34838\,
            in3 => \N__37095\,
            lcout => \tok.n265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_134_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35507\,
            in2 => \_gnd_net_\,
            in3 => \N__33252\,
            lcout => \tok.n156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i338_4_lut_adj_143_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110100000"
        )
    port map (
            in0 => \N__31300\,
            in1 => \N__36319\,
            in2 => \N__33298\,
            in3 => \N__34811\,
            lcout => OPEN,
            ltout => \tok.n211_adj_741_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_3_lut_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110101"
        )
    port map (
            in0 => \N__37096\,
            in1 => \_gnd_net_\,
            in2 => \N__25165\,
            in3 => \N__32133\,
            lcout => OPEN,
            ltout => \tok.n277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_150_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__31301\,
            in1 => \N__35509\,
            in2 => \N__25162\,
            in3 => \N__25159\,
            lcout => \tok.n6_adj_748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i361_4_lut_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__26863\,
            in1 => \N__32132\,
            in2 => \N__25138\,
            in3 => \N__33253\,
            lcout => OPEN,
            ltout => \tok.n238_adj_855_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_295_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__35508\,
            in1 => \N__36317\,
            in2 => \N__25123\,
            in3 => \N__25075\,
            lcout => \tok.n4_adj_859\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_289_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111011101"
        )
    port map (
            in0 => \N__37094\,
            in1 => \N__34781\,
            in2 => \N__25111\,
            in3 => \N__31299\,
            lcout => \tok.n298_adj_856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_i0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__29346\,
            in1 => \_gnd_net_\,
            in2 => \N__29818\,
            in3 => \_gnd_net_\,
            lcout => \tok.depth_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38487\,
            ce => 'H',
            sr => \N__29168\
        );

    \tok.i1_2_lut_adj_288_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29814\,
            in2 => \_gnd_net_\,
            in3 => \N__29345\,
            lcout => OPEN,
            ltout => \tok.n53_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7015_4_lut_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__25378\,
            in1 => \N__25409\,
            in2 => \N__25654\,
            in3 => \N__29305\,
            lcout => \tok.n992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_3__I_0_389_i2_2_lut_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29759\,
            in2 => \_gnd_net_\,
            in3 => \N__28979\,
            lcout => OPEN,
            ltout => \tok.n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_287_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31312\,
            in1 => \N__26500\,
            in2 => \N__25522\,
            in3 => \N__25216\,
            lcout => \tok.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2566_2_lut_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29344\,
            in2 => \_gnd_net_\,
            in3 => \N__29395\,
            lcout => \tok.n174\,
            ltout => \tok.n174_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_i2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__28980\,
            in1 => \_gnd_net_\,
            in2 => \N__25381\,
            in3 => \N__29287\,
            lcout => \tok.depth_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38487\,
            ce => 'H',
            sr => \N__29168\
        );

    \tok.i6106_2_lut_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25377\,
            in2 => \_gnd_net_\,
            in3 => \N__29396\,
            lcout => \tok.n6189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_adj_118_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__37087\,
            in1 => \N__35506\,
            in2 => \N__29851\,
            in3 => \N__36301\,
            lcout => \tok.n6_adj_722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i965_3_lut_3_lut_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101100110"
        )
    port map (
            in0 => \N__36300\,
            in1 => \N__32092\,
            in2 => \_gnd_net_\,
            in3 => \N__33249\,
            lcout => OPEN,
            ltout => \tok.n10_adj_773_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_174_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__33250\,
            in1 => \N__25828\,
            in2 => \N__25819\,
            in3 => \N__31307\,
            lcout => OPEN,
            ltout => \tok.n6146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_178_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__25660\,
            in1 => \N__28973\,
            in2 => \N__25816\,
            in3 => \N__37086\,
            lcout => \tok.n86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i349_4_lut_4_lut_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010100000101"
        )
    port map (
            in0 => \N__33251\,
            in1 => \N__36302\,
            in2 => \N__37128\,
            in3 => \N__31308\,
            lcout => OPEN,
            ltout => \tok.n369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_109_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__31309\,
            in1 => \N__25738\,
            in2 => \N__25705\,
            in3 => \N__34812\,
            lcout => OPEN,
            ltout => \tok.n233_adj_716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_114_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__32093\,
            in1 => \N__25702\,
            in2 => \N__25690\,
            in3 => \N__25687\,
            lcout => \tok.n6156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_adj_177_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29847\,
            in2 => \_gnd_net_\,
            in3 => \N__29757\,
            lcout => \tok.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6858_4_lut_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__26496\,
            in1 => \N__26842\,
            in2 => \N__26074\,
            in3 => \N__31314\,
            lcout => \tok.n6639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6753_2_lut_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28189\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32115\,
            lcout => OPEN,
            ltout => \tok.n6653_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6982_4_lut_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010100000"
        )
    port map (
            in0 => \N__26130\,
            in1 => \N__26098\,
            in2 => \N__26080\,
            in3 => \N__34809\,
            lcout => OPEN,
            ltout => \tok.n6646_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i341_4_lut_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__35514\,
            in1 => \N__27091\,
            in2 => \N__26077\,
            in3 => \N__33190\,
            lcout => \tok.n280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_221_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34808\,
            in2 => \_gnd_net_\,
            in3 => \N__35510\,
            lcout => \tok.n6167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6989_4_lut_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__31315\,
            in1 => \N__26065\,
            in2 => \N__26053\,
            in3 => \N__33191\,
            lcout => OPEN,
            ltout => \tok.n6638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6963_4_lut_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__26038\,
            in1 => \N__26032\,
            in2 => \N__26026\,
            in3 => \N__37068\,
            lcout => \tok.n6636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i345_3_lut_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31313\,
            in2 => \N__35524\,
            in3 => \N__26014\,
            lcout => \tok.n367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i317_4_lut_adj_210_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110100000"
        )
    port map (
            in0 => \N__36988\,
            in1 => \N__30026\,
            in2 => \N__25992\,
            in3 => \N__31188\,
            lcout => OPEN,
            ltout => \tok.n177_adj_799_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i303_4_lut_adj_213_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__25882\,
            in1 => \N__25840\,
            in2 => \N__25831\,
            in3 => \N__35485\,
            lcout => OPEN,
            ltout => \tok.n252_adj_801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_215_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__35486\,
            in1 => \N__26266\,
            in2 => \N__26395\,
            in3 => \N__34816\,
            lcout => \tok.n4_adj_804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_223_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__34815\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36986\,
            lcout => \tok.n5_adj_745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i314_4_lut_adj_198_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__36987\,
            in1 => \N__26445\,
            in2 => \N__26391\,
            in3 => \N__26350\,
            lcout => OPEN,
            ltout => \tok.n255_adj_793_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_212_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__26446\,
            in1 => \N__26287\,
            in2 => \N__26269\,
            in3 => \N__36258\,
            lcout => \tok.n258_adj_800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_263_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000001000"
        )
    port map (
            in0 => \N__36985\,
            in1 => \N__34814\,
            in2 => \N__29412\,
            in3 => \N__31187\,
            lcout => OPEN,
            ltout => \tok.n6162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_264_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__26483\,
            in1 => \N__26259\,
            in2 => \N__26236\,
            in3 => \N__36257\,
            lcout => \tok.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__34094\,
            in1 => \N__35488\,
            in2 => \N__32594\,
            in3 => \N__27536\,
            lcout => OPEN,
            ltout => \tok.n865_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6776_4_lut_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101000"
        )
    port map (
            in0 => \N__32547\,
            in1 => \N__30027\,
            in2 => \N__26233\,
            in3 => \N__32585\,
            lcout => \tok.n6496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_3_lut_adj_260_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__36259\,
            in1 => \N__34817\,
            in2 => \_gnd_net_\,
            in3 => \N__33257\,
            lcout => \tok.n222\,
            ltout => \tok.n222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i11_3_lut_4_lut_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011111100"
        )
    port map (
            in0 => \N__34818\,
            in1 => \N__27083\,
            in2 => \N__26230\,
            in3 => \N__36260\,
            lcout => \tok.n245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_208_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__36261\,
            in1 => \N__29890\,
            in2 => \N__26641\,
            in3 => \N__33258\,
            lcout => OPEN,
            ltout => \tok.n186_adj_798_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i315_4_lut_adj_216_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__34819\,
            in1 => \N__35489\,
            in2 => \N__26629\,
            in3 => \N__26626\,
            lcout => OPEN,
            ltout => \tok.n338_adj_805_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6759_4_lut_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__30028\,
            in1 => \N__26608\,
            in2 => \N__26530\,
            in3 => \N__26416\,
            lcout => \tok.n6608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_286_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37043\,
            in2 => \_gnd_net_\,
            in3 => \N__31229\,
            lcout => \tok.n4_adj_712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_36_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31744\,
            in2 => \_gnd_net_\,
            in3 => \N__33102\,
            lcout => \tok.n219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_adj_256_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__31745\,
            in1 => \N__31225\,
            in2 => \N__27558\,
            in3 => \N__35481\,
            lcout => \tok.n190_adj_792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_217_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000100"
        )
    port map (
            in0 => \N__34078\,
            in1 => \N__26434\,
            in2 => \N__33299\,
            in3 => \N__26425\,
            lcout => \tok.n205_adj_806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i317_4_lut_adj_233_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110100000"
        )
    port map (
            in0 => \N__28338\,
            in1 => \N__37455\,
            in2 => \N__36936\,
            in3 => \N__31226\,
            lcout => \tok.n177_adj_813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_220_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__33259\,
            in1 => \_gnd_net_\,
            in2 => \N__31957\,
            in3 => \N__36784\,
            lcout => \tok.n821\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2575_2_lut_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34077\,
            in2 => \_gnd_net_\,
            in3 => \N__37456\,
            lcout => OPEN,
            ltout => \tok.n2598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i310_4_lut_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__31227\,
            in1 => \N__33467\,
            in2 => \N__27046\,
            in3 => \N__27037\,
            lcout => OPEN,
            ltout => \tok.n215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6831_4_lut_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__26947\,
            in1 => \N__26906\,
            in2 => \N__26878\,
            in3 => \N__35482\,
            lcout => \tok.n6547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6966_2_lut_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26856\,
            in2 => \_gnd_net_\,
            in3 => \N__26838\,
            lcout => OPEN,
            ltout => \tok.n6650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i337_4_lut_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__35356\,
            in1 => \N__27609\,
            in2 => \N__26806\,
            in3 => \N__26779\,
            lcout => OPEN,
            ltout => \tok.n211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6969_3_lut_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34698\,
            in2 => \N__26671\,
            in3 => \N__34053\,
            lcout => \tok.n6641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_105_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010100"
        )
    port map (
            in0 => \N__35357\,
            in1 => \N__34699\,
            in2 => \N__26668\,
            in3 => \N__33233\,
            lcout => OPEN,
            ltout => \tok.n260_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_106_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110010"
        )
    port map (
            in0 => \N__34700\,
            in1 => \N__37067\,
            in2 => \N__26644\,
            in3 => \N__27540\,
            lcout => OPEN,
            ltout => \tok.n266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_115_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111100"
        )
    port map (
            in0 => \N__27400\,
            in1 => \N__27619\,
            in2 => \N__27613\,
            in3 => \N__36177\,
            lcout => OPEN,
            ltout => \tok.n4_adj_718_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_318_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__27610\,
            in1 => \N__27592\,
            in2 => \N__27580\,
            in3 => \N__32078\,
            lcout => \tok.n221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i344_4_lut_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__34052\,
            in1 => \N__37066\,
            in2 => \N__27559\,
            in3 => \N__33232\,
            lcout => \tok.n2637\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i7_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37534\,
            in1 => \N__27190\,
            in2 => \_gnd_net_\,
            in3 => \N__27382\,
            lcout => \tok.uart.sender_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38506\,
            ce => \N__27178\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i8_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27184\,
            in1 => \N__37535\,
            in2 => \_gnd_net_\,
            in3 => \N__30346\,
            lcout => \tok.uart.sender_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38506\,
            ce => \N__27178\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i9_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37536\,
            in1 => \N__37299\,
            in2 => \_gnd_net_\,
            in3 => \N__30062\,
            lcout => \tok.uart.sender_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38506\,
            ce => \N__27178\,
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_126_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34764\,
            in2 => \_gnd_net_\,
            in3 => \N__33124\,
            lcout => \tok.n274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_68_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32079\,
            in2 => \_gnd_net_\,
            in3 => \N__31228\,
            lcout => \tok.n185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_rep_284_2_lut_2_lut_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36282\,
            in2 => \_gnd_net_\,
            in3 => \N__32080\,
            lcout => \tok.n7410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.reset_I_0_1_lut_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27787\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.reset_N_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i58_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__27759\,
            in1 => \N__28835\,
            in2 => \N__27777\,
            in3 => \N__28674\,
            lcout => \tok.tail_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i6_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28616\,
            in1 => \N__27649\,
            in2 => \_gnd_net_\,
            in3 => \N__27672\,
            lcout => \tok.C_stk.tail_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38481\,
            ce => \N__28910\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i6149_3_lut_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27657\,
            in1 => \N__28123\,
            in2 => \_gnd_net_\,
            in3 => \N__27748\,
            lcout => OPEN,
            ltout => \tok.C_stk.n6233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i6_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__28048\,
            in1 => \N__27943\,
            in2 => \N__27718\,
            in3 => \N__27715\,
            lcout => \tok.c_stk_r_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38481\,
            ce => \N__28910\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i14_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27658\,
            in1 => \_gnd_net_\,
            in2 => \N__27640\,
            in3 => \N__28611\,
            lcout => \tok.tail_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38481\,
            ce => \N__28910\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i22_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28612\,
            in1 => \N__27628\,
            in2 => \_gnd_net_\,
            in3 => \N__27648\,
            lcout => \tok.C_stk.tail_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38481\,
            ce => \N__28910\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i30_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27636\,
            in1 => \N__28144\,
            in2 => \_gnd_net_\,
            in3 => \N__28613\,
            lcout => \tok.tail_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38481\,
            ce => \N__28910\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i38_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28614\,
            in1 => \N__28135\,
            in2 => \_gnd_net_\,
            in3 => \N__27627\,
            lcout => \tok.C_stk.tail_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38481\,
            ce => \N__28910\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i46_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28158\,
            in1 => \N__28143\,
            in2 => \_gnd_net_\,
            in3 => \N__28615\,
            lcout => \tok.tail_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38481\,
            ce => \N__28910\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i7_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28665\,
            in1 => \N__27826\,
            in2 => \_gnd_net_\,
            in3 => \N__27853\,
            lcout => \tok.C_stk.tail_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38484\,
            ce => \N__28917\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i6143_3_lut_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27834\,
            in1 => \N__28118\,
            in2 => \_gnd_net_\,
            in3 => \N__28380\,
            lcout => OPEN,
            ltout => \tok.C_stk.n6227_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i7_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__28052\,
            in1 => \N__27978\,
            in2 => \N__27946\,
            in3 => \N__27942\,
            lcout => \tok.c_stk_r_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38484\,
            ce => \N__28917\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i15_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27835\,
            in1 => \_gnd_net_\,
            in2 => \N__27817\,
            in3 => \N__28660\,
            lcout => \tok.tail_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38484\,
            ce => \N__28917\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i23_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28661\,
            in1 => \N__27805\,
            in2 => \_gnd_net_\,
            in3 => \N__27825\,
            lcout => \tok.C_stk.tail_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38484\,
            ce => \N__28917\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i31_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27813\,
            in1 => \N__27796\,
            in2 => \_gnd_net_\,
            in3 => \N__28662\,
            lcout => \tok.tail_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38484\,
            ce => \N__28917\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i39_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28663\,
            in1 => \N__28935\,
            in2 => \_gnd_net_\,
            in3 => \N__27804\,
            lcout => \tok.C_stk.tail_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38484\,
            ce => \N__28917\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i47_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28776\,
            in1 => \N__27795\,
            in2 => \_gnd_net_\,
            in3 => \N__28664\,
            lcout => \tok.tail_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38484\,
            ce => \N__28917\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i63_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__28862\,
            in1 => \N__28494\,
            in2 => \N__28780\,
            in3 => \N__28735\,
            lcout => \tok.tail_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i1608_3_lut_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28472\,
            in1 => \N__28381\,
            in2 => \_gnd_net_\,
            in3 => \N__28339\,
            lcout => \tok.table_wr_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i1_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28174\,
            in1 => \N__37808\,
            in2 => \_gnd_net_\,
            in3 => \N__38217\,
            lcout => capture_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37270\,
            in1 => \N__37790\,
            in2 => \_gnd_net_\,
            in3 => \N__28221\,
            lcout => uart_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i2_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37789\,
            in1 => \_gnd_net_\,
            in2 => \N__37288\,
            in3 => \N__28203\,
            lcout => uart_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i1_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28173\,
            in1 => \N__37788\,
            in2 => \_gnd_net_\,
            in3 => \N__28188\,
            lcout => uart_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i2_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37284\,
            in1 => \N__28172\,
            in2 => \_gnd_net_\,
            in3 => \N__38218\,
            lcout => capture_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_87_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100101101100"
        )
    port map (
            in0 => \N__29285\,
            in1 => \N__29753\,
            in2 => \N__28981\,
            in3 => \N__29297\,
            lcout => \tok.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_i1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001111101100000"
        )
    port map (
            in0 => \N__29401\,
            in1 => \N__29798\,
            in2 => \N__29359\,
            in3 => \N__29873\,
            lcout => \tok.depth_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38492\,
            ce => 'H',
            sr => \N__29116\
        );

    \tok.i2_4_lut_4_lut_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011001101010"
        )
    port map (
            in0 => \N__29872\,
            in1 => \N__29355\,
            in2 => \N__29811\,
            in3 => \N__29400\,
            lcout => \tok.n52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_adj_72_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28971\,
            in1 => \N__29794\,
            in2 => \N__29760\,
            in3 => \N__29870\,
            lcout => \tok.A_stk_delta_1__N_4\,
            ltout => \tok.A_stk_delta_1__N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_252_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__29871\,
            in1 => \N__29813\,
            in2 => \N__29362\,
            in3 => \N__29354\,
            lcout => \tok.n4_adj_702\,
            ltout => \tok.n4_adj_702_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__29298\,
            in1 => \_gnd_net_\,
            in2 => \N__29323\,
            in3 => \N__28977\,
            lcout => OPEN,
            ltout => \tok.n51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29320\,
            in2 => \N__29314\,
            in3 => \N__29311\,
            lcout => \tok.n8_adj_854\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_i3_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011010011010010"
        )
    port map (
            in0 => \N__29299\,
            in1 => \N__29286\,
            in2 => \N__29761\,
            in3 => \N__28978\,
            lcout => \tok.depth_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38492\,
            ce => 'H',
            sr => \N__29116\
        );

    \tok.i1_4_lut_adj_151_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__29008\,
            in1 => \N__28999\,
            in2 => \N__32134\,
            in3 => \N__34763\,
            lcout => \tok.n215_adj_750\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6129_2_lut_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28972\,
            in2 => \_gnd_net_\,
            in3 => \N__29875\,
            lcout => \tok.n6213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_4_lut_adj_335_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__29874\,
            in1 => \N__34108\,
            in2 => \N__29812\,
            in3 => \N__34760\,
            lcout => \tok.n741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_199_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__34761\,
            in1 => \_gnd_net_\,
            in2 => \N__34114\,
            in3 => \N__37084\,
            lcout => \tok.n806\,
            ltout => \tok.n806_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_173_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__29802\,
            in1 => \N__29770\,
            in2 => \N__29764\,
            in3 => \N__29758\,
            lcout => \tok.n748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i299_4_lut_adj_119_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__34762\,
            in1 => \N__29626\,
            in2 => \N__29476\,
            in3 => \N__31310\,
            lcout => OPEN,
            ltout => \tok.n158_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6851_3_lut_4_lut_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__37085\,
            in1 => \N__32127\,
            in2 => \N__29461\,
            in3 => \N__33280\,
            lcout => \tok.n6627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i8_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38208\,
            in1 => \N__37661\,
            in2 => \_gnd_net_\,
            in3 => \N__37870\,
            lcout => capture_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__29428\,
            in1 => \N__37720\,
            in2 => \N__29422\,
            in3 => \N__30146\,
            lcout => \tok.uart_stall_N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_373_i9_2_lut_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33244\,
            in2 => \_gnd_net_\,
            in3 => \N__30937\,
            lcout => \tok.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_i10_2_lut_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34807\,
            in2 => \_gnd_net_\,
            in3 => \N__32113\,
            lcout => \tok.n10\,
            ltout => \tok.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7025_2_lut_3_lut_4_lut_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__30148\,
            in1 => \N__33248\,
            in2 => \N__30172\,
            in3 => \N__30939\,
            lcout => \tok.write_flag\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i4_4_lut_adj_21_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__30938\,
            in1 => \N__37721\,
            in2 => \N__33297\,
            in3 => \N__30147\,
            lcout => OPEN,
            ltout => \tok.uart.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i7042_3_lut_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__32114\,
            in1 => \_gnd_net_\,
            in2 => \N__30094\,
            in3 => \N__34810\,
            lcout => n23,
            ltout => \n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i7022_2_lut_3_lut_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37616\,
            in2 => \N__30091\,
            in3 => \N__37722\,
            lcout => \tok.uart.n1013\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_3_lut_adj_25_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__37723\,
            in1 => \_gnd_net_\,
            in2 => \N__37623\,
            in3 => \N__37500\,
            lcout => \tok.uart.n994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i320_4_lut_4_lut_4_lut_adj_102_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010110000000"
        )
    port map (
            in0 => \N__31305\,
            in1 => \N__29883\,
            in2 => \N__32131\,
            in3 => \N__32378\,
            lcout => OPEN,
            ltout => \tok.n168_adj_710_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6945_4_lut_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__32476\,
            in1 => \N__36364\,
            in2 => \N__30088\,
            in3 => \N__30064\,
            lcout => \tok.n6502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i6_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37791\,
            in1 => \N__37152\,
            in2 => \_gnd_net_\,
            in3 => \N__29884\,
            lcout => uart_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i7_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37151\,
            in1 => \N__37668\,
            in2 => \_gnd_net_\,
            in3 => \N__38184\,
            lcout => capture_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_105_i15_1_lut_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32377\,
            lcout => \tok.n311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_adj_204_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001001000"
        )
    port map (
            in0 => \N__33607\,
            in1 => \N__32087\,
            in2 => \N__34112\,
            in3 => \N__31304\,
            lcout => \tok.n190_adj_797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i320_4_lut_4_lut_4_lut_adj_75_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000100010"
        )
    port map (
            in0 => \N__32230\,
            in1 => \N__32091\,
            in2 => \N__37834\,
            in3 => \N__31306\,
            lcout => \tok.n168_adj_690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6949_4_lut_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__32470\,
            in1 => \N__36374\,
            in2 => \N__30577\,
            in3 => \N__30314\,
            lcout => OPEN,
            ltout => \tok.n6526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_180_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__30568\,
            in1 => \N__36269\,
            in2 => \N__30553\,
            in3 => \N__33294\,
            lcout => OPEN,
            ltout => \tok.n186_adj_777_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i315_4_lut_adj_190_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__30178\,
            in1 => \N__35487\,
            in2 => \N__30550\,
            in3 => \N__34779\,
            lcout => \tok.n338_adj_787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_adj_61_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__30525\,
            in1 => \N__34095\,
            in2 => \N__32593\,
            in3 => \N__37044\,
            lcout => OPEN,
            ltout => \tok.n866_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6793_4_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__30313\,
            in1 => \N__32549\,
            in2 => \N__30181\,
            in3 => \N__32581\,
            lcout => \tok.n6520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i271_2_lut_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35951\,
            in2 => \_gnd_net_\,
            in3 => \N__36753\,
            lcout => \tok.n317\,
            ltout => \tok.n317_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_98_i8_3_lut_4_lut_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101001"
        )
    port map (
            in0 => \N__34092\,
            in1 => \N__35483\,
            in2 => \N__36559\,
            in3 => \N__36549\,
            lcout => \tok.n205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6934_4_lut_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__36388\,
            in1 => \N__32472\,
            in2 => \N__36376\,
            in3 => \N__37476\,
            lcout => OPEN,
            ltout => \tok.n6478_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i308_4_lut_adj_232_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__35952\,
            in1 => \N__32386\,
            in2 => \N__35527\,
            in3 => \N__33293\,
            lcout => OPEN,
            ltout => \tok.n186_adj_812_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i315_4_lut_adj_241_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__35484\,
            in1 => \N__32482\,
            in2 => \N__34849\,
            in3 => \N__34778\,
            lcout => \tok.n338_adj_819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_4_lut_adj_290_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__34093\,
            in1 => \N__33644\,
            in2 => \N__33483\,
            in3 => \N__33292\,
            lcout => OPEN,
            ltout => \tok.n863_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6758_4_lut_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__32586\,
            in1 => \N__32548\,
            in2 => \N__32485\,
            in3 => \N__37475\,
            lcout => \tok.n6472\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6760_2_lut_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32471\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32400\,
            lcout => \tok.n6477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i7_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37669\,
            in1 => \N__37795\,
            in2 => \_gnd_net_\,
            in3 => \N__37641\,
            lcout => uart_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i10_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__37627\,
            in1 => \N__37515\,
            in2 => \N__37303\,
            in3 => \N__37474\,
            lcout => sender_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i3_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37911\,
            in1 => \N__37283\,
            in2 => \_gnd_net_\,
            in3 => \N__38214\,
            lcout => capture_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_3_lut_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__37787\,
            in1 => \N__37190\,
            in2 => \_gnd_net_\,
            in3 => \N__37242\,
            lcout => \tok.uart.n922\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i4_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37266\,
            in1 => \N__37910\,
            in2 => \_gnd_net_\,
            in3 => \N__38215\,
            lcout => capture_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i5_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__38216\,
            in1 => \N__37855\,
            in2 => \_gnd_net_\,
            in3 => \N__37265\,
            lcout => capture_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.valid_54_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37191\,
            in2 => \_gnd_net_\,
            in3 => \N__37252\,
            lcout => \tok.uart_rx_valid\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38498\,
            ce => \N__37171\,
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i6_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38206\,
            in1 => \N__37847\,
            in2 => \_gnd_net_\,
            in3 => \N__37159\,
            lcout => capture_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i0_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37815\,
            in1 => \N__37924\,
            in2 => \_gnd_net_\,
            in3 => \N__38205\,
            lcout => capture_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i2_3_lut_adj_24_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__37923\,
            in1 => \N__37868\,
            in2 => \_gnd_net_\,
            in3 => \N__37984\,
            lcout => \rx_data_7__N_510\,
            ltout => \rx_data_7__N_510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i3_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37915\,
            in2 => \N__37894\,
            in3 => \N__37884\,
            lcout => uart_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i9_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__38207\,
            in1 => \N__38010\,
            in2 => \_gnd_net_\,
            in3 => \N__37869\,
            lcout => capture_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i5_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37780\,
            in1 => \_gnd_net_\,
            in2 => \N__37854\,
            in3 => \N__37830\,
            lcout => uart_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i0_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37816\,
            in1 => \N__37779\,
            in2 => \_gnd_net_\,
            in3 => \N__37737\,
            lcout => uart_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i2_4_lut_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__37707\,
            in1 => \N__38046\,
            in2 => \N__37699\,
            in3 => \N__37681\,
            lcout => \tok.uart_tx_busy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sentbits_143__i3_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__37684\,
            in1 => \N__37698\,
            in2 => \N__38056\,
            in3 => \N__37708\,
            lcout => \tok.uart.sentbits_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38504\,
            ce => \N__38032\,
            sr => \N__38020\
        );

    \tok.uart.sentbits_143__i2_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__37697\,
            in1 => \N__38051\,
            in2 => \_gnd_net_\,
            in3 => \N__37683\,
            lcout => \tok.uart.sentbits_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38504\,
            ce => \N__38032\,
            sr => \N__38020\
        );

    \tok.uart.sentbits_143__i1_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__37682\,
            in1 => \_gnd_net_\,
            in2 => \N__38055\,
            in3 => \_gnd_net_\,
            lcout => \tok.uart.sentbits_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38504\,
            ce => \N__38032\,
            sr => \N__38020\
        );

    \tok.uart.sentbits_143__i0_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38047\,
            lcout => \tok.uart.sentbits_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38504\,
            ce => \N__38032\,
            sr => \N__38020\
        );

    \tok.uart.i3_4_lut_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__38232\,
            in1 => \N__37962\,
            in2 => \N__38011\,
            in3 => \N__37941\,
            lcout => \tok.uart.n809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i3_4_lut_adj_23_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__37940\,
            in1 => \N__38231\,
            in2 => \N__37966\,
            in3 => \N__38629\,
            lcout => \tok.uart.n4977\,
            ltout => \tok.uart.n4977_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rxstop_I_0_60_4_lut_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__38115\,
            in1 => \N__38128\,
            in2 => \N__37978\,
            in3 => \N__38652\,
            lcout => \bytephase_5__N_509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.bytephase__i0_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38076\,
            in2 => \_gnd_net_\,
            in3 => \N__37975\,
            lcout => \tok.uart.bytephase_0\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \tok.uart.n4819\,
            clk => \N__38505\,
            ce => \N__38140\,
            sr => \N__38158\
        );

    \tok.uart.bytephase__i1_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38653\,
            in2 => \_gnd_net_\,
            in3 => \N__37972\,
            lcout => \tok.uart.bytephase_1\,
            ltout => OPEN,
            carryin => \tok.uart.n4819\,
            carryout => \tok.uart.n4820\,
            clk => \N__38505\,
            ce => \N__38140\,
            sr => \N__38158\
        );

    \tok.uart.bytephase__i2_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38092\,
            in2 => \_gnd_net_\,
            in3 => \N__37969\,
            lcout => \tok.uart.bytephase_2\,
            ltout => OPEN,
            carryin => \tok.uart.n4820\,
            carryout => \tok.uart.n4821\,
            clk => \N__38505\,
            ce => \N__38140\,
            sr => \N__38158\
        );

    \tok.uart.bytephase__i3_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37961\,
            in2 => \_gnd_net_\,
            in3 => \N__37945\,
            lcout => \tok.uart.bytephase_3\,
            ltout => OPEN,
            carryin => \tok.uart.n4821\,
            carryout => \tok.uart.n4822\,
            clk => \N__38505\,
            ce => \N__38140\,
            sr => \N__38158\
        );

    \tok.uart.bytephase__i4_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37942\,
            in2 => \_gnd_net_\,
            in3 => \N__37927\,
            lcout => \tok.uart.bytephase_4\,
            ltout => OPEN,
            carryin => \tok.uart.n4822\,
            carryout => \tok.uart.n4823\,
            clk => \N__38505\,
            ce => \N__38140\,
            sr => \N__38158\
        );

    \tok.uart.bytephase__i5_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38233\,
            in2 => \_gnd_net_\,
            in3 => \N__38236\,
            lcout => \tok.uart.bytephase_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38505\,
            ce => \N__38140\,
            sr => \N__38158\
        );

    \tok.uart.i2_3_lut_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__38650\,
            in1 => \_gnd_net_\,
            in2 => \N__38077\,
            in3 => \N__38100\,
            lcout => n4928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__38520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38571\,
            lcout => OPEN,
            ltout => \tok.uart.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i4_4_lut_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__38605\,
            in1 => \N__38619\,
            in2 => \N__38164\,
            in3 => \N__38134\,
            lcout => n746,
            ltout => \n746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38161\,
            in3 => \N__38157\,
            lcout => n974,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i6127_3_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__38586\,
            in1 => \_gnd_net_\,
            in2 => \N__38557\,
            in3 => \N__38538\,
            lcout => \tok.uart.n6211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_adj_22_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__38091\,
            in1 => \N__38072\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tok.uart.n2356\,
            ltout => \tok.uart.n2356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rxrst_I_0_3_lut_4_lut_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011111111"
        )
    port map (
            in0 => \N__38651\,
            in1 => \N__38119\,
            in2 => \N__38104\,
            in3 => \N__38101\,
            lcout => \tok.uart.rxclkcounter_6__N_476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_3_lut_adj_20_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__38090\,
            in1 => \N__38071\,
            in2 => \_gnd_net_\,
            in3 => \N__38649\,
            lcout => \tok.uart.n2357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rxclkcounter_144__i0_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38620\,
            in2 => \_gnd_net_\,
            in3 => \N__38608\,
            lcout => \tok.uart.rxclkcounter_0\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \tok.uart.n4824\,
            clk => \N__38508\,
            ce => 'H',
            sr => \N__38251\
        );

    \tok.uart.rxclkcounter_144__i1_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38604\,
            in2 => \_gnd_net_\,
            in3 => \N__38590\,
            lcout => \tok.uart.rxclkcounter_1\,
            ltout => OPEN,
            carryin => \tok.uart.n4824\,
            carryout => \tok.uart.n4825\,
            clk => \N__38508\,
            ce => 'H',
            sr => \N__38251\
        );

    \tok.uart.rxclkcounter_144__i2_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38587\,
            in2 => \_gnd_net_\,
            in3 => \N__38575\,
            lcout => \tok.uart.rxclkcounter_2\,
            ltout => OPEN,
            carryin => \tok.uart.n4825\,
            carryout => \tok.uart.n4826\,
            clk => \N__38508\,
            ce => 'H',
            sr => \N__38251\
        );

    \tok.uart.rxclkcounter_144__i3_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38572\,
            in2 => \_gnd_net_\,
            in3 => \N__38560\,
            lcout => \tok.uart.rxclkcounter_3\,
            ltout => OPEN,
            carryin => \tok.uart.n4826\,
            carryout => \tok.uart.n4827\,
            clk => \N__38508\,
            ce => 'H',
            sr => \N__38251\
        );

    \tok.uart.rxclkcounter_144__i4_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38556\,
            in2 => \_gnd_net_\,
            in3 => \N__38542\,
            lcout => \tok.uart.rxclkcounter_4\,
            ltout => OPEN,
            carryin => \tok.uart.n4827\,
            carryout => \tok.uart.n4828\,
            clk => \N__38508\,
            ce => 'H',
            sr => \N__38251\
        );

    \tok.uart.rxclkcounter_144__i5_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38539\,
            in2 => \_gnd_net_\,
            in3 => \N__38527\,
            lcout => \tok.uart.rxclkcounter_5\,
            ltout => OPEN,
            carryin => \tok.uart.n4828\,
            carryout => \tok.uart.n4829\,
            clk => \N__38508\,
            ce => 'H',
            sr => \N__38251\
        );

    \tok.uart.rxclkcounter_144__i6_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38521\,
            in2 => \_gnd_net_\,
            in3 => \N__38524\,
            lcout => \tok.uart.rxclkcounter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38508\,
            ce => 'H',
            sr => \N__38251\
        );
end \INTERFACE\;
