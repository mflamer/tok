// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Dec 31 2020 17:42:06

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    tx,
    rx,
    reset);

    output tx;
    input rx;
    input reset;

    wire N__38690;
    wire N__38689;
    wire N__38688;
    wire N__38681;
    wire N__38680;
    wire N__38679;
    wire N__38672;
    wire N__38671;
    wire N__38670;
    wire N__38653;
    wire N__38652;
    wire N__38651;
    wire N__38650;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38636;
    wire N__38629;
    wire N__38626;
    wire N__38623;
    wire N__38620;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38608;
    wire N__38605;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38590;
    wire N__38587;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38575;
    wire N__38572;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38560;
    wire N__38557;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38542;
    wire N__38539;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38520;
    wire N__38517;
    wire N__38514;
    wire N__38509;
    wire N__38508;
    wire N__38507;
    wire N__38506;
    wire N__38505;
    wire N__38504;
    wire N__38503;
    wire N__38502;
    wire N__38501;
    wire N__38500;
    wire N__38499;
    wire N__38498;
    wire N__38497;
    wire N__38496;
    wire N__38495;
    wire N__38494;
    wire N__38493;
    wire N__38492;
    wire N__38491;
    wire N__38490;
    wire N__38489;
    wire N__38488;
    wire N__38487;
    wire N__38486;
    wire N__38485;
    wire N__38484;
    wire N__38483;
    wire N__38482;
    wire N__38481;
    wire N__38480;
    wire N__38479;
    wire N__38478;
    wire N__38477;
    wire N__38476;
    wire N__38475;
    wire N__38474;
    wire N__38473;
    wire N__38472;
    wire N__38471;
    wire N__38470;
    wire N__38469;
    wire N__38468;
    wire N__38467;
    wire N__38466;
    wire N__38465;
    wire N__38464;
    wire N__38463;
    wire N__38462;
    wire N__38461;
    wire N__38460;
    wire N__38459;
    wire N__38458;
    wire N__38457;
    wire N__38456;
    wire N__38455;
    wire N__38454;
    wire N__38453;
    wire N__38452;
    wire N__38451;
    wire N__38450;
    wire N__38449;
    wire N__38448;
    wire N__38447;
    wire N__38446;
    wire N__38445;
    wire N__38444;
    wire N__38443;
    wire N__38442;
    wire N__38441;
    wire N__38440;
    wire N__38439;
    wire N__38438;
    wire N__38437;
    wire N__38436;
    wire N__38435;
    wire N__38434;
    wire N__38433;
    wire N__38432;
    wire N__38431;
    wire N__38430;
    wire N__38429;
    wire N__38428;
    wire N__38427;
    wire N__38426;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38232;
    wire N__38231;
    wire N__38228;
    wire N__38223;
    wire N__38218;
    wire N__38217;
    wire N__38216;
    wire N__38215;
    wire N__38214;
    wire N__38209;
    wire N__38208;
    wire N__38207;
    wire N__38206;
    wire N__38205;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38185;
    wire N__38184;
    wire N__38181;
    wire N__38174;
    wire N__38171;
    wire N__38164;
    wire N__38161;
    wire N__38158;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38145;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38104;
    wire N__38101;
    wire N__38100;
    wire N__38095;
    wire N__38092;
    wire N__38091;
    wire N__38090;
    wire N__38087;
    wire N__38082;
    wire N__38077;
    wire N__38076;
    wire N__38073;
    wire N__38072;
    wire N__38071;
    wire N__38068;
    wire N__38061;
    wire N__38056;
    wire N__38055;
    wire N__38052;
    wire N__38051;
    wire N__38048;
    wire N__38047;
    wire N__38046;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37981;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37962;
    wire N__37961;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37945;
    wire N__37942;
    wire N__37941;
    wire N__37940;
    wire N__37937;
    wire N__37932;
    wire N__37927;
    wire N__37924;
    wire N__37923;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37911;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37870;
    wire N__37869;
    wire N__37868;
    wire N__37865;
    wire N__37860;
    wire N__37855;
    wire N__37854;
    wire N__37851;
    wire N__37848;
    wire N__37847;
    wire N__37844;
    wire N__37839;
    wire N__37834;
    wire N__37831;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37816;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37808;
    wire N__37803;
    wire N__37800;
    wire N__37795;
    wire N__37792;
    wire N__37791;
    wire N__37790;
    wire N__37789;
    wire N__37788;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37780;
    wire N__37779;
    wire N__37772;
    wire N__37769;
    wire N__37764;
    wire N__37759;
    wire N__37754;
    wire N__37747;
    wire N__37744;
    wire N__37741;
    wire N__37738;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37723;
    wire N__37722;
    wire N__37721;
    wire N__37720;
    wire N__37711;
    wire N__37708;
    wire N__37707;
    wire N__37702;
    wire N__37699;
    wire N__37698;
    wire N__37697;
    wire N__37694;
    wire N__37687;
    wire N__37684;
    wire N__37683;
    wire N__37682;
    wire N__37681;
    wire N__37672;
    wire N__37669;
    wire N__37668;
    wire N__37665;
    wire N__37662;
    wire N__37661;
    wire N__37658;
    wire N__37655;
    wire N__37652;
    wire N__37645;
    wire N__37642;
    wire N__37641;
    wire N__37638;
    wire N__37635;
    wire N__37632;
    wire N__37627;
    wire N__37624;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37616;
    wire N__37613;
    wire N__37608;
    wire N__37607;
    wire N__37602;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37591;
    wire N__37588;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37574;
    wire N__37567;
    wire N__37566;
    wire N__37565;
    wire N__37562;
    wire N__37561;
    wire N__37558;
    wire N__37557;
    wire N__37556;
    wire N__37549;
    wire N__37546;
    wire N__37541;
    wire N__37540;
    wire N__37537;
    wire N__37536;
    wire N__37535;
    wire N__37534;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37516;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37504;
    wire N__37501;
    wire N__37500;
    wire N__37497;
    wire N__37490;
    wire N__37487;
    wire N__37484;
    wire N__37477;
    wire N__37476;
    wire N__37475;
    wire N__37474;
    wire N__37471;
    wire N__37470;
    wire N__37469;
    wire N__37468;
    wire N__37467;
    wire N__37466;
    wire N__37465;
    wire N__37460;
    wire N__37457;
    wire N__37456;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37446;
    wire N__37445;
    wire N__37444;
    wire N__37443;
    wire N__37442;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37406;
    wire N__37403;
    wire N__37402;
    wire N__37401;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37387;
    wire N__37386;
    wire N__37383;
    wire N__37380;
    wire N__37375;
    wire N__37372;
    wire N__37365;
    wire N__37360;
    wire N__37359;
    wire N__37356;
    wire N__37349;
    wire N__37346;
    wire N__37341;
    wire N__37334;
    wire N__37329;
    wire N__37326;
    wire N__37321;
    wire N__37316;
    wire N__37303;
    wire N__37300;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37288;
    wire N__37285;
    wire N__37284;
    wire N__37283;
    wire N__37278;
    wire N__37275;
    wire N__37270;
    wire N__37267;
    wire N__37266;
    wire N__37265;
    wire N__37262;
    wire N__37257;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37242;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37234;
    wire N__37231;
    wire N__37230;
    wire N__37227;
    wire N__37224;
    wire N__37221;
    wire N__37216;
    wire N__37207;
    wire N__37204;
    wire N__37203;
    wire N__37202;
    wire N__37195;
    wire N__37192;
    wire N__37191;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37171;
    wire N__37168;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37152;
    wire N__37151;
    wire N__37148;
    wire N__37143;
    wire N__37138;
    wire N__37137;
    wire N__37136;
    wire N__37135;
    wire N__37134;
    wire N__37131;
    wire N__37130;
    wire N__37129;
    wire N__37128;
    wire N__37127;
    wire N__37126;
    wire N__37125;
    wire N__37124;
    wire N__37123;
    wire N__37122;
    wire N__37117;
    wire N__37114;
    wire N__37113;
    wire N__37112;
    wire N__37111;
    wire N__37110;
    wire N__37107;
    wire N__37100;
    wire N__37099;
    wire N__37098;
    wire N__37097;
    wire N__37096;
    wire N__37095;
    wire N__37094;
    wire N__37093;
    wire N__37092;
    wire N__37091;
    wire N__37088;
    wire N__37087;
    wire N__37086;
    wire N__37085;
    wire N__37084;
    wire N__37083;
    wire N__37082;
    wire N__37079;
    wire N__37078;
    wire N__37077;
    wire N__37076;
    wire N__37075;
    wire N__37074;
    wire N__37073;
    wire N__37070;
    wire N__37069;
    wire N__37068;
    wire N__37067;
    wire N__37066;
    wire N__37065;
    wire N__37064;
    wire N__37063;
    wire N__37058;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37046;
    wire N__37045;
    wire N__37044;
    wire N__37043;
    wire N__37042;
    wire N__37039;
    wire N__37034;
    wire N__37031;
    wire N__37026;
    wire N__37023;
    wire N__37018;
    wire N__37011;
    wire N__37004;
    wire N__37003;
    wire N__37002;
    wire N__37001;
    wire N__36994;
    wire N__36989;
    wire N__36988;
    wire N__36987;
    wire N__36986;
    wire N__36985;
    wire N__36984;
    wire N__36983;
    wire N__36982;
    wire N__36981;
    wire N__36980;
    wire N__36979;
    wire N__36978;
    wire N__36973;
    wire N__36970;
    wire N__36959;
    wire N__36958;
    wire N__36957;
    wire N__36956;
    wire N__36955;
    wire N__36954;
    wire N__36953;
    wire N__36952;
    wire N__36951;
    wire N__36950;
    wire N__36949;
    wire N__36948;
    wire N__36947;
    wire N__36946;
    wire N__36945;
    wire N__36942;
    wire N__36937;
    wire N__36936;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36918;
    wire N__36909;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36897;
    wire N__36894;
    wire N__36889;
    wire N__36884;
    wire N__36881;
    wire N__36874;
    wire N__36867;
    wire N__36862;
    wire N__36853;
    wire N__36852;
    wire N__36845;
    wire N__36842;
    wire N__36841;
    wire N__36838;
    wire N__36833;
    wire N__36826;
    wire N__36819;
    wire N__36810;
    wire N__36805;
    wire N__36798;
    wire N__36797;
    wire N__36796;
    wire N__36795;
    wire N__36790;
    wire N__36785;
    wire N__36784;
    wire N__36781;
    wire N__36780;
    wire N__36777;
    wire N__36774;
    wire N__36771;
    wire N__36768;
    wire N__36759;
    wire N__36754;
    wire N__36753;
    wire N__36750;
    wire N__36749;
    wire N__36748;
    wire N__36747;
    wire N__36746;
    wire N__36733;
    wire N__36728;
    wire N__36727;
    wire N__36724;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36704;
    wire N__36699;
    wire N__36698;
    wire N__36697;
    wire N__36694;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36678;
    wire N__36673;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36627;
    wire N__36622;
    wire N__36617;
    wire N__36596;
    wire N__36591;
    wire N__36588;
    wire N__36571;
    wire N__36568;
    wire N__36565;
    wire N__36562;
    wire N__36559;
    wire N__36556;
    wire N__36555;
    wire N__36554;
    wire N__36553;
    wire N__36550;
    wire N__36549;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36541;
    wire N__36536;
    wire N__36535;
    wire N__36534;
    wire N__36533;
    wire N__36532;
    wire N__36529;
    wire N__36528;
    wire N__36525;
    wire N__36520;
    wire N__36517;
    wire N__36514;
    wire N__36513;
    wire N__36510;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36457;
    wire N__36456;
    wire N__36455;
    wire N__36454;
    wire N__36453;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36435;
    wire N__36430;
    wire N__36425;
    wire N__36422;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36375;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36342;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36325;
    wire N__36324;
    wire N__36323;
    wire N__36322;
    wire N__36321;
    wire N__36320;
    wire N__36319;
    wire N__36318;
    wire N__36317;
    wire N__36316;
    wire N__36315;
    wire N__36312;
    wire N__36311;
    wire N__36310;
    wire N__36307;
    wire N__36306;
    wire N__36305;
    wire N__36304;
    wire N__36303;
    wire N__36302;
    wire N__36301;
    wire N__36300;
    wire N__36299;
    wire N__36298;
    wire N__36297;
    wire N__36296;
    wire N__36295;
    wire N__36294;
    wire N__36293;
    wire N__36292;
    wire N__36291;
    wire N__36288;
    wire N__36287;
    wire N__36286;
    wire N__36285;
    wire N__36284;
    wire N__36283;
    wire N__36282;
    wire N__36281;
    wire N__36280;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36269;
    wire N__36262;
    wire N__36261;
    wire N__36260;
    wire N__36259;
    wire N__36258;
    wire N__36257;
    wire N__36256;
    wire N__36255;
    wire N__36254;
    wire N__36253;
    wire N__36252;
    wire N__36251;
    wire N__36250;
    wire N__36249;
    wire N__36246;
    wire N__36239;
    wire N__36236;
    wire N__36235;
    wire N__36234;
    wire N__36233;
    wire N__36232;
    wire N__36231;
    wire N__36230;
    wire N__36229;
    wire N__36228;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36220;
    wire N__36219;
    wire N__36216;
    wire N__36215;
    wire N__36214;
    wire N__36213;
    wire N__36210;
    wire N__36207;
    wire N__36206;
    wire N__36199;
    wire N__36196;
    wire N__36191;
    wire N__36186;
    wire N__36185;
    wire N__36184;
    wire N__36183;
    wire N__36180;
    wire N__36179;
    wire N__36178;
    wire N__36177;
    wire N__36174;
    wire N__36169;
    wire N__36166;
    wire N__36157;
    wire N__36156;
    wire N__36155;
    wire N__36154;
    wire N__36153;
    wire N__36152;
    wire N__36151;
    wire N__36150;
    wire N__36149;
    wire N__36148;
    wire N__36147;
    wire N__36146;
    wire N__36145;
    wire N__36144;
    wire N__36143;
    wire N__36142;
    wire N__36139;
    wire N__36138;
    wire N__36135;
    wire N__36132;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36108;
    wire N__36103;
    wire N__36102;
    wire N__36099;
    wire N__36098;
    wire N__36097;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36079;
    wire N__36074;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36052;
    wire N__36051;
    wire N__36050;
    wire N__36049;
    wire N__36048;
    wire N__36045;
    wire N__36044;
    wire N__36041;
    wire N__36036;
    wire N__36033;
    wire N__36032;
    wire N__36031;
    wire N__36030;
    wire N__36029;
    wire N__36024;
    wire N__36019;
    wire N__36018;
    wire N__36017;
    wire N__36016;
    wire N__36015;
    wire N__36014;
    wire N__36011;
    wire N__36010;
    wire N__36009;
    wire N__36002;
    wire N__35999;
    wire N__35992;
    wire N__35989;
    wire N__35986;
    wire N__35983;
    wire N__35976;
    wire N__35973;
    wire N__35972;
    wire N__35969;
    wire N__35962;
    wire N__35953;
    wire N__35952;
    wire N__35951;
    wire N__35944;
    wire N__35939;
    wire N__35936;
    wire N__35927;
    wire N__35922;
    wire N__35919;
    wire N__35918;
    wire N__35915;
    wire N__35910;
    wire N__35901;
    wire N__35896;
    wire N__35891;
    wire N__35882;
    wire N__35875;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35839;
    wire N__35836;
    wire N__35835;
    wire N__35832;
    wire N__35831;
    wire N__35830;
    wire N__35829;
    wire N__35828;
    wire N__35825;
    wire N__35822;
    wire N__35817;
    wire N__35804;
    wire N__35799;
    wire N__35792;
    wire N__35783;
    wire N__35780;
    wire N__35779;
    wire N__35778;
    wire N__35775;
    wire N__35768;
    wire N__35767;
    wire N__35766;
    wire N__35765;
    wire N__35764;
    wire N__35763;
    wire N__35758;
    wire N__35749;
    wire N__35746;
    wire N__35741;
    wire N__35734;
    wire N__35725;
    wire N__35724;
    wire N__35723;
    wire N__35722;
    wire N__35721;
    wire N__35718;
    wire N__35717;
    wire N__35716;
    wire N__35715;
    wire N__35712;
    wire N__35707;
    wire N__35704;
    wire N__35701;
    wire N__35692;
    wire N__35689;
    wire N__35676;
    wire N__35671;
    wire N__35668;
    wire N__35659;
    wire N__35656;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35632;
    wire N__35629;
    wire N__35618;
    wire N__35613;
    wire N__35612;
    wire N__35611;
    wire N__35610;
    wire N__35607;
    wire N__35598;
    wire N__35595;
    wire N__35592;
    wire N__35573;
    wire N__35552;
    wire N__35549;
    wire N__35544;
    wire N__35527;
    wire N__35524;
    wire N__35523;
    wire N__35522;
    wire N__35521;
    wire N__35520;
    wire N__35519;
    wire N__35518;
    wire N__35517;
    wire N__35516;
    wire N__35515;
    wire N__35514;
    wire N__35511;
    wire N__35510;
    wire N__35509;
    wire N__35508;
    wire N__35507;
    wire N__35506;
    wire N__35505;
    wire N__35504;
    wire N__35503;
    wire N__35502;
    wire N__35501;
    wire N__35500;
    wire N__35497;
    wire N__35496;
    wire N__35495;
    wire N__35494;
    wire N__35493;
    wire N__35492;
    wire N__35491;
    wire N__35490;
    wire N__35489;
    wire N__35488;
    wire N__35487;
    wire N__35486;
    wire N__35485;
    wire N__35484;
    wire N__35483;
    wire N__35482;
    wire N__35481;
    wire N__35480;
    wire N__35479;
    wire N__35478;
    wire N__35475;
    wire N__35474;
    wire N__35469;
    wire N__35468;
    wire N__35467;
    wire N__35466;
    wire N__35465;
    wire N__35460;
    wire N__35459;
    wire N__35458;
    wire N__35457;
    wire N__35456;
    wire N__35455;
    wire N__35452;
    wire N__35447;
    wire N__35446;
    wire N__35445;
    wire N__35444;
    wire N__35443;
    wire N__35442;
    wire N__35435;
    wire N__35432;
    wire N__35427;
    wire N__35424;
    wire N__35423;
    wire N__35420;
    wire N__35419;
    wire N__35416;
    wire N__35415;
    wire N__35412;
    wire N__35409;
    wire N__35406;
    wire N__35403;
    wire N__35398;
    wire N__35397;
    wire N__35396;
    wire N__35395;
    wire N__35394;
    wire N__35391;
    wire N__35390;
    wire N__35389;
    wire N__35388;
    wire N__35387;
    wire N__35386;
    wire N__35385;
    wire N__35384;
    wire N__35383;
    wire N__35382;
    wire N__35381;
    wire N__35380;
    wire N__35379;
    wire N__35378;
    wire N__35377;
    wire N__35376;
    wire N__35375;
    wire N__35374;
    wire N__35373;
    wire N__35372;
    wire N__35371;
    wire N__35370;
    wire N__35367;
    wire N__35358;
    wire N__35357;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35347;
    wire N__35342;
    wire N__35337;
    wire N__35332;
    wire N__35331;
    wire N__35330;
    wire N__35329;
    wire N__35326;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35305;
    wire N__35302;
    wire N__35301;
    wire N__35300;
    wire N__35297;
    wire N__35288;
    wire N__35285;
    wire N__35280;
    wire N__35279;
    wire N__35278;
    wire N__35273;
    wire N__35272;
    wire N__35269;
    wire N__35268;
    wire N__35267;
    wire N__35266;
    wire N__35265;
    wire N__35264;
    wire N__35261;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35247;
    wire N__35242;
    wire N__35239;
    wire N__35238;
    wire N__35237;
    wire N__35234;
    wire N__35229;
    wire N__35222;
    wire N__35219;
    wire N__35214;
    wire N__35207;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35199;
    wire N__35198;
    wire N__35187;
    wire N__35180;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35159;
    wire N__35152;
    wire N__35147;
    wire N__35142;
    wire N__35137;
    wire N__35128;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35110;
    wire N__35103;
    wire N__35100;
    wire N__35095;
    wire N__35090;
    wire N__35085;
    wire N__35080;
    wire N__35077;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35058;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35044;
    wire N__35039;
    wire N__35034;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__34999;
    wire N__34986;
    wire N__34979;
    wire N__34976;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34960;
    wire N__34949;
    wire N__34942;
    wire N__34935;
    wire N__34932;
    wire N__34927;
    wire N__34918;
    wire N__34917;
    wire N__34910;
    wire N__34907;
    wire N__34896;
    wire N__34893;
    wire N__34880;
    wire N__34877;
    wire N__34872;
    wire N__34869;
    wire N__34862;
    wire N__34849;
    wire N__34846;
    wire N__34845;
    wire N__34844;
    wire N__34843;
    wire N__34842;
    wire N__34841;
    wire N__34840;
    wire N__34839;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34827;
    wire N__34822;
    wire N__34821;
    wire N__34820;
    wire N__34819;
    wire N__34818;
    wire N__34817;
    wire N__34816;
    wire N__34815;
    wire N__34814;
    wire N__34813;
    wire N__34812;
    wire N__34811;
    wire N__34810;
    wire N__34809;
    wire N__34808;
    wire N__34807;
    wire N__34804;
    wire N__34803;
    wire N__34802;
    wire N__34801;
    wire N__34800;
    wire N__34799;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34795;
    wire N__34794;
    wire N__34793;
    wire N__34792;
    wire N__34791;
    wire N__34790;
    wire N__34787;
    wire N__34786;
    wire N__34785;
    wire N__34782;
    wire N__34781;
    wire N__34780;
    wire N__34779;
    wire N__34778;
    wire N__34773;
    wire N__34768;
    wire N__34765;
    wire N__34764;
    wire N__34763;
    wire N__34762;
    wire N__34761;
    wire N__34760;
    wire N__34759;
    wire N__34758;
    wire N__34755;
    wire N__34754;
    wire N__34753;
    wire N__34752;
    wire N__34751;
    wire N__34750;
    wire N__34743;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34723;
    wire N__34722;
    wire N__34717;
    wire N__34714;
    wire N__34713;
    wire N__34712;
    wire N__34711;
    wire N__34710;
    wire N__34707;
    wire N__34706;
    wire N__34705;
    wire N__34704;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34698;
    wire N__34697;
    wire N__34690;
    wire N__34683;
    wire N__34682;
    wire N__34681;
    wire N__34680;
    wire N__34677;
    wire N__34676;
    wire N__34675;
    wire N__34672;
    wire N__34665;
    wire N__34662;
    wire N__34661;
    wire N__34660;
    wire N__34657;
    wire N__34654;
    wire N__34649;
    wire N__34644;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34627;
    wire N__34624;
    wire N__34615;
    wire N__34614;
    wire N__34613;
    wire N__34612;
    wire N__34611;
    wire N__34610;
    wire N__34607;
    wire N__34606;
    wire N__34603;
    wire N__34600;
    wire N__34595;
    wire N__34590;
    wire N__34587;
    wire N__34582;
    wire N__34579;
    wire N__34574;
    wire N__34571;
    wire N__34566;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34551;
    wire N__34548;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34537;
    wire N__34536;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34528;
    wire N__34527;
    wire N__34524;
    wire N__34523;
    wire N__34518;
    wire N__34515;
    wire N__34514;
    wire N__34511;
    wire N__34506;
    wire N__34497;
    wire N__34492;
    wire N__34487;
    wire N__34484;
    wire N__34483;
    wire N__34482;
    wire N__34481;
    wire N__34476;
    wire N__34467;
    wire N__34462;
    wire N__34461;
    wire N__34460;
    wire N__34451;
    wire N__34448;
    wire N__34443;
    wire N__34436;
    wire N__34429;
    wire N__34428;
    wire N__34425;
    wire N__34420;
    wire N__34415;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34397;
    wire N__34394;
    wire N__34391;
    wire N__34384;
    wire N__34381;
    wire N__34376;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34360;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34344;
    wire N__34341;
    wire N__34334;
    wire N__34331;
    wire N__34326;
    wire N__34321;
    wire N__34318;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34300;
    wire N__34293;
    wire N__34290;
    wire N__34281;
    wire N__34276;
    wire N__34275;
    wire N__34274;
    wire N__34273;
    wire N__34272;
    wire N__34271;
    wire N__34270;
    wire N__34269;
    wire N__34268;
    wire N__34267;
    wire N__34266;
    wire N__34265;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34253;
    wire N__34246;
    wire N__34237;
    wire N__34226;
    wire N__34219;
    wire N__34212;
    wire N__34205;
    wire N__34202;
    wire N__34197;
    wire N__34190;
    wire N__34185;
    wire N__34176;
    wire N__34169;
    wire N__34156;
    wire N__34149;
    wire N__34144;
    wire N__34129;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34113;
    wire N__34112;
    wire N__34109;
    wire N__34108;
    wire N__34107;
    wire N__34106;
    wire N__34105;
    wire N__34104;
    wire N__34103;
    wire N__34102;
    wire N__34101;
    wire N__34100;
    wire N__34097;
    wire N__34096;
    wire N__34095;
    wire N__34094;
    wire N__34093;
    wire N__34092;
    wire N__34089;
    wire N__34084;
    wire N__34083;
    wire N__34082;
    wire N__34081;
    wire N__34080;
    wire N__34079;
    wire N__34078;
    wire N__34077;
    wire N__34076;
    wire N__34075;
    wire N__34072;
    wire N__34071;
    wire N__34070;
    wire N__34069;
    wire N__34064;
    wire N__34063;
    wire N__34062;
    wire N__34061;
    wire N__34060;
    wire N__34059;
    wire N__34056;
    wire N__34055;
    wire N__34054;
    wire N__34053;
    wire N__34052;
    wire N__34049;
    wire N__34048;
    wire N__34047;
    wire N__34046;
    wire N__34045;
    wire N__34042;
    wire N__34041;
    wire N__34040;
    wire N__34037;
    wire N__34036;
    wire N__34035;
    wire N__34032;
    wire N__34031;
    wire N__34030;
    wire N__34027;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34005;
    wire N__34004;
    wire N__34003;
    wire N__33996;
    wire N__33995;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33987;
    wire N__33986;
    wire N__33981;
    wire N__33980;
    wire N__33979;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33963;
    wire N__33960;
    wire N__33953;
    wire N__33952;
    wire N__33951;
    wire N__33950;
    wire N__33947;
    wire N__33946;
    wire N__33945;
    wire N__33942;
    wire N__33937;
    wire N__33936;
    wire N__33935;
    wire N__33934;
    wire N__33931;
    wire N__33926;
    wire N__33923;
    wire N__33916;
    wire N__33909;
    wire N__33906;
    wire N__33899;
    wire N__33892;
    wire N__33889;
    wire N__33884;
    wire N__33873;
    wire N__33872;
    wire N__33871;
    wire N__33868;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33837;
    wire N__33834;
    wire N__33827;
    wire N__33822;
    wire N__33813;
    wire N__33808;
    wire N__33803;
    wire N__33802;
    wire N__33799;
    wire N__33798;
    wire N__33797;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33779;
    wire N__33770;
    wire N__33765;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33746;
    wire N__33733;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33711;
    wire N__33696;
    wire N__33693;
    wire N__33682;
    wire N__33675;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33646;
    wire N__33645;
    wire N__33644;
    wire N__33643;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33635;
    wire N__33634;
    wire N__33633;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33611;
    wire N__33610;
    wire N__33609;
    wire N__33608;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33586;
    wire N__33583;
    wire N__33582;
    wire N__33581;
    wire N__33578;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33564;
    wire N__33563;
    wire N__33562;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33552;
    wire N__33547;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33525;
    wire N__33516;
    wire N__33505;
    wire N__33490;
    wire N__33489;
    wire N__33486;
    wire N__33485;
    wire N__33484;
    wire N__33483;
    wire N__33480;
    wire N__33479;
    wire N__33476;
    wire N__33475;
    wire N__33472;
    wire N__33471;
    wire N__33468;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33432;
    wire N__33431;
    wire N__33430;
    wire N__33429;
    wire N__33428;
    wire N__33421;
    wire N__33418;
    wire N__33417;
    wire N__33416;
    wire N__33415;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33383;
    wire N__33378;
    wire N__33373;
    wire N__33372;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33352;
    wire N__33347;
    wire N__33344;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33326;
    wire N__33317;
    wire N__33312;
    wire N__33301;
    wire N__33300;
    wire N__33299;
    wire N__33298;
    wire N__33297;
    wire N__33296;
    wire N__33295;
    wire N__33294;
    wire N__33293;
    wire N__33292;
    wire N__33291;
    wire N__33290;
    wire N__33289;
    wire N__33288;
    wire N__33287;
    wire N__33284;
    wire N__33283;
    wire N__33282;
    wire N__33281;
    wire N__33280;
    wire N__33279;
    wire N__33276;
    wire N__33275;
    wire N__33274;
    wire N__33273;
    wire N__33272;
    wire N__33271;
    wire N__33270;
    wire N__33269;
    wire N__33268;
    wire N__33267;
    wire N__33266;
    wire N__33265;
    wire N__33264;
    wire N__33263;
    wire N__33260;
    wire N__33259;
    wire N__33258;
    wire N__33257;
    wire N__33254;
    wire N__33253;
    wire N__33252;
    wire N__33251;
    wire N__33250;
    wire N__33249;
    wire N__33248;
    wire N__33245;
    wire N__33244;
    wire N__33241;
    wire N__33240;
    wire N__33237;
    wire N__33236;
    wire N__33235;
    wire N__33234;
    wire N__33233;
    wire N__33232;
    wire N__33229;
    wire N__33224;
    wire N__33223;
    wire N__33220;
    wire N__33219;
    wire N__33218;
    wire N__33217;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33199;
    wire N__33198;
    wire N__33197;
    wire N__33196;
    wire N__33193;
    wire N__33192;
    wire N__33191;
    wire N__33190;
    wire N__33187;
    wire N__33186;
    wire N__33185;
    wire N__33184;
    wire N__33183;
    wire N__33176;
    wire N__33169;
    wire N__33168;
    wire N__33167;
    wire N__33166;
    wire N__33165;
    wire N__33164;
    wire N__33163;
    wire N__33162;
    wire N__33161;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33143;
    wire N__33138;
    wire N__33137;
    wire N__33136;
    wire N__33135;
    wire N__33130;
    wire N__33125;
    wire N__33124;
    wire N__33117;
    wire N__33110;
    wire N__33103;
    wire N__33102;
    wire N__33101;
    wire N__33100;
    wire N__33099;
    wire N__33098;
    wire N__33097;
    wire N__33094;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33084;
    wire N__33079;
    wire N__33074;
    wire N__33069;
    wire N__33066;
    wire N__33065;
    wire N__33064;
    wire N__33061;
    wire N__33056;
    wire N__33053;
    wire N__33044;
    wire N__33041;
    wire N__33032;
    wire N__33031;
    wire N__33026;
    wire N__33023;
    wire N__33022;
    wire N__33015;
    wire N__33012;
    wire N__33007;
    wire N__33000;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32978;
    wire N__32973;
    wire N__32968;
    wire N__32967;
    wire N__32966;
    wire N__32965;
    wire N__32962;
    wire N__32961;
    wire N__32960;
    wire N__32959;
    wire N__32958;
    wire N__32957;
    wire N__32956;
    wire N__32955;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32907;
    wire N__32904;
    wire N__32899;
    wire N__32892;
    wire N__32887;
    wire N__32878;
    wire N__32877;
    wire N__32874;
    wire N__32869;
    wire N__32866;
    wire N__32857;
    wire N__32854;
    wire N__32853;
    wire N__32852;
    wire N__32851;
    wire N__32848;
    wire N__32845;
    wire N__32842;
    wire N__32833;
    wire N__32828;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32816;
    wire N__32811;
    wire N__32804;
    wire N__32799;
    wire N__32790;
    wire N__32789;
    wire N__32788;
    wire N__32787;
    wire N__32786;
    wire N__32785;
    wire N__32782;
    wire N__32781;
    wire N__32780;
    wire N__32779;
    wire N__32778;
    wire N__32775;
    wire N__32766;
    wire N__32761;
    wire N__32750;
    wire N__32747;
    wire N__32736;
    wire N__32731;
    wire N__32728;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32701;
    wire N__32696;
    wire N__32695;
    wire N__32694;
    wire N__32691;
    wire N__32686;
    wire N__32683;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32667;
    wire N__32658;
    wire N__32651;
    wire N__32644;
    wire N__32635;
    wire N__32630;
    wire N__32605;
    wire N__32602;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32594;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32586;
    wire N__32585;
    wire N__32582;
    wire N__32581;
    wire N__32578;
    wire N__32573;
    wire N__32570;
    wire N__32565;
    wire N__32560;
    wire N__32551;
    wire N__32550;
    wire N__32549;
    wire N__32548;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32472;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32466;
    wire N__32461;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32449;
    wire N__32446;
    wire N__32443;
    wire N__32438;
    wire N__32435;
    wire N__32434;
    wire N__32433;
    wire N__32426;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32407;
    wire N__32404;
    wire N__32401;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32386;
    wire N__32383;
    wire N__32380;
    wire N__32379;
    wire N__32378;
    wire N__32377;
    wire N__32374;
    wire N__32373;
    wire N__32372;
    wire N__32369;
    wire N__32368;
    wire N__32363;
    wire N__32360;
    wire N__32357;
    wire N__32356;
    wire N__32355;
    wire N__32354;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32331;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32308;
    wire N__32305;
    wire N__32302;
    wire N__32295;
    wire N__32290;
    wire N__32281;
    wire N__32278;
    wire N__32275;
    wire N__32274;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32251;
    wire N__32248;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32236;
    wire N__32233;
    wire N__32232;
    wire N__32231;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32210;
    wire N__32207;
    wire N__32204;
    wire N__32201;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32190;
    wire N__32189;
    wire N__32188;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32170;
    wire N__32169;
    wire N__32164;
    wire N__32161;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32134;
    wire N__32133;
    wire N__32132;
    wire N__32131;
    wire N__32128;
    wire N__32127;
    wire N__32126;
    wire N__32125;
    wire N__32124;
    wire N__32123;
    wire N__32122;
    wire N__32121;
    wire N__32120;
    wire N__32119;
    wire N__32118;
    wire N__32117;
    wire N__32116;
    wire N__32115;
    wire N__32114;
    wire N__32113;
    wire N__32112;
    wire N__32111;
    wire N__32110;
    wire N__32109;
    wire N__32108;
    wire N__32107;
    wire N__32106;
    wire N__32101;
    wire N__32100;
    wire N__32099;
    wire N__32098;
    wire N__32097;
    wire N__32096;
    wire N__32095;
    wire N__32094;
    wire N__32093;
    wire N__32092;
    wire N__32091;
    wire N__32088;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32080;
    wire N__32079;
    wire N__32078;
    wire N__32077;
    wire N__32076;
    wire N__32075;
    wire N__32072;
    wire N__32071;
    wire N__32066;
    wire N__32065;
    wire N__32064;
    wire N__32063;
    wire N__32060;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32046;
    wire N__32045;
    wire N__32044;
    wire N__32043;
    wire N__32042;
    wire N__32041;
    wire N__32038;
    wire N__32035;
    wire N__32034;
    wire N__32033;
    wire N__32030;
    wire N__32025;
    wire N__32024;
    wire N__32023;
    wire N__32022;
    wire N__32021;
    wire N__32020;
    wire N__32019;
    wire N__32018;
    wire N__32015;
    wire N__32012;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31996;
    wire N__31989;
    wire N__31982;
    wire N__31981;
    wire N__31980;
    wire N__31979;
    wire N__31978;
    wire N__31975;
    wire N__31974;
    wire N__31973;
    wire N__31968;
    wire N__31961;
    wire N__31960;
    wire N__31959;
    wire N__31958;
    wire N__31957;
    wire N__31956;
    wire N__31955;
    wire N__31950;
    wire N__31945;
    wire N__31944;
    wire N__31943;
    wire N__31942;
    wire N__31941;
    wire N__31940;
    wire N__31939;
    wire N__31938;
    wire N__31937;
    wire N__31936;
    wire N__31935;
    wire N__31934;
    wire N__31933;
    wire N__31932;
    wire N__31931;
    wire N__31928;
    wire N__31923;
    wire N__31922;
    wire N__31921;
    wire N__31920;
    wire N__31919;
    wire N__31918;
    wire N__31917;
    wire N__31916;
    wire N__31915;
    wire N__31914;
    wire N__31913;
    wire N__31912;
    wire N__31909;
    wire N__31908;
    wire N__31907;
    wire N__31906;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31898;
    wire N__31897;
    wire N__31896;
    wire N__31893;
    wire N__31886;
    wire N__31885;
    wire N__31884;
    wire N__31881;
    wire N__31880;
    wire N__31879;
    wire N__31878;
    wire N__31877;
    wire N__31876;
    wire N__31875;
    wire N__31872;
    wire N__31865;
    wire N__31858;
    wire N__31855;
    wire N__31844;
    wire N__31839;
    wire N__31834;
    wire N__31829;
    wire N__31828;
    wire N__31827;
    wire N__31826;
    wire N__31823;
    wire N__31818;
    wire N__31815;
    wire N__31810;
    wire N__31801;
    wire N__31798;
    wire N__31789;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31769;
    wire N__31766;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31746;
    wire N__31745;
    wire N__31744;
    wire N__31743;
    wire N__31738;
    wire N__31735;
    wire N__31730;
    wire N__31725;
    wire N__31720;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31704;
    wire N__31699;
    wire N__31694;
    wire N__31691;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31672;
    wire N__31671;
    wire N__31666;
    wire N__31661;
    wire N__31658;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31642;
    wire N__31639;
    wire N__31634;
    wire N__31625;
    wire N__31618;
    wire N__31611;
    wire N__31606;
    wire N__31601;
    wire N__31598;
    wire N__31593;
    wire N__31582;
    wire N__31573;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31555;
    wire N__31550;
    wire N__31549;
    wire N__31548;
    wire N__31547;
    wire N__31546;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31538;
    wire N__31535;
    wire N__31528;
    wire N__31525;
    wire N__31520;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31499;
    wire N__31494;
    wire N__31487;
    wire N__31476;
    wire N__31471;
    wire N__31470;
    wire N__31469;
    wire N__31468;
    wire N__31463;
    wire N__31458;
    wire N__31455;
    wire N__31448;
    wire N__31445;
    wire N__31436;
    wire N__31431;
    wire N__31428;
    wire N__31423;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31409;
    wire N__31398;
    wire N__31389;
    wire N__31384;
    wire N__31377;
    wire N__31372;
    wire N__31365;
    wire N__31362;
    wire N__31333;
    wire N__31332;
    wire N__31331;
    wire N__31330;
    wire N__31329;
    wire N__31328;
    wire N__31327;
    wire N__31326;
    wire N__31325;
    wire N__31324;
    wire N__31323;
    wire N__31322;
    wire N__31321;
    wire N__31320;
    wire N__31319;
    wire N__31318;
    wire N__31317;
    wire N__31316;
    wire N__31315;
    wire N__31314;
    wire N__31313;
    wire N__31312;
    wire N__31311;
    wire N__31310;
    wire N__31309;
    wire N__31308;
    wire N__31307;
    wire N__31306;
    wire N__31305;
    wire N__31304;
    wire N__31303;
    wire N__31302;
    wire N__31301;
    wire N__31300;
    wire N__31299;
    wire N__31298;
    wire N__31297;
    wire N__31296;
    wire N__31291;
    wire N__31286;
    wire N__31285;
    wire N__31276;
    wire N__31271;
    wire N__31262;
    wire N__31253;
    wire N__31252;
    wire N__31251;
    wire N__31250;
    wire N__31249;
    wire N__31244;
    wire N__31241;
    wire N__31240;
    wire N__31239;
    wire N__31238;
    wire N__31237;
    wire N__31236;
    wire N__31235;
    wire N__31232;
    wire N__31231;
    wire N__31230;
    wire N__31229;
    wire N__31228;
    wire N__31227;
    wire N__31226;
    wire N__31225;
    wire N__31224;
    wire N__31223;
    wire N__31222;
    wire N__31221;
    wire N__31220;
    wire N__31217;
    wire N__31216;
    wire N__31215;
    wire N__31214;
    wire N__31213;
    wire N__31212;
    wire N__31211;
    wire N__31210;
    wire N__31209;
    wire N__31208;
    wire N__31207;
    wire N__31206;
    wire N__31203;
    wire N__31196;
    wire N__31189;
    wire N__31188;
    wire N__31187;
    wire N__31182;
    wire N__31175;
    wire N__31174;
    wire N__31173;
    wire N__31168;
    wire N__31167;
    wire N__31166;
    wire N__31165;
    wire N__31164;
    wire N__31163;
    wire N__31162;
    wire N__31161;
    wire N__31160;
    wire N__31159;
    wire N__31156;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31138;
    wire N__31131;
    wire N__31130;
    wire N__31127;
    wire N__31122;
    wire N__31113;
    wire N__31112;
    wire N__31111;
    wire N__31110;
    wire N__31105;
    wire N__31102;
    wire N__31097;
    wire N__31096;
    wire N__31095;
    wire N__31094;
    wire N__31093;
    wire N__31092;
    wire N__31091;
    wire N__31090;
    wire N__31089;
    wire N__31088;
    wire N__31087;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31073;
    wire N__31072;
    wire N__31071;
    wire N__31070;
    wire N__31069;
    wire N__31068;
    wire N__31065;
    wire N__31058;
    wire N__31051;
    wire N__31050;
    wire N__31049;
    wire N__31048;
    wire N__31045;
    wire N__31042;
    wire N__31041;
    wire N__31036;
    wire N__31031;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31008;
    wire N__31003;
    wire N__30998;
    wire N__30995;
    wire N__30986;
    wire N__30975;
    wire N__30974;
    wire N__30973;
    wire N__30972;
    wire N__30971;
    wire N__30970;
    wire N__30967;
    wire N__30956;
    wire N__30955;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30943;
    wire N__30940;
    wire N__30939;
    wire N__30938;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30926;
    wire N__30923;
    wire N__30916;
    wire N__30913;
    wire N__30908;
    wire N__30907;
    wire N__30906;
    wire N__30901;
    wire N__30898;
    wire N__30893;
    wire N__30886;
    wire N__30881;
    wire N__30874;
    wire N__30867;
    wire N__30860;
    wire N__30859;
    wire N__30858;
    wire N__30857;
    wire N__30854;
    wire N__30851;
    wire N__30848;
    wire N__30843;
    wire N__30832;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30808;
    wire N__30803;
    wire N__30798;
    wire N__30789;
    wire N__30788;
    wire N__30787;
    wire N__30786;
    wire N__30785;
    wire N__30778;
    wire N__30775;
    wire N__30764;
    wire N__30761;
    wire N__30756;
    wire N__30747;
    wire N__30738;
    wire N__30733;
    wire N__30730;
    wire N__30729;
    wire N__30728;
    wire N__30727;
    wire N__30722;
    wire N__30721;
    wire N__30720;
    wire N__30719;
    wire N__30718;
    wire N__30717;
    wire N__30716;
    wire N__30715;
    wire N__30714;
    wire N__30711;
    wire N__30704;
    wire N__30701;
    wire N__30694;
    wire N__30689;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30668;
    wire N__30659;
    wire N__30656;
    wire N__30649;
    wire N__30646;
    wire N__30641;
    wire N__30636;
    wire N__30629;
    wire N__30626;
    wire N__30621;
    wire N__30614;
    wire N__30607;
    wire N__30598;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30534;
    wire N__30533;
    wire N__30532;
    wire N__30531;
    wire N__30528;
    wire N__30527;
    wire N__30526;
    wire N__30525;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30515;
    wire N__30512;
    wire N__30511;
    wire N__30510;
    wire N__30509;
    wire N__30508;
    wire N__30507;
    wire N__30504;
    wire N__30503;
    wire N__30500;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30488;
    wire N__30487;
    wire N__30482;
    wire N__30479;
    wire N__30478;
    wire N__30475;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30414;
    wire N__30411;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30395;
    wire N__30394;
    wire N__30393;
    wire N__30392;
    wire N__30391;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30369;
    wire N__30360;
    wire N__30357;
    wire N__30346;
    wire N__30345;
    wire N__30344;
    wire N__30343;
    wire N__30342;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30329;
    wire N__30328;
    wire N__30327;
    wire N__30326;
    wire N__30325;
    wire N__30324;
    wire N__30323;
    wire N__30322;
    wire N__30321;
    wire N__30320;
    wire N__30319;
    wire N__30318;
    wire N__30315;
    wire N__30314;
    wire N__30313;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30293;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30277;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30260;
    wire N__30259;
    wire N__30258;
    wire N__30255;
    wire N__30250;
    wire N__30247;
    wire N__30240;
    wire N__30237;
    wire N__30232;
    wire N__30227;
    wire N__30222;
    wire N__30219;
    wire N__30214;
    wire N__30211;
    wire N__30206;
    wire N__30203;
    wire N__30194;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30147;
    wire N__30146;
    wire N__30145;
    wire N__30144;
    wire N__30143;
    wire N__30142;
    wire N__30135;
    wire N__30134;
    wire N__30131;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30113;
    wire N__30110;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30084;
    wire N__30083;
    wire N__30080;
    wire N__30075;
    wire N__30074;
    wire N__30073;
    wire N__30072;
    wire N__30067;
    wire N__30066;
    wire N__30065;
    wire N__30064;
    wire N__30063;
    wire N__30062;
    wire N__30059;
    wire N__30058;
    wire N__30055;
    wire N__30054;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30043;
    wire N__30042;
    wire N__30039;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30028;
    wire N__30027;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30010;
    wire N__30005;
    wire N__30000;
    wire N__29997;
    wire N__29994;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29932;
    wire N__29931;
    wire N__29926;
    wire N__29917;
    wire N__29912;
    wire N__29907;
    wire N__29904;
    wire N__29899;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29883;
    wire N__29878;
    wire N__29875;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29871;
    wire N__29870;
    wire N__29865;
    wire N__29856;
    wire N__29851;
    wire N__29848;
    wire N__29847;
    wire N__29842;
    wire N__29839;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29827;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29814;
    wire N__29813;
    wire N__29812;
    wire N__29811;
    wire N__29806;
    wire N__29803;
    wire N__29802;
    wire N__29799;
    wire N__29798;
    wire N__29795;
    wire N__29794;
    wire N__29789;
    wire N__29784;
    wire N__29777;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29760;
    wire N__29759;
    wire N__29758;
    wire N__29757;
    wire N__29754;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29734;
    wire N__29725;
    wire N__29724;
    wire N__29723;
    wire N__29720;
    wire N__29719;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29711;
    wire N__29710;
    wire N__29707;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29661;
    wire N__29658;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29634;
    wire N__29629;
    wire N__29628;
    wire N__29627;
    wire N__29626;
    wire N__29623;
    wire N__29622;
    wire N__29621;
    wire N__29620;
    wire N__29619;
    wire N__29618;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29600;
    wire N__29597;
    wire N__29596;
    wire N__29595;
    wire N__29592;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29577;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29549;
    wire N__29548;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29529;
    wire N__29526;
    wire N__29521;
    wire N__29516;
    wire N__29509;
    wire N__29504;
    wire N__29501;
    wire N__29496;
    wire N__29491;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29448;
    wire N__29447;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29412;
    wire N__29409;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29401;
    wire N__29400;
    wire N__29397;
    wire N__29396;
    wire N__29395;
    wire N__29392;
    wire N__29389;
    wire N__29384;
    wire N__29381;
    wire N__29376;
    wire N__29373;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29355;
    wire N__29354;
    wire N__29347;
    wire N__29346;
    wire N__29345;
    wire N__29344;
    wire N__29341;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29298;
    wire N__29297;
    wire N__29290;
    wire N__29287;
    wire N__29286;
    wire N__29285;
    wire N__29282;
    wire N__29277;
    wire N__29272;
    wire N__29271;
    wire N__29270;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29262;
    wire N__29261;
    wire N__29260;
    wire N__29259;
    wire N__29256;
    wire N__29255;
    wire N__29254;
    wire N__29251;
    wire N__29246;
    wire N__29243;
    wire N__29242;
    wire N__29241;
    wire N__29238;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29220;
    wire N__29217;
    wire N__29216;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29184;
    wire N__29181;
    wire N__29180;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29169;
    wire N__29168;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29152;
    wire N__29149;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29117;
    wire N__29116;
    wire N__29113;
    wire N__29108;
    wire N__29105;
    wire N__29100;
    wire N__29097;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29067;
    wire N__29062;
    wire N__29057;
    wire N__29054;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29029;
    wire N__29024;
    wire N__29019;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28980;
    wire N__28979;
    wire N__28978;
    wire N__28977;
    wire N__28974;
    wire N__28973;
    wire N__28972;
    wire N__28971;
    wire N__28966;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28939;
    wire N__28936;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28921;
    wire N__28920;
    wire N__28919;
    wire N__28918;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28910;
    wire N__28909;
    wire N__28906;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28889;
    wire N__28886;
    wire N__28883;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28873;
    wire N__28866;
    wire N__28863;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28839;
    wire N__28836;
    wire N__28835;
    wire N__28834;
    wire N__28833;
    wire N__28832;
    wire N__28831;
    wire N__28830;
    wire N__28827;
    wire N__28822;
    wire N__28817;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28795;
    wire N__28780;
    wire N__28777;
    wire N__28776;
    wire N__28773;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28753;
    wire N__28752;
    wire N__28751;
    wire N__28750;
    wire N__28749;
    wire N__28748;
    wire N__28747;
    wire N__28746;
    wire N__28745;
    wire N__28744;
    wire N__28743;
    wire N__28742;
    wire N__28741;
    wire N__28740;
    wire N__28739;
    wire N__28738;
    wire N__28737;
    wire N__28736;
    wire N__28735;
    wire N__28734;
    wire N__28733;
    wire N__28720;
    wire N__28707;
    wire N__28694;
    wire N__28693;
    wire N__28692;
    wire N__28691;
    wire N__28690;
    wire N__28689;
    wire N__28686;
    wire N__28681;
    wire N__28680;
    wire N__28679;
    wire N__28678;
    wire N__28677;
    wire N__28676;
    wire N__28675;
    wire N__28674;
    wire N__28671;
    wire N__28666;
    wire N__28665;
    wire N__28664;
    wire N__28663;
    wire N__28662;
    wire N__28661;
    wire N__28660;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28630;
    wire N__28629;
    wire N__28628;
    wire N__28627;
    wire N__28626;
    wire N__28625;
    wire N__28624;
    wire N__28623;
    wire N__28622;
    wire N__28621;
    wire N__28620;
    wire N__28619;
    wire N__28618;
    wire N__28617;
    wire N__28616;
    wire N__28615;
    wire N__28614;
    wire N__28613;
    wire N__28612;
    wire N__28611;
    wire N__28610;
    wire N__28609;
    wire N__28608;
    wire N__28607;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28584;
    wire N__28581;
    wire N__28574;
    wire N__28559;
    wire N__28546;
    wire N__28533;
    wire N__28522;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28483;
    wire N__28480;
    wire N__28479;
    wire N__28478;
    wire N__28477;
    wire N__28476;
    wire N__28475;
    wire N__28474;
    wire N__28473;
    wire N__28472;
    wire N__28469;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28451;
    wire N__28450;
    wire N__28449;
    wire N__28448;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28438;
    wire N__28435;
    wire N__28426;
    wire N__28425;
    wire N__28424;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28381;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28352;
    wire N__28349;
    wire N__28344;
    wire N__28339;
    wire N__28338;
    wire N__28335;
    wire N__28334;
    wire N__28331;
    wire N__28330;
    wire N__28329;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28302;
    wire N__28299;
    wire N__28298;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28266;
    wire N__28263;
    wire N__28258;
    wire N__28253;
    wire N__28250;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28207;
    wire N__28204;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28189;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28174;
    wire N__28173;
    wire N__28172;
    wire N__28169;
    wire N__28164;
    wire N__28159;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28144;
    wire N__28143;
    wire N__28138;
    wire N__28135;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28123;
    wire N__28122;
    wire N__28119;
    wire N__28118;
    wire N__28117;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28103;
    wire N__28102;
    wire N__28099;
    wire N__28098;
    wire N__28095;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28071;
    wire N__28066;
    wire N__28061;
    wire N__28054;
    wire N__28053;
    wire N__28052;
    wire N__28051;
    wire N__28050;
    wire N__28049;
    wire N__28048;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28015;
    wire N__28010;
    wire N__28005;
    wire N__28004;
    wire N__28001;
    wire N__27996;
    wire N__27991;
    wire N__27988;
    wire N__27979;
    wire N__27978;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27970;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27946;
    wire N__27943;
    wire N__27942;
    wire N__27941;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27933;
    wire N__27930;
    wire N__27929;
    wire N__27926;
    wire N__27925;
    wire N__27924;
    wire N__27923;
    wire N__27918;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27859;
    wire N__27858;
    wire N__27855;
    wire N__27854;
    wire N__27853;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27835;
    wire N__27834;
    wire N__27829;
    wire N__27826;
    wire N__27825;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27813;
    wire N__27808;
    wire N__27805;
    wire N__27804;
    wire N__27799;
    wire N__27796;
    wire N__27795;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27760;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27738;
    wire N__27737;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27725;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27711;
    wire N__27708;
    wire N__27707;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27695;
    wire N__27692;
    wire N__27685;
    wire N__27684;
    wire N__27681;
    wire N__27680;
    wire N__27673;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27658;
    wire N__27657;
    wire N__27652;
    wire N__27649;
    wire N__27648;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27636;
    wire N__27631;
    wire N__27628;
    wire N__27627;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27609;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27561;
    wire N__27560;
    wire N__27559;
    wire N__27558;
    wire N__27555;
    wire N__27554;
    wire N__27553;
    wire N__27552;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27537;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27525;
    wire N__27524;
    wire N__27523;
    wire N__27520;
    wire N__27515;
    wire N__27514;
    wire N__27511;
    wire N__27510;
    wire N__27509;
    wire N__27506;
    wire N__27501;
    wire N__27498;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27482;
    wire N__27477;
    wire N__27472;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27461;
    wire N__27458;
    wire N__27457;
    wire N__27452;
    wire N__27449;
    wire N__27442;
    wire N__27435;
    wire N__27432;
    wire N__27425;
    wire N__27418;
    wire N__27409;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27393;
    wire N__27392;
    wire N__27391;
    wire N__27390;
    wire N__27389;
    wire N__27388;
    wire N__27387;
    wire N__27386;
    wire N__27383;
    wire N__27382;
    wire N__27379;
    wire N__27378;
    wire N__27375;
    wire N__27374;
    wire N__27371;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27363;
    wire N__27362;
    wire N__27359;
    wire N__27358;
    wire N__27357;
    wire N__27354;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27346;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27325;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27277;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27262;
    wire N__27255;
    wire N__27250;
    wire N__27245;
    wire N__27242;
    wire N__27233;
    wire N__27226;
    wire N__27223;
    wire N__27218;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27171;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27163;
    wire N__27160;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27133;
    wire N__27130;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27099;
    wire N__27096;
    wire N__27091;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27039;
    wire N__27038;
    wire N__27037;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27023;
    wire N__27022;
    wire N__27019;
    wire N__27018;
    wire N__27013;
    wire N__27012;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26962;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26937;
    wire N__26934;
    wire N__26933;
    wire N__26932;
    wire N__26931;
    wire N__26928;
    wire N__26927;
    wire N__26926;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26912;
    wire N__26907;
    wire N__26906;
    wire N__26899;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26883;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26802;
    wire N__26799;
    wire N__26798;
    wire N__26797;
    wire N__26794;
    wire N__26793;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26781;
    wire N__26780;
    wire N__26779;
    wire N__26776;
    wire N__26775;
    wire N__26774;
    wire N__26773;
    wire N__26772;
    wire N__26769;
    wire N__26768;
    wire N__26767;
    wire N__26762;
    wire N__26759;
    wire N__26758;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26739;
    wire N__26738;
    wire N__26737;
    wire N__26736;
    wire N__26733;
    wire N__26728;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26698;
    wire N__26689;
    wire N__26680;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26616;
    wire N__26615;
    wire N__26612;
    wire N__26611;
    wire N__26610;
    wire N__26609;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26587;
    wire N__26586;
    wire N__26585;
    wire N__26584;
    wire N__26583;
    wire N__26578;
    wire N__26575;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26556;
    wire N__26553;
    wire N__26548;
    wire N__26543;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26504;
    wire N__26501;
    wire N__26500;
    wire N__26497;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26484;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26458;
    wire N__26453;
    wire N__26446;
    wire N__26445;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26384;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26360;
    wire N__26355;
    wire N__26350;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26317;
    wire N__26316;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26293;
    wire N__26288;
    wire N__26287;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26259;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26226;
    wire N__26223;
    wire N__26222;
    wire N__26221;
    wire N__26218;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26183;
    wire N__26182;
    wire N__26181;
    wire N__26176;
    wire N__26173;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26152;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26131;
    wire N__26130;
    wire N__26129;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26106;
    wire N__26103;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26047;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25992;
    wire N__25989;
    wire N__25988;
    wire N__25985;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25937;
    wire N__25936;
    wire N__25933;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25903;
    wire N__25894;
    wire N__25893;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25845;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25809;
    wire N__25808;
    wire N__25807;
    wire N__25806;
    wire N__25805;
    wire N__25804;
    wire N__25801;
    wire N__25798;
    wire N__25797;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25768;
    wire N__25763;
    wire N__25756;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25738;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25650;
    wire N__25649;
    wire N__25646;
    wire N__25645;
    wire N__25644;
    wire N__25643;
    wire N__25642;
    wire N__25641;
    wire N__25640;
    wire N__25639;
    wire N__25636;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25563;
    wire N__25560;
    wire N__25555;
    wire N__25552;
    wire N__25547;
    wire N__25544;
    wire N__25537;
    wire N__25532;
    wire N__25527;
    wire N__25522;
    wire N__25519;
    wire N__25518;
    wire N__25517;
    wire N__25516;
    wire N__25515;
    wire N__25512;
    wire N__25507;
    wire N__25504;
    wire N__25501;
    wire N__25500;
    wire N__25499;
    wire N__25494;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25482;
    wire N__25481;
    wire N__25480;
    wire N__25479;
    wire N__25478;
    wire N__25477;
    wire N__25468;
    wire N__25467;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25455;
    wire N__25450;
    wire N__25449;
    wire N__25446;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25395;
    wire N__25392;
    wire N__25381;
    wire N__25378;
    wire N__25377;
    wire N__25376;
    wire N__25375;
    wire N__25374;
    wire N__25369;
    wire N__25368;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25360;
    wire N__25359;
    wire N__25358;
    wire N__25355;
    wire N__25354;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25343;
    wire N__25340;
    wire N__25339;
    wire N__25338;
    wire N__25333;
    wire N__25330;
    wire N__25329;
    wire N__25326;
    wire N__25325;
    wire N__25320;
    wire N__25317;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25298;
    wire N__25295;
    wire N__25290;
    wire N__25285;
    wire N__25282;
    wire N__25275;
    wire N__25270;
    wire N__25255;
    wire N__25254;
    wire N__25249;
    wire N__25248;
    wire N__25247;
    wire N__25244;
    wire N__25239;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25221;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25195;
    wire N__25194;
    wire N__25189;
    wire N__25186;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25110;
    wire N__25107;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25083;
    wire N__25080;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25068;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25050;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25000;
    wire N__24997;
    wire N__24996;
    wire N__24995;
    wire N__24992;
    wire N__24987;
    wire N__24986;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24963;
    wire N__24960;
    wire N__24959;
    wire N__24956;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24934;
    wire N__24933;
    wire N__24930;
    wire N__24929;
    wire N__24928;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24910;
    wire N__24909;
    wire N__24904;
    wire N__24901;
    wire N__24900;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24888;
    wire N__24883;
    wire N__24880;
    wire N__24879;
    wire N__24874;
    wire N__24871;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24856;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24844;
    wire N__24841;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24817;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24805;
    wire N__24802;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24784;
    wire N__24781;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24751;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24733;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24721;
    wire N__24718;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24706;
    wire N__24705;
    wire N__24700;
    wire N__24697;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24682;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24652;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24640;
    wire N__24637;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24622;
    wire N__24619;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24555;
    wire N__24554;
    wire N__24553;
    wire N__24552;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24541;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24502;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24462;
    wire N__24461;
    wire N__24460;
    wire N__24459;
    wire N__24458;
    wire N__24455;
    wire N__24454;
    wire N__24453;
    wire N__24452;
    wire N__24449;
    wire N__24448;
    wire N__24445;
    wire N__24442;
    wire N__24441;
    wire N__24438;
    wire N__24437;
    wire N__24434;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24426;
    wire N__24425;
    wire N__24422;
    wire N__24413;
    wire N__24410;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24391;
    wire N__24384;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24333;
    wire N__24330;
    wire N__24329;
    wire N__24328;
    wire N__24325;
    wire N__24324;
    wire N__24323;
    wire N__24322;
    wire N__24319;
    wire N__24318;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24290;
    wire N__24289;
    wire N__24288;
    wire N__24287;
    wire N__24284;
    wire N__24279;
    wire N__24274;
    wire N__24269;
    wire N__24266;
    wire N__24259;
    wire N__24256;
    wire N__24249;
    wire N__24246;
    wire N__24237;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24219;
    wire N__24218;
    wire N__24215;
    wire N__24210;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24198;
    wire N__24197;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24186;
    wire N__24185;
    wire N__24184;
    wire N__24181;
    wire N__24180;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24169;
    wire N__24166;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24144;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24094;
    wire N__24091;
    wire N__24086;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24031;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__24000;
    wire N__23999;
    wire N__23996;
    wire N__23995;
    wire N__23994;
    wire N__23993;
    wire N__23992;
    wire N__23989;
    wire N__23988;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23968;
    wire N__23967;
    wire N__23966;
    wire N__23965;
    wire N__23962;
    wire N__23957;
    wire N__23954;
    wire N__23953;
    wire N__23952;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23929;
    wire N__23926;
    wire N__23921;
    wire N__23916;
    wire N__23913;
    wire N__23906;
    wire N__23903;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23856;
    wire N__23853;
    wire N__23852;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23844;
    wire N__23843;
    wire N__23840;
    wire N__23839;
    wire N__23836;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23800;
    wire N__23797;
    wire N__23790;
    wire N__23785;
    wire N__23782;
    wire N__23777;
    wire N__23774;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23742;
    wire N__23741;
    wire N__23738;
    wire N__23733;
    wire N__23732;
    wire N__23731;
    wire N__23730;
    wire N__23729;
    wire N__23728;
    wire N__23727;
    wire N__23726;
    wire N__23721;
    wire N__23720;
    wire N__23719;
    wire N__23716;
    wire N__23711;
    wire N__23706;
    wire N__23701;
    wire N__23698;
    wire N__23693;
    wire N__23690;
    wire N__23677;
    wire N__23676;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23616;
    wire N__23613;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23586;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23553;
    wire N__23550;
    wire N__23549;
    wire N__23548;
    wire N__23547;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23496;
    wire N__23495;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23263;
    wire N__23260;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23217;
    wire N__23216;
    wire N__23215;
    wire N__23212;
    wire N__23211;
    wire N__23210;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23178;
    wire N__23173;
    wire N__23170;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23150;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22971;
    wire N__22966;
    wire N__22963;
    wire N__22962;
    wire N__22957;
    wire N__22954;
    wire N__22953;
    wire N__22948;
    wire N__22945;
    wire N__22944;
    wire N__22943;
    wire N__22940;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22932;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22915;
    wire N__22914;
    wire N__22911;
    wire N__22906;
    wire N__22903;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22885;
    wire N__22876;
    wire N__22875;
    wire N__22874;
    wire N__22871;
    wire N__22870;
    wire N__22869;
    wire N__22868;
    wire N__22865;
    wire N__22864;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22832;
    wire N__22827;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22807;
    wire N__22806;
    wire N__22803;
    wire N__22802;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22791;
    wire N__22790;
    wire N__22787;
    wire N__22780;
    wire N__22779;
    wire N__22776;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22702;
    wire N__22699;
    wire N__22698;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22686;
    wire N__22681;
    wire N__22678;
    wire N__22677;
    wire N__22672;
    wire N__22669;
    wire N__22668;
    wire N__22663;
    wire N__22660;
    wire N__22659;
    wire N__22656;
    wire N__22655;
    wire N__22650;
    wire N__22647;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22610;
    wire N__22607;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22585;
    wire N__22584;
    wire N__22583;
    wire N__22582;
    wire N__22579;
    wire N__22572;
    wire N__22567;
    wire N__22566;
    wire N__22561;
    wire N__22558;
    wire N__22557;
    wire N__22552;
    wire N__22549;
    wire N__22548;
    wire N__22543;
    wire N__22540;
    wire N__22539;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22527;
    wire N__22522;
    wire N__22519;
    wire N__22518;
    wire N__22513;
    wire N__22510;
    wire N__22509;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22497;
    wire N__22496;
    wire N__22491;
    wire N__22488;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22468;
    wire N__22465;
    wire N__22464;
    wire N__22461;
    wire N__22460;
    wire N__22457;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22435;
    wire N__22434;
    wire N__22433;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22421;
    wire N__22418;
    wire N__22411;
    wire N__22410;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22334;
    wire N__22333;
    wire N__22328;
    wire N__22323;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22308;
    wire N__22307;
    wire N__22306;
    wire N__22303;
    wire N__22298;
    wire N__22295;
    wire N__22288;
    wire N__22287;
    wire N__22286;
    wire N__22279;
    wire N__22278;
    wire N__22275;
    wire N__22272;
    wire N__22269;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22251;
    wire N__22250;
    wire N__22249;
    wire N__22246;
    wire N__22245;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22233;
    wire N__22232;
    wire N__22229;
    wire N__22228;
    wire N__22225;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22195;
    wire N__22192;
    wire N__22191;
    wire N__22190;
    wire N__22189;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22168;
    wire N__22167;
    wire N__22162;
    wire N__22159;
    wire N__22154;
    wire N__22149;
    wire N__22144;
    wire N__22139;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22123;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22029;
    wire N__22028;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22014;
    wire N__22011;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21992;
    wire N__21991;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21955;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21841;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21774;
    wire N__21773;
    wire N__21772;
    wire N__21769;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21646;
    wire N__21643;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21486;
    wire N__21481;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21381;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21352;
    wire N__21349;
    wire N__21348;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21244;
    wire N__21243;
    wire N__21240;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21219;
    wire N__21214;
    wire N__21211;
    wire N__21210;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21171;
    wire N__21168;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21146;
    wire N__21143;
    wire N__21138;
    wire N__21133;
    wire N__21130;
    wire N__21129;
    wire N__21128;
    wire N__21125;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21103;
    wire N__21102;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21090;
    wire N__21089;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21073;
    wire N__21070;
    wire N__21069;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21057;
    wire N__21056;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21044;
    wire N__21037;
    wire N__21034;
    wire N__21033;
    wire N__21030;
    wire N__21029;
    wire N__21028;
    wire N__21025;
    wire N__21020;
    wire N__21017;
    wire N__21010;
    wire N__21009;
    wire N__21008;
    wire N__21005;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20993;
    wire N__20986;
    wire N__20985;
    wire N__20980;
    wire N__20977;
    wire N__20976;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20964;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20793;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20785;
    wire N__20782;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20770;
    wire N__20769;
    wire N__20768;
    wire N__20767;
    wire N__20766;
    wire N__20765;
    wire N__20762;
    wire N__20761;
    wire N__20760;
    wire N__20759;
    wire N__20758;
    wire N__20751;
    wire N__20748;
    wire N__20741;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20724;
    wire N__20721;
    wire N__20716;
    wire N__20713;
    wire N__20698;
    wire N__20695;
    wire N__20692;
    wire N__20691;
    wire N__20690;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20670;
    wire N__20665;
    wire N__20660;
    wire N__20657;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20574;
    wire N__20573;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20559;
    wire N__20558;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20541;
    wire N__20538;
    wire N__20535;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20426;
    wire N__20425;
    wire N__20422;
    wire N__20417;
    wire N__20416;
    wire N__20413;
    wire N__20412;
    wire N__20407;
    wire N__20406;
    wire N__20405;
    wire N__20404;
    wire N__20401;
    wire N__20400;
    wire N__20397;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20377;
    wire N__20374;
    wire N__20369;
    wire N__20366;
    wire N__20361;
    wire N__20356;
    wire N__20347;
    wire N__20344;
    wire N__20343;
    wire N__20342;
    wire N__20341;
    wire N__20340;
    wire N__20339;
    wire N__20336;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20322;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20291;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20259;
    wire N__20258;
    wire N__20253;
    wire N__20250;
    wire N__20249;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20238;
    wire N__20235;
    wire N__20230;
    wire N__20227;
    wire N__20226;
    wire N__20223;
    wire N__20216;
    wire N__20213;
    wire N__20208;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20180;
    wire N__20179;
    wire N__20178;
    wire N__20177;
    wire N__20174;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20094;
    wire N__20091;
    wire N__20090;
    wire N__20089;
    wire N__20088;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20077;
    wire N__20076;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20042;
    wire N__20037;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19906;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19881;
    wire N__19878;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19752;
    wire N__19751;
    wire N__19750;
    wire N__19749;
    wire N__19748;
    wire N__19739;
    wire N__19738;
    wire N__19737;
    wire N__19732;
    wire N__19731;
    wire N__19730;
    wire N__19729;
    wire N__19728;
    wire N__19725;
    wire N__19720;
    wire N__19719;
    wire N__19718;
    wire N__19717;
    wire N__19716;
    wire N__19713;
    wire N__19708;
    wire N__19703;
    wire N__19698;
    wire N__19689;
    wire N__19686;
    wire N__19681;
    wire N__19676;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19504;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19487;
    wire N__19482;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19470;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19389;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19335;
    wire N__19334;
    wire N__19333;
    wire N__19330;
    wire N__19325;
    wire N__19322;
    wire N__19321;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19304;
    wire N__19301;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19278;
    wire N__19275;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19251;
    wire N__19248;
    wire N__19247;
    wire N__19246;
    wire N__19245;
    wire N__19244;
    wire N__19241;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19218;
    wire N__19215;
    wire N__19214;
    wire N__19209;
    wire N__19206;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19180;
    wire N__19177;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18972;
    wire N__18969;
    wire N__18964;
    wire N__18963;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18955;
    wire N__18952;
    wire N__18951;
    wire N__18950;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18928;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18912;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18834;
    wire N__18833;
    wire N__18832;
    wire N__18829;
    wire N__18828;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18813;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18776;
    wire N__18773;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18753;
    wire N__18750;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18729;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18705;
    wire N__18702;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18688;
    wire N__18687;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18592;
    wire N__18589;
    wire N__18588;
    wire N__18587;
    wire N__18586;
    wire N__18585;
    wire N__18584;
    wire N__18583;
    wire N__18582;
    wire N__18581;
    wire N__18578;
    wire N__18573;
    wire N__18570;
    wire N__18569;
    wire N__18566;
    wire N__18565;
    wire N__18564;
    wire N__18563;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18551;
    wire N__18550;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18519;
    wire N__18516;
    wire N__18511;
    wire N__18506;
    wire N__18503;
    wire N__18496;
    wire N__18491;
    wire N__18486;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18457;
    wire N__18456;
    wire N__18455;
    wire N__18454;
    wire N__18453;
    wire N__18452;
    wire N__18451;
    wire N__18450;
    wire N__18449;
    wire N__18448;
    wire N__18447;
    wire N__18446;
    wire N__18445;
    wire N__18444;
    wire N__18443;
    wire N__18442;
    wire N__18441;
    wire N__18440;
    wire N__18439;
    wire N__18424;
    wire N__18409;
    wire N__18398;
    wire N__18397;
    wire N__18396;
    wire N__18395;
    wire N__18394;
    wire N__18393;
    wire N__18392;
    wire N__18391;
    wire N__18390;
    wire N__18389;
    wire N__18388;
    wire N__18387;
    wire N__18386;
    wire N__18385;
    wire N__18384;
    wire N__18383;
    wire N__18382;
    wire N__18381;
    wire N__18380;
    wire N__18379;
    wire N__18378;
    wire N__18377;
    wire N__18376;
    wire N__18375;
    wire N__18374;
    wire N__18373;
    wire N__18372;
    wire N__18371;
    wire N__18370;
    wire N__18369;
    wire N__18368;
    wire N__18367;
    wire N__18366;
    wire N__18365;
    wire N__18364;
    wire N__18363;
    wire N__18362;
    wire N__18361;
    wire N__18360;
    wire N__18359;
    wire N__18358;
    wire N__18357;
    wire N__18356;
    wire N__18355;
    wire N__18354;
    wire N__18353;
    wire N__18352;
    wire N__18351;
    wire N__18350;
    wire N__18349;
    wire N__18348;
    wire N__18347;
    wire N__18346;
    wire N__18345;
    wire N__18338;
    wire N__18323;
    wire N__18322;
    wire N__18321;
    wire N__18320;
    wire N__18319;
    wire N__18318;
    wire N__18317;
    wire N__18316;
    wire N__18299;
    wire N__18282;
    wire N__18277;
    wire N__18260;
    wire N__18255;
    wire N__18254;
    wire N__18253;
    wire N__18238;
    wire N__18223;
    wire N__18220;
    wire N__18219;
    wire N__18218;
    wire N__18217;
    wire N__18216;
    wire N__18209;
    wire N__18204;
    wire N__18203;
    wire N__18202;
    wire N__18201;
    wire N__18200;
    wire N__18199;
    wire N__18198;
    wire N__18197;
    wire N__18196;
    wire N__18195;
    wire N__18194;
    wire N__18193;
    wire N__18192;
    wire N__18191;
    wire N__18190;
    wire N__18189;
    wire N__18188;
    wire N__18187;
    wire N__18186;
    wire N__18185;
    wire N__18184;
    wire N__18183;
    wire N__18182;
    wire N__18181;
    wire N__18180;
    wire N__18179;
    wire N__18178;
    wire N__18177;
    wire N__18176;
    wire N__18175;
    wire N__18174;
    wire N__18173;
    wire N__18172;
    wire N__18171;
    wire N__18170;
    wire N__18169;
    wire N__18168;
    wire N__18167;
    wire N__18152;
    wire N__18145;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18127;
    wire N__18118;
    wire N__18117;
    wire N__18116;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18108;
    wire N__18101;
    wire N__18088;
    wire N__18073;
    wire N__18058;
    wire N__18045;
    wire N__18028;
    wire N__18021;
    wire N__18016;
    wire N__18011;
    wire N__18008;
    wire N__17999;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17956;
    wire N__17955;
    wire N__17952;
    wire N__17949;
    wire N__17948;
    wire N__17947;
    wire N__17946;
    wire N__17943;
    wire N__17940;
    wire N__17937;
    wire N__17936;
    wire N__17935;
    wire N__17934;
    wire N__17933;
    wire N__17932;
    wire N__17931;
    wire N__17928;
    wire N__17927;
    wire N__17926;
    wire N__17925;
    wire N__17924;
    wire N__17923;
    wire N__17920;
    wire N__17919;
    wire N__17916;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17904;
    wire N__17903;
    wire N__17902;
    wire N__17901;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17887;
    wire N__17886;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17875;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17828;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17814;
    wire N__17813;
    wire N__17812;
    wire N__17811;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17795;
    wire N__17792;
    wire N__17787;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17767;
    wire N__17758;
    wire N__17757;
    wire N__17754;
    wire N__17753;
    wire N__17750;
    wire N__17749;
    wire N__17746;
    wire N__17741;
    wire N__17734;
    wire N__17729;
    wire N__17722;
    wire N__17719;
    wire N__17710;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17535;
    wire N__17532;
    wire N__17529;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17518;
    wire N__17517;
    wire N__17516;
    wire N__17515;
    wire N__17510;
    wire N__17509;
    wire N__17508;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17497;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17448;
    wire N__17445;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17425;
    wire N__17422;
    wire N__17421;
    wire N__17418;
    wire N__17415;
    wire N__17414;
    wire N__17409;
    wire N__17406;
    wire N__17403;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17319;
    wire N__17318;
    wire N__17315;
    wire N__17314;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17299;
    wire N__17298;
    wire N__17289;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17266;
    wire N__17265;
    wire N__17262;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17251;
    wire N__17250;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17235;
    wire N__17232;
    wire N__17229;
    wire N__17224;
    wire N__17221;
    wire N__17220;
    wire N__17217;
    wire N__17214;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17198;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17013;
    wire N__17012;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17000;
    wire N__16997;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16981;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16909;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16884;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16858;
    wire N__16855;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16825;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16794;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16782;
    wire N__16781;
    wire N__16780;
    wire N__16779;
    wire N__16776;
    wire N__16775;
    wire N__16772;
    wire N__16771;
    wire N__16770;
    wire N__16769;
    wire N__16766;
    wire N__16761;
    wire N__16758;
    wire N__16755;
    wire N__16748;
    wire N__16745;
    wire N__16740;
    wire N__16729;
    wire N__16728;
    wire N__16727;
    wire N__16720;
    wire N__16717;
    wire N__16716;
    wire N__16715;
    wire N__16714;
    wire N__16711;
    wire N__16704;
    wire N__16699;
    wire N__16696;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16678;
    wire N__16677;
    wire N__16672;
    wire N__16671;
    wire N__16670;
    wire N__16669;
    wire N__16668;
    wire N__16667;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16657;
    wire N__16648;
    wire N__16643;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16599;
    wire N__16594;
    wire N__16591;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16579;
    wire N__16576;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16552;
    wire N__16549;
    wire N__16546;
    wire N__16543;
    wire N__16540;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16528;
    wire N__16527;
    wire N__16524;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16405;
    wire N__16404;
    wire N__16399;
    wire N__16396;
    wire N__16393;
    wire N__16390;
    wire N__16389;
    wire N__16386;
    wire N__16383;
    wire N__16378;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16366;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16354;
    wire N__16351;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16260;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16243;
    wire N__16240;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16228;
    wire N__16227;
    wire N__16222;
    wire N__16219;
    wire N__16218;
    wire N__16213;
    wire N__16210;
    wire N__16209;
    wire N__16204;
    wire N__16201;
    wire N__16200;
    wire N__16195;
    wire N__16192;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16119;
    wire N__16118;
    wire N__16117;
    wire N__16116;
    wire N__16115;
    wire N__16114;
    wire N__16113;
    wire N__16108;
    wire N__16101;
    wire N__16094;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16021;
    wire N__16018;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15963;
    wire N__15958;
    wire N__15955;
    wire N__15954;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15933;
    wire N__15928;
    wire N__15925;
    wire N__15924;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15845;
    wire N__15844;
    wire N__15841;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15817;
    wire N__15814;
    wire N__15809;
    wire N__15802;
    wire N__15801;
    wire N__15798;
    wire N__15797;
    wire N__15796;
    wire N__15789;
    wire N__15788;
    wire N__15787;
    wire N__15784;
    wire N__15783;
    wire N__15780;
    wire N__15773;
    wire N__15772;
    wire N__15771;
    wire N__15768;
    wire N__15767;
    wire N__15766;
    wire N__15763;
    wire N__15760;
    wire N__15749;
    wire N__15742;
    wire N__15741;
    wire N__15740;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15726;
    wire N__15725;
    wire N__15724;
    wire N__15723;
    wire N__15714;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15686;
    wire N__15681;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15632;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15608;
    wire N__15603;
    wire N__15602;
    wire N__15599;
    wire N__15596;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15542;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15517;
    wire N__15514;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15502;
    wire N__15499;
    wire N__15494;
    wire N__15491;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15461;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15441;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15419;
    wire N__15412;
    wire N__15411;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15398;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15379;
    wire N__15378;
    wire N__15373;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15352;
    wire N__15351;
    wire N__15346;
    wire N__15343;
    wire N__15340;
    wire N__15339;
    wire N__15334;
    wire N__15331;
    wire N__15328;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15286;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15274;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15259;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15247;
    wire N__15246;
    wire N__15241;
    wire N__15238;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15226;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15214;
    wire N__15213;
    wire N__15210;
    wire N__15207;
    wire N__15202;
    wire N__15201;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15184;
    wire N__15181;
    wire N__15180;
    wire N__15175;
    wire N__15172;
    wire N__15171;
    wire N__15166;
    wire N__15163;
    wire N__15162;
    wire N__15157;
    wire N__15154;
    wire N__15153;
    wire N__15148;
    wire N__15145;
    wire N__15144;
    wire N__15139;
    wire N__15136;
    wire N__15135;
    wire N__15130;
    wire N__15127;
    wire N__15126;
    wire N__15121;
    wire N__15118;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15106;
    wire N__15105;
    wire N__15100;
    wire N__15097;
    wire N__15096;
    wire N__15091;
    wire N__15088;
    wire N__15087;
    wire N__15082;
    wire N__15079;
    wire N__15078;
    wire N__15073;
    wire N__15070;
    wire N__15069;
    wire N__15064;
    wire N__15061;
    wire N__15060;
    wire N__15055;
    wire N__15052;
    wire N__15049;
    wire N__15048;
    wire N__15043;
    wire N__15040;
    wire N__15039;
    wire N__15034;
    wire N__15031;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15016;
    wire N__15015;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__15001;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14964;
    wire N__14961;
    wire N__14958;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14835;
    wire N__14830;
    wire N__14827;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14799;
    wire N__14794;
    wire N__14791;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14779;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14752;
    wire N__14751;
    wire N__14748;
    wire N__14745;
    wire N__14740;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14725;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14684;
    wire N__14683;
    wire N__14682;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14520;
    wire N__14517;
    wire N__14516;
    wire N__14515;
    wire N__14514;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14478;
    wire N__14475;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14463;
    wire N__14460;
    wire N__14457;
    wire N__14454;
    wire N__14453;
    wire N__14452;
    wire N__14451;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14425;
    wire N__14424;
    wire N__14419;
    wire N__14416;
    wire N__14415;
    wire N__14410;
    wire N__14407;
    wire N__14406;
    wire N__14401;
    wire N__14398;
    wire N__14397;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14376;
    wire N__14373;
    wire N__14370;
    wire N__14365;
    wire N__14364;
    wire N__14361;
    wire N__14358;
    wire N__14355;
    wire N__14350;
    wire N__14347;
    wire N__14346;
    wire N__14343;
    wire N__14340;
    wire N__14335;
    wire N__14332;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14313;
    wire N__14310;
    wire N__14307;
    wire N__14302;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14290;
    wire N__14289;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14277;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14265;
    wire N__14260;
    wire N__14257;
    wire N__14256;
    wire N__14251;
    wire N__14248;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14236;
    wire N__14235;
    wire N__14232;
    wire N__14229;
    wire N__14224;
    wire N__14223;
    wire N__14220;
    wire N__14217;
    wire N__14212;
    wire N__14211;
    wire N__14206;
    wire N__14203;
    wire N__14202;
    wire N__14197;
    wire N__14194;
    wire N__14193;
    wire N__14188;
    wire N__14185;
    wire N__14184;
    wire N__14179;
    wire N__14176;
    wire N__14175;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14157;
    wire N__14154;
    wire N__14151;
    wire N__14146;
    wire N__14145;
    wire N__14142;
    wire N__14139;
    wire N__14134;
    wire N__14131;
    wire N__14130;
    wire N__14127;
    wire N__14124;
    wire N__14119;
    wire N__14116;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14104;
    wire N__14101;
    wire N__14100;
    wire N__14097;
    wire N__14094;
    wire N__14089;
    wire N__14086;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14074;
    wire N__14071;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14059;
    wire N__14056;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14013;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13992;
    wire N__13989;
    wire N__13986;
    wire N__13983;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13956;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13878;
    wire N__13875;
    wire N__13872;
    wire N__13869;
    wire N__13864;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13852;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13840;
    wire N__13839;
    wire N__13834;
    wire N__13831;
    wire N__13830;
    wire N__13825;
    wire N__13822;
    wire N__13821;
    wire N__13816;
    wire N__13813;
    wire N__13812;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13800;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13777;
    wire N__13776;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13729;
    wire N__13726;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13695;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13681;
    wire N__13678;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13666;
    wire N__13665;
    wire N__13662;
    wire N__13659;
    wire N__13654;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13642;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13630;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13609;
    wire N__13608;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13594;
    wire N__13593;
    wire N__13588;
    wire N__13585;
    wire N__13584;
    wire N__13579;
    wire N__13576;
    wire N__13573;
    wire N__13572;
    wire N__13567;
    wire N__13564;
    wire N__13563;
    wire N__13560;
    wire N__13557;
    wire N__13554;
    wire N__13549;
    wire N__13548;
    wire N__13543;
    wire N__13540;
    wire N__13539;
    wire N__13536;
    wire N__13533;
    wire N__13528;
    wire N__13527;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13515;
    wire N__13510;
    wire N__13507;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13495;
    wire N__13494;
    wire N__13491;
    wire N__13488;
    wire N__13483;
    wire N__13480;
    wire N__13477;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13465;
    wire N__13464;
    wire N__13461;
    wire N__13458;
    wire N__13455;
    wire N__13452;
    wire N__13447;
    wire N__13444;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13432;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13420;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13402;
    wire N__13401;
    wire N__13398;
    wire N__13395;
    wire N__13392;
    wire N__13389;
    wire N__13384;
    wire N__13381;
    wire N__13378;
    wire N__13375;
    wire N__13372;
    wire N__13369;
    wire N__13368;
    wire N__13365;
    wire N__13362;
    wire N__13359;
    wire N__13354;
    wire N__13353;
    wire N__13350;
    wire N__13347;
    wire N__13342;
    wire N__13341;
    wire N__13336;
    wire N__13333;
    wire N__13332;
    wire N__13327;
    wire N__13324;
    wire N__13323;
    wire N__13318;
    wire N__13315;
    wire N__13314;
    wire N__13309;
    wire N__13306;
    wire N__13305;
    wire N__13300;
    wire N__13297;
    wire N__13296;
    wire N__13291;
    wire N__13288;
    wire N__13287;
    wire N__13282;
    wire N__13279;
    wire N__13276;
    wire N__13273;
    wire N__13272;
    wire N__13269;
    wire N__13266;
    wire N__13261;
    wire N__13260;
    wire N__13257;
    wire N__13254;
    wire N__13251;
    wire N__13248;
    wire N__13245;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13219;
    wire N__13218;
    wire N__13213;
    wire N__13210;
    wire N__13209;
    wire N__13204;
    wire N__13201;
    wire N__13200;
    wire N__13195;
    wire N__13192;
    wire N__13191;
    wire N__13186;
    wire N__13183;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13171;
    wire N__13168;
    wire N__13167;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13155;
    wire N__13152;
    wire N__13149;
    wire N__13144;
    wire N__13143;
    wire N__13138;
    wire N__13135;
    wire N__13132;
    wire N__13131;
    wire N__13126;
    wire N__13123;
    wire N__13122;
    wire N__13117;
    wire N__13114;
    wire N__13113;
    wire N__13108;
    wire N__13105;
    wire N__13104;
    wire N__13099;
    wire N__13096;
    wire N__13095;
    wire N__13090;
    wire N__13087;
    wire N__13086;
    wire N__13081;
    wire N__13078;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13066;
    wire N__13065;
    wire N__13060;
    wire N__13057;
    wire N__13056;
    wire N__13051;
    wire N__13048;
    wire N__13047;
    wire N__13042;
    wire VCCG0;
    wire \tok.A_stk.tail_73 ;
    wire \tok.A_stk.tail_93 ;
    wire \tok.A_stk.tail_77 ;
    wire \tok.A_stk.tail_61 ;
    wire \tok.A_stk.tail_45 ;
    wire \tok.A_stk.tail_29 ;
    wire \tok.A_stk.tail_13 ;
    wire \tok.A_stk.tail_75 ;
    wire \tok.A_stk.tail_59 ;
    wire \tok.A_stk.tail_43 ;
    wire \tok.A_stk.tail_27 ;
    wire \tok.A_stk.tail_85 ;
    wire \tok.A_stk.tail_69 ;
    wire \tok.A_stk.tail_53 ;
    wire \tok.A_stk.tail_37 ;
    wire \tok.A_stk.tail_21 ;
    wire \tok.A_stk.tail_5 ;
    wire \tok.A_stk.tail_11 ;
    wire \tok.A_stk.tail_9 ;
    wire \tok.A_stk.tail_25 ;
    wire \tok.A_stk.tail_57 ;
    wire \tok.A_stk.tail_41 ;
    wire \tok.table_rd_10 ;
    wire \tok.n203_adj_866_cascade_ ;
    wire \tok.n212_adj_867_cascade_ ;
    wire \tok.n6426_cascade_ ;
    wire tail_80;
    wire \tok.A_stk.tail_64 ;
    wire tail_48;
    wire \tok.A_stk.tail_32 ;
    wire tail_16;
    wire tail_96;
    wire tail_112;
    wire tail_118;
    wire \tok.table_wr_data_8 ;
    wire \tok.A_stk.tail_89 ;
    wire tail_122;
    wire tail_106;
    wire \tok.A_stk.tail_90 ;
    wire \tok.A_stk.tail_74 ;
    wire \tok.A_stk.tail_58 ;
    wire \tok.A_stk.tail_42 ;
    wire tail_109;
    wire tail_125;
    wire \tok.n6274 ;
    wire \tok.n34_cascade_ ;
    wire A_stk_delta_1_cascade_;
    wire tail_105;
    wire tail_121;
    wire tail_101;
    wire tail_117;
    wire \tok.n34 ;
    wire tail_100;
    wire rd_15__N_300_cascade_;
    wire tail_116;
    wire \tok.A_stk.tail_91 ;
    wire tail_123;
    wire tail_107;
    wire \tok.A_stk.tail_84 ;
    wire \tok.A_stk.tail_68 ;
    wire \tok.A_stk.tail_52 ;
    wire \tok.A_stk.tail_36 ;
    wire \tok.A_stk.tail_20 ;
    wire \tok.A_stk.tail_0 ;
    wire \tok.A_stk.tail_4 ;
    wire bfn_1_7_0_;
    wire \tok.n4767 ;
    wire \tok.n4768 ;
    wire \tok.n4769 ;
    wire \tok.n4770 ;
    wire \tok.n4771 ;
    wire \tok.n4772 ;
    wire \tok.n4773 ;
    wire tail_120;
    wire tail_104;
    wire \tok.A_stk.tail_88 ;
    wire \tok.A_stk.tail_72 ;
    wire \tok.A_stk.tail_56 ;
    wire \tok.A_stk.tail_40 ;
    wire \tok.A_stk.tail_24 ;
    wire \tok.A_stk.tail_8 ;
    wire \tok.table_rd_13 ;
    wire \tok.n226_cascade_ ;
    wire \tok.n203_adj_643_cascade_ ;
    wire \tok.n226 ;
    wire \tok.n212_adj_646_cascade_ ;
    wire \tok.n6448_cascade_ ;
    wire \tok.n6388 ;
    wire \tok.n206_adj_649 ;
    wire \tok.table_rd_9 ;
    wire \tok.n203_adj_833_cascade_ ;
    wire \tok.n212_adj_835_cascade_ ;
    wire \tok.n206_adj_834 ;
    wire \tok.n6443_cascade_ ;
    wire \tok.n242_adj_839_cascade_ ;
    wire \tok.n230 ;
    wire \tok.n242_adj_874 ;
    wire \tok.n6431_cascade_ ;
    wire \tok.n206_adj_869 ;
    wire \tok.n206_adj_691 ;
    wire \tok.n212_adj_689_cascade_ ;
    wire \tok.n229_adj_863 ;
    wire \tok.uart.n6223_cascade_ ;
    wire txtick_cascade_;
    wire \tok.uart.n12 ;
    wire \tok.uart.txclkcounter_0 ;
    wire bfn_1_13_0_;
    wire \tok.uart.txclkcounter_1 ;
    wire \tok.uart.n4830 ;
    wire \tok.uart.txclkcounter_2 ;
    wire \tok.uart.n4831 ;
    wire \tok.uart.txclkcounter_3 ;
    wire \tok.uart.n4832 ;
    wire \tok.uart.txclkcounter_4 ;
    wire \tok.uart.n4833 ;
    wire \tok.uart.txclkcounter_5 ;
    wire \tok.uart.n4834 ;
    wire \tok.uart.txclkcounter_6 ;
    wire \tok.uart.n4835 ;
    wire \tok.uart.txclkcounter_7 ;
    wire \tok.uart.n4836 ;
    wire \tok.uart.n4837 ;
    wire bfn_1_14_0_;
    wire \tok.uart.txclkcounter_8 ;
    wire tail_127;
    wire tail_111;
    wire \tok.A_stk.tail_95 ;
    wire \tok.A_stk.tail_79 ;
    wire \tok.A_stk.tail_63 ;
    wire \tok.A_stk.tail_47 ;
    wire \tok.A_stk.tail_31 ;
    wire \tok.A_stk.tail_15 ;
    wire \tok.A_stk.tail_26 ;
    wire tail_126;
    wire tail_110;
    wire \tok.A_stk.tail_94 ;
    wire \tok.A_stk.tail_78 ;
    wire \tok.A_stk.tail_62 ;
    wire \tok.A_stk.tail_46 ;
    wire \tok.A_stk.tail_30 ;
    wire \tok.A_stk.tail_14 ;
    wire \tok.A_stk.tail_34 ;
    wire \tok.A_stk.tail_50 ;
    wire \tok.A_stk.tail_66 ;
    wire \tok.A_stk.tail_82 ;
    wire table_wr_data_0;
    wire tail_98;
    wire tail_114;
    wire \tok.n4_adj_642_cascade_ ;
    wire \tok.table_wr_data_13 ;
    wire \tok.table_wr_data_10 ;
    wire \tok.table_wr_data_15 ;
    wire \tok.n33_adj_631 ;
    wire \tok.n27_cascade_ ;
    wire \tok.n41 ;
    wire \tok.n33_adj_662 ;
    wire \tok.n27_adj_709_cascade_ ;
    wire \tok.n19 ;
    wire \tok.n33_adj_634 ;
    wire \tok.n27_adj_706_cascade_ ;
    wire \tok.n35 ;
    wire \tok.n6667_cascade_ ;
    wire \tok.n2532 ;
    wire \tok.n4_adj_642 ;
    wire \tok.found_slot_cascade_ ;
    wire \tok.write_slot ;
    wire \tok.n21_cascade_ ;
    wire \tok.n30_adj_647 ;
    wire \tok.key_rd_10 ;
    wire \tok.key_rd_12 ;
    wire \tok.n26 ;
    wire \tok.n27_adj_639_cascade_ ;
    wire \tok.found_slot_N_144 ;
    wire \tok.n6322 ;
    wire \tok.n313_cascade_ ;
    wire \tok.key_rd_2 ;
    wire \tok.key_rd_7 ;
    wire \tok.n22 ;
    wire \tok.table_rd_12 ;
    wire \tok.n227 ;
    wire \tok.n203_cascade_ ;
    wire \tok.n212_cascade_ ;
    wire \tok.n206 ;
    wire bfn_2_10_0_;
    wire \tok.n4774 ;
    wire \tok.n4775 ;
    wire \tok.n4776 ;
    wire \tok.n4777 ;
    wire \tok.n4778 ;
    wire \tok.n4779 ;
    wire \tok.n4780 ;
    wire \tok.n4781 ;
    wire bfn_2_11_0_;
    wire \tok.n214_cascade_ ;
    wire \tok.n6358 ;
    wire \tok.n6402 ;
    wire \tok.table_rd_14 ;
    wire \tok.n225_cascade_ ;
    wire \tok.n203_adj_664_cascade_ ;
    wire \tok.n225 ;
    wire \tok.n224 ;
    wire \tok.table_rd_15 ;
    wire \tok.n224_cascade_ ;
    wire \tok.n203_adj_688 ;
    wire \tok.n6373_cascade_ ;
    wire \tok.n206_adj_666_cascade_ ;
    wire \tok.n212_adj_665 ;
    wire \tok.n281_cascade_ ;
    wire \tok.n236_adj_864_cascade_ ;
    wire \tok.n2648_cascade_ ;
    wire \tok.n226_adj_865 ;
    wire \tok.n6334 ;
    wire \tok.n4_adj_762 ;
    wire \tok.n6316 ;
    wire sender_1;
    wire tx_c;
    wire \tok.A_stk.tail_65 ;
    wire tail_49;
    wire tail_81;
    wire \tok.A_stk.tail_33 ;
    wire tail_17;
    wire \tok.A_stk.tail_1 ;
    wire tail_102;
    wire \tok.A_stk.tail_86 ;
    wire \tok.A_stk.tail_70 ;
    wire \tok.A_stk.tail_54 ;
    wire \tok.A_stk.tail_38 ;
    wire \tok.A_stk.tail_22 ;
    wire \tok.A_stk.tail_28 ;
    wire \tok.A_stk.tail_44 ;
    wire \tok.A_stk.tail_92 ;
    wire \tok.A_stk.tail_60 ;
    wire \tok.A_stk.tail_76 ;
    wire \tok.A_stk.tail_6 ;
    wire \tok.A_stk.tail_12 ;
    wire \tok.A_stk.tail_10 ;
    wire \tok.A_stk.tail_83 ;
    wire \tok.A_stk.tail_67 ;
    wire \tok.A_stk.tail_51 ;
    wire \tok.A_stk.tail_35 ;
    wire \tok.A_stk.tail_19 ;
    wire \tok.A_stk.tail_3 ;
    wire \tok.n4_cascade_ ;
    wire \tok.n6273 ;
    wire \tok.table_wr_data_9 ;
    wire \tok.n4 ;
    wire \tok.n6252 ;
    wire \tok.n6253_cascade_ ;
    wire tail_99;
    wire tail_115;
    wire \tok.n33_adj_633 ;
    wire \tok.n27_adj_704_cascade_ ;
    wire \tok.n38 ;
    wire \tok.n33_adj_632 ;
    wire \tok.n33_adj_661 ;
    wire \tok.n27_adj_705_cascade_ ;
    wire \tok.n36 ;
    wire \tok.n27_adj_703 ;
    wire \tok.n40 ;
    wire \tok.n32 ;
    wire \tok.n33 ;
    wire \tok.n27_adj_707 ;
    wire \tok.n33_adj_663 ;
    wire \tok.n27_adj_708_cascade_ ;
    wire \tok.n29 ;
    wire \tok.search_clk ;
    wire \tok.found_slot ;
    wire \tok.n6670 ;
    wire \tok.key_rd_6 ;
    wire \tok.key_rd_0 ;
    wire \tok.n25 ;
    wire \tok.key_rd_4 ;
    wire \tok.key_rd_1 ;
    wire \tok.n18 ;
    wire \tok.n6575_cascade_ ;
    wire \tok.n177 ;
    wire bfn_4_9_0_;
    wire \tok.n4797 ;
    wire \tok.n4798 ;
    wire \tok.n4799 ;
    wire \tok.n6556 ;
    wire \tok.n4800 ;
    wire \tok.n4801 ;
    wire \tok.n4802 ;
    wire \tok.n4803 ;
    wire \tok.n4803_THRU_CRY_0_THRU_CO ;
    wire bfn_4_10_0_;
    wire \tok.n4804 ;
    wire \tok.n6437 ;
    wire \tok.n4805 ;
    wire \tok.n4806 ;
    wire \tok.n4807 ;
    wire \tok.n4808 ;
    wire \tok.n6377 ;
    wire \tok.n4809 ;
    wire \tok.n4810 ;
    wire \tok.n4810_THRU_CRY_0_THRU_CO ;
    wire bfn_4_11_0_;
    wire \tok.n4811 ;
    wire \tok.n6362 ;
    wire \tok.n83 ;
    wire \tok.n161_adj_836 ;
    wire \tok.n197_adj_837_cascade_ ;
    wire \tok.n248_adj_838 ;
    wire \tok.n161_adj_650 ;
    wire \tok.n6386_cascade_ ;
    wire \tok.n197_adj_652_cascade_ ;
    wire \tok.table_rd_11 ;
    wire \tok.n228_cascade_ ;
    wire \tok.n203_adj_879_cascade_ ;
    wire \tok.n228 ;
    wire \tok.n212_adj_880_cascade_ ;
    wire \tok.n6339 ;
    wire \tok.n161_adj_692_cascade_ ;
    wire \tok.n6356 ;
    wire \tok.n6417 ;
    wire \tok.n206_adj_881 ;
    wire \tok.n6412 ;
    wire tail_119;
    wire tail_103;
    wire \tok.A_stk.tail_87 ;
    wire \tok.A_stk.tail_71 ;
    wire \tok.A_stk.tail_55 ;
    wire \tok.A_stk.tail_39 ;
    wire \tok.A_stk.tail_23 ;
    wire \tok.A_stk.tail_7 ;
    wire tail_97;
    wire tail_113;
    wire tail_108;
    wire tail_124;
    wire \tok.table_wr_data_3 ;
    wire table_wr_data_1;
    wire \tok.table_wr_data_6 ;
    wire \tok.table_wr_data_4 ;
    wire \tok.table_wr_data_2 ;
    wire \tok.ram.n6266_cascade_ ;
    wire \tok.n1495_cascade_ ;
    wire \tok.n13_adj_766 ;
    wire n10_adj_907;
    wire n10_adj_907_cascade_;
    wire \tok.tc_6 ;
    wire \tok.n83_adj_765_cascade_ ;
    wire \tok.n6435 ;
    wire \tok.n6283_cascade_ ;
    wire \tok.n80_cascade_ ;
    wire \tok.n89_cascade_ ;
    wire \tok.n83_adj_734_cascade_ ;
    wire \tok.n6279 ;
    wire \tok.table_rd_0 ;
    wire \tok.table_wr_data_14 ;
    wire \tok.table_wr_data_11 ;
    wire \tok.table_wr_data_12 ;
    wire \tok.n2696 ;
    wire \tok.n9_adj_651_cascade_ ;
    wire \tok.n13 ;
    wire n15_cascade_;
    wire \tok.n6_adj_687_cascade_ ;
    wire \tok.n4_adj_641 ;
    wire \tok.n5 ;
    wire \tok.n796_cascade_ ;
    wire \tok.n12 ;
    wire \tok.n796 ;
    wire \tok.n2702 ;
    wire \tok.uart_stall ;
    wire \tok.n6203 ;
    wire \tok.search_clk_N_137 ;
    wire \tok.n31_adj_637_cascade_ ;
    wire \tok.n6170 ;
    wire \tok.n30 ;
    wire \tok.n221_adj_753_cascade_ ;
    wire \tok.key_rd_3 ;
    wire \tok.key_rd_5 ;
    wire \tok.key_rd_8 ;
    wire \tok.n20_cascade_ ;
    wire \tok.n26_adj_645 ;
    wire \tok.key_rd_13 ;
    wire \tok.n14_adj_644 ;
    wire bfn_5_8_0_;
    wire \tok.n4782 ;
    wire \tok.n4783 ;
    wire \tok.n127 ;
    wire \tok.n4784 ;
    wire \tok.n6557 ;
    wire \tok.n4785 ;
    wire \tok.n320 ;
    wire \tok.n4786 ;
    wire \tok.n4787 ;
    wire GNDG0;
    wire \tok.n4788 ;
    wire \tok.n4788_THRU_CRY_0_THRU_CO ;
    wire \tok.n21_adj_660 ;
    wire \tok.n318 ;
    wire bfn_5_9_0_;
    wire \tok.n4789 ;
    wire \tok.n4790 ;
    wire \tok.n315 ;
    wire \tok.n4791 ;
    wire \tok.n4792 ;
    wire \tok.n313 ;
    wire \tok.n4793 ;
    wire \tok.n312 ;
    wire \tok.n295 ;
    wire \tok.n4794 ;
    wire \tok.n4795 ;
    wire \tok.n4796 ;
    wire bfn_5_10_0_;
    wire \tok.n293 ;
    wire \tok.n297 ;
    wire \tok.n310 ;
    wire \tok.n6452 ;
    wire \tok.n2579 ;
    wire \tok.n6392 ;
    wire \tok.n6421 ;
    wire \tok.n300 ;
    wire \tok.n6460 ;
    wire \tok.n161_adj_825 ;
    wire \tok.n197_adj_826 ;
    wire \tok.n18_adj_850 ;
    wire \tok.n17_adj_853 ;
    wire \tok.n31_cascade_ ;
    wire \tok.n299 ;
    wire \tok.n6446 ;
    wire \tok.n308 ;
    wire \tok.n294 ;
    wire \tok.n161_adj_667 ;
    wire \tok.n6371_cascade_ ;
    wire \tok.n248_adj_653 ;
    wire \tok.n200_adj_655_cascade_ ;
    wire \tok.n6_adj_658_cascade_ ;
    wire \tok.n6_adj_832_cascade_ ;
    wire \tok.n6383 ;
    wire \tok.n242_adj_654 ;
    wire \tok.S_13 ;
    wire \tok.S_8 ;
    wire \tok.n14_adj_844_cascade_ ;
    wire \tok.n20_adj_845 ;
    wire \tok.n26_adj_851 ;
    wire \tok.n6324_cascade_ ;
    wire \tok.n262_adj_858_cascade_ ;
    wire \tok.n268 ;
    wire \tok.n6315 ;
    wire CONSTANT_ONE_NET;
    wire CONSTANT_ONE_NET_cascade_;
    wire \tok.n239 ;
    wire sender_2;
    wire \tok.n6347 ;
    wire \tok.n197_adj_693 ;
    wire \tok.n248_adj_694_cascade_ ;
    wire \tok.n242_adj_695 ;
    wire \tok.n200_adj_696_cascade_ ;
    wire \tok.n6_adj_699_cascade_ ;
    wire bfn_6_2_0_;
    wire \tok.n4812 ;
    wire \tok.n4813 ;
    wire \tok.n4814 ;
    wire \tok.n4815 ;
    wire \tok.n4816 ;
    wire \tok.n4817 ;
    wire \tok.n4818 ;
    wire \tok.n13_adj_760_cascade_ ;
    wire n10_adj_905_cascade_;
    wire \tok.tc_5 ;
    wire \tok.ram.n6263_cascade_ ;
    wire \tok.n1530 ;
    wire \tok.n83_adj_759_cascade_ ;
    wire \tok.n6660 ;
    wire n10_adj_905;
    wire \tok.n83_adj_764_cascade_ ;
    wire \tok.ram.n6277_cascade_ ;
    wire n10_cascade_;
    wire \tok.tc_7 ;
    wire \tok.n1635 ;
    wire \tok.n6662 ;
    wire \tok.n13_adj_790 ;
    wire n10;
    wire \tok.n5_adj_675 ;
    wire \tok.n6205_cascade_ ;
    wire \tok.n270 ;
    wire \tok.n270_cascade_ ;
    wire \tok.A_stk.tail_18 ;
    wire A_stk_delta_1;
    wire \tok.A_stk.tail_2 ;
    wire rd_15__N_300;
    wire \tok.n283_cascade_ ;
    wire \tok.n223_cascade_ ;
    wire \tok.n4_adj_752 ;
    wire \tok.n6586_cascade_ ;
    wire \tok.n226_adj_744 ;
    wire \tok.n254 ;
    wire \tok.n319 ;
    wire \tok.n6326 ;
    wire \tok.n387_cascade_ ;
    wire \tok.n254_adj_860_cascade_ ;
    wire \tok.n163 ;
    wire \tok.n256_adj_862 ;
    wire \tok.n5_adj_871 ;
    wire \tok.n6_adj_868_cascade_ ;
    wire S_0;
    wire \tok.n28 ;
    wire \tok.key_rd_11 ;
    wire \tok.key_rd_14 ;
    wire \tok.n23_adj_638 ;
    wire \tok.key_rd_15 ;
    wire \tok.key_rd_9 ;
    wire \tok.n24 ;
    wire \tok.n26_adj_781 ;
    wire \tok.n28_adj_778_cascade_ ;
    wire \tok.n25_adj_788 ;
    wire \tok.S_15 ;
    wire \tok.n6634 ;
    wire \tok.n23_adj_848 ;
    wire \tok.n21_adj_849_cascade_ ;
    wire \tok.n24_adj_846 ;
    wire \tok.n30_adj_852 ;
    wire \tok.n323 ;
    wire \tok.n22_adj_847 ;
    wire \tok.n27_adj_782 ;
    wire \tok.n298 ;
    wire \tok.n161_adj_870 ;
    wire \tok.n6429_cascade_ ;
    wire \tok.n197_adj_872_cascade_ ;
    wire \tok.n248_adj_873 ;
    wire \tok.n296 ;
    wire \tok.n6400_cascade_ ;
    wire \tok.n161 ;
    wire \tok.n6406 ;
    wire \tok.n6415 ;
    wire \tok.n161_adj_882_cascade_ ;
    wire \tok.n208_adj_857 ;
    wire \tok.n6328 ;
    wire \tok.n250 ;
    wire \tok.n190_adj_774_cascade_ ;
    wire \tok.n6514 ;
    wire \tok.n833_cascade_ ;
    wire \tok.n6515 ;
    wire \tok.n6534_cascade_ ;
    wire \tok.n252_adj_783_cascade_ ;
    wire \tok.n255_adj_775 ;
    wire \tok.n190_adj_774 ;
    wire \tok.n258_adj_780 ;
    wire \tok.n177_adj_779 ;
    wire \tok.n6368 ;
    wire \tok.n197_adj_668 ;
    wire \tok.n248_adj_669_cascade_ ;
    wire \tok.n242_adj_670 ;
    wire \tok.n200_adj_671_cascade_ ;
    wire \tok.S_14 ;
    wire \tok.n6_adj_674_cascade_ ;
    wire \tok.table_rd_8 ;
    wire \tok.n7269 ;
    wire \tok.n203_adj_822_cascade_ ;
    wire \tok.n212_adj_824_cascade_ ;
    wire \tok.n6457_cascade_ ;
    wire \tok.n248_adj_827 ;
    wire \tok.n242_adj_828_cascade_ ;
    wire \tok.n200_adj_829 ;
    wire \tok.n231 ;
    wire \tok.n242_adj_885 ;
    wire \tok.n200_adj_886_cascade_ ;
    wire \tok.n6_adj_889_cascade_ ;
    wire \tok.n8_cascade_ ;
    wire \tok.S_11 ;
    wire \tok.n197_adj_883 ;
    wire \tok.n248_adj_884 ;
    wire \tok.n83_adj_756_cascade_ ;
    wire \tok.ram.n6260_cascade_ ;
    wire \tok.n6295 ;
    wire \tok.n1565_cascade_ ;
    wire \tok.n13_adj_757_cascade_ ;
    wire n10_adj_906_cascade_;
    wire \tok.tc_4 ;
    wire n10_adj_906;
    wire \tok.n324_cascade_ ;
    wire \tok.n225_adj_678 ;
    wire \tok.n225_adj_678_cascade_ ;
    wire \tok.n6351 ;
    wire \tok.n6632 ;
    wire \tok.n7456_cascade_ ;
    wire \tok.n176 ;
    wire \tok.n8_adj_686 ;
    wire \tok.n6622 ;
    wire \tok.n237_adj_724_cascade_ ;
    wire \tok.n4893 ;
    wire \tok.n286 ;
    wire \tok.n286_cascade_ ;
    wire \tok.n877 ;
    wire \tok.n394_cascade_ ;
    wire \tok.n6143 ;
    wire \tok.tc_3 ;
    wire \tok.tc_1 ;
    wire n92_adj_897;
    wire \tok.tc_0 ;
    wire stall_;
    wire \tok.tc_2 ;
    wire \tok.n6140 ;
    wire \tok.n6582 ;
    wire \tok.table_wr_data_5 ;
    wire \tok.n199_cascade_ ;
    wire \tok.n262 ;
    wire \tok.n4_adj_648_cascade_ ;
    wire \tok.n326 ;
    wire \tok.n234 ;
    wire \tok.table_rd_5 ;
    wire \tok.n4842_cascade_ ;
    wire \tok.n7451_cascade_ ;
    wire \tok.n6616 ;
    wire \tok.S_2 ;
    wire \tok.n164 ;
    wire \tok.n6597 ;
    wire \tok.n4_adj_711 ;
    wire \tok.n307 ;
    wire \tok.n6397 ;
    wire \tok.n242_cascade_ ;
    wire \tok.n197 ;
    wire \tok.n248 ;
    wire \tok.n6606_cascade_ ;
    wire \tok.n200 ;
    wire \tok.n6_cascade_ ;
    wire \tok.S_12 ;
    wire \tok.n200_adj_875 ;
    wire \tok.n6_adj_878_cascade_ ;
    wire \tok.S_10 ;
    wire \tok.n2600_cascade_ ;
    wire \tok.n6610_cascade_ ;
    wire \tok.n6344 ;
    wire \tok.n269_cascade_ ;
    wire \tok.n4_adj_786 ;
    wire \tok.n205_adj_789 ;
    wire \tok.n4_adj_635 ;
    wire \tok.n6341_cascade_ ;
    wire \tok.n170 ;
    wire \tok.n321 ;
    wire \tok.n4_adj_640 ;
    wire \tok.n4_adj_680 ;
    wire \tok.n239_adj_679 ;
    wire \tok.n238_adj_681_cascade_ ;
    wire \tok.n900 ;
    wire \tok.n317_adj_659 ;
    wire \tok.n2663 ;
    wire \tok.uart.sender_5 ;
    wire \tok.uart.sender_4 ;
    wire \tok.uart.sender_3 ;
    wire \tok.n2602 ;
    wire \tok.n6450 ;
    wire \tok.n215_adj_830_cascade_ ;
    wire \tok.n6605_cascade_ ;
    wire \tok.n6604 ;
    wire \tok.n6456 ;
    wire \tok.n179_adj_831 ;
    wire \tok.n214 ;
    wire \tok.n6462_cascade_ ;
    wire \tok.n786 ;
    wire \tok.n206_adj_823 ;
    wire \tok.n314 ;
    wire \tok.n6425 ;
    wire \tok.n6346 ;
    wire \tok.n215_adj_876 ;
    wire \tok.n179_adj_877 ;
    wire \tok.n6553_cascade_ ;
    wire \tok.n6552 ;
    wire \tok.n179_adj_698 ;
    wire \tok.n6537 ;
    wire \tok.n6541_cascade_ ;
    wire \tok.n6540 ;
    wire \tok.n6367 ;
    wire \tok.n179_adj_673 ;
    wire tc_plus_1_0;
    wire \tok.C_stk.n6230_cascade_ ;
    wire tc_0;
    wire c_stk_r_0;
    wire \tok.C_stk.tail_0 ;
    wire \tok.tc_plus_1_4 ;
    wire \tok.C_stk.n6239_cascade_ ;
    wire tc_4;
    wire \tok.c_stk_r_4 ;
    wire \tok.C_stk.tail_4 ;
    wire \tok.tail_12 ;
    wire \tok.C_stk.tail_20 ;
    wire \tok.tail_28 ;
    wire \tok.C_stk.tail_36 ;
    wire \tok.n83_adj_723_cascade_ ;
    wire n10_adj_908;
    wire \tok.n4_adj_726_cascade_ ;
    wire \tok.ram.n6257_cascade_ ;
    wire \tok.n6664 ;
    wire \tok.n1600_cascade_ ;
    wire \tok.n13_adj_742 ;
    wire \tok.n6301_cascade_ ;
    wire \tok.n80_adj_751_cascade_ ;
    wire \tok.n83_adj_746_cascade_ ;
    wire \tok.n6297 ;
    wire \tok.n89_adj_754 ;
    wire n92_adj_898;
    wire \tok.table_rd_3 ;
    wire \tok.n14_adj_683_cascade_ ;
    wire \tok.n9_adj_651 ;
    wire \tok.n15_adj_807_cascade_ ;
    wire \tok.n903 ;
    wire \tok.n14_adj_683 ;
    wire \tok.n6621 ;
    wire \tok.n241_adj_747 ;
    wire \tok.n6593 ;
    wire \tok.n236 ;
    wire \tok.n4925 ;
    wire \tok.n288 ;
    wire \tok.n2613 ;
    wire \tok.n6578_cascade_ ;
    wire \tok.n6581 ;
    wire \tok.n4_adj_739 ;
    wire \tok.n2611 ;
    wire \tok.n6580 ;
    wire \tok.n4_adj_684 ;
    wire \tok.n6620_cascade_ ;
    wire \tok.n311_adj_721 ;
    wire \tok.n167_cascade_ ;
    wire \tok.n6567 ;
    wire \tok.table_rd_2 ;
    wire \tok.n209_cascade_ ;
    wire \tok.n6625_cascade_ ;
    wire \tok.n6624 ;
    wire \tok.n168_adj_700_cascade_ ;
    wire \tok.n6569 ;
    wire \tok.n2548 ;
    wire \tok.n6396 ;
    wire \tok.n179_cascade_ ;
    wire \tok.n6546 ;
    wire \tok.table_rd_7 ;
    wire \tok.table_rd_4 ;
    wire \tok.n258_adj_814 ;
    wire \tok.n252_adj_815_cascade_ ;
    wire \tok.n232 ;
    wire \tok.n255_adj_808 ;
    wire \tok.n210_adj_816 ;
    wire \tok.n872_cascade_ ;
    wire \tok.n174_adj_817_cascade_ ;
    wire \tok.n4_adj_818 ;
    wire \tok.n205_adj_820 ;
    wire \tok.n200_adj_840 ;
    wire \tok.n6_adj_843_cascade_ ;
    wire \tok.S_9 ;
    wire \tok.n6440_cascade_ ;
    wire \tok.n6612_cascade_ ;
    wire \tok.n6365 ;
    wire \tok.n215_adj_672 ;
    wire \tok.n252 ;
    wire \tok.n4_adj_769_cascade_ ;
    wire \tok.n205_adj_770 ;
    wire \tok.n235 ;
    wire \tok.n190_cascade_ ;
    wire \tok.n190 ;
    wire \tok.n255_cascade_ ;
    wire \tok.n258 ;
    wire \tok.n6508_cascade_ ;
    wire \tok.n6532 ;
    wire \tok.n207_adj_771_cascade_ ;
    wire \tok.n6583 ;
    wire \tok.S_5 ;
    wire \tok.n213 ;
    wire \tok.n207_adj_776_cascade_ ;
    wire \tok.n6529_cascade_ ;
    wire \tok.n210_adj_784 ;
    wire \tok.n174_adj_785 ;
    wire \tok.n229_adj_861 ;
    wire \tok.n6320 ;
    wire \tok.n49 ;
    wire \tok.n6380_cascade_ ;
    wire \tok.n215_adj_656_cascade_ ;
    wire \tok.n2665 ;
    wire \tok.n4_adj_719 ;
    wire \tok.n4_adj_719_cascade_ ;
    wire \tok.n10_adj_809 ;
    wire \tok.n6411 ;
    wire \tok.n6404_cascade_ ;
    wire \tok.n179_adj_888 ;
    wire \tok.n6550_cascade_ ;
    wire \tok.n6549 ;
    wire \tok.n6419 ;
    wire \tok.n215_adj_697 ;
    wire \tok.n6337_cascade_ ;
    wire \tok.n6538 ;
    wire \tok.tc_plus_1_5 ;
    wire \tok.C_stk.n6236_cascade_ ;
    wire tc_5;
    wire \tok.c_stk_r_5 ;
    wire \tok.C_stk.tail_5 ;
    wire \tok.tail_13 ;
    wire \tok.C_stk.tail_21 ;
    wire \tok.tail_29 ;
    wire \tok.C_stk.tail_37 ;
    wire \tok.tc_plus_1_2 ;
    wire \tok.C_stk.n6245_cascade_ ;
    wire tc_2;
    wire \tok.c_stk_r_2 ;
    wire \tok.C_stk.tail_2 ;
    wire \tok.tail_10 ;
    wire \tok.C_stk.tail_18 ;
    wire \tok.tail_26 ;
    wire \tok.C_stk.tail_34 ;
    wire \tok.tc_plus_1_3 ;
    wire \tok.C_stk.n6242_cascade_ ;
    wire tc_3;
    wire \tok.c_stk_r_3 ;
    wire \tok.C_stk.tail_3 ;
    wire \tok.C_stk.tail_11 ;
    wire \tok.C_stk.tail_19 ;
    wire \tok.C_stk.tail_27 ;
    wire \tok.C_stk.tail_35 ;
    wire \tok.n4_adj_726 ;
    wire \tok.tc__7__N_133 ;
    wire \tok.n2573 ;
    wire \tok.n6291_cascade_ ;
    wire \tok.n80_adj_735_cascade_ ;
    wire \tok.n83_adj_725_cascade_ ;
    wire \tok.n6287 ;
    wire \tok.n89_adj_736 ;
    wire n92;
    wire \tok.n4926 ;
    wire \tok.n2692_cascade_ ;
    wire \tok.n217 ;
    wire \tok.n7154 ;
    wire \tok.n6_adj_701 ;
    wire \tok.n2700 ;
    wire \tok.n236_adj_737 ;
    wire \tok.n239_adj_738 ;
    wire \tok.n17 ;
    wire \tok.n5_adj_821 ;
    wire \tok.n2679 ;
    wire \tok.n17_cascade_ ;
    wire \tok.n864 ;
    wire \tok.n186 ;
    wire \tok.n6562_cascade_ ;
    wire \tok.n338 ;
    wire \tok.n162 ;
    wire \tok.n179_adj_730 ;
    wire \tok.n197_adj_729_cascade_ ;
    wire \tok.n7458 ;
    wire \tok.n2544 ;
    wire \tok.table_rd_1 ;
    wire \tok.n7475_cascade_ ;
    wire \tok.n237 ;
    wire \tok.n180 ;
    wire \tok.n6628 ;
    wire \tok.S_3 ;
    wire \tok.n241 ;
    wire \tok.n6637 ;
    wire \tok.n284_cascade_ ;
    wire \tok.n244_cascade_ ;
    wire \tok.n4_adj_720_cascade_ ;
    wire \tok.n145 ;
    wire \tok.n251 ;
    wire \tok.n2557 ;
    wire \tok.n4_adj_714_cascade_ ;
    wire \tok.n218 ;
    wire \tok.n39 ;
    wire \tok.n6269_cascade_ ;
    wire \tok.n6466 ;
    wire \tok.n6467 ;
    wire \tok.n6486 ;
    wire \tok.n833 ;
    wire \tok.n6490 ;
    wire \tok.n6491 ;
    wire S_1;
    wire \tok.n208 ;
    wire \tok.n6589 ;
    wire \tok.n239_adj_727 ;
    wire \tok.n6_adj_728_cascade_ ;
    wire \tok.n200_adj_732_cascade_ ;
    wire \tok.n203_adj_731 ;
    wire \tok.n6_adj_733 ;
    wire \tok.n206_adj_794 ;
    wire \tok.n207_adj_811_cascade_ ;
    wire \tok.n6481 ;
    wire \tok.n6484 ;
    wire \tok.n213_adj_810 ;
    wire \tok.S_4 ;
    wire \tok.n207_cascade_ ;
    wire \tok.n210 ;
    wire \tok.n6572_cascade_ ;
    wire \tok.n174_adj_768 ;
    wire \tok.n31 ;
    wire \tok.n26_adj_763 ;
    wire \tok.n26_adj_763_cascade_ ;
    wire \tok.n4_adj_636 ;
    wire \tok.n213_adj_795 ;
    wire \tok.n207_adj_796_cascade_ ;
    wire \tok.n872 ;
    wire \tok.n6505_cascade_ ;
    wire \tok.n42 ;
    wire \tok.n6360 ;
    wire \tok.table_rd_6 ;
    wire \tok.n210_adj_802 ;
    wire \tok.n316 ;
    wire \tok.n6409_cascade_ ;
    wire \tok.n46 ;
    wire \tok.n215_adj_887 ;
    wire \tok.n6442 ;
    wire \tok.n6433_cascade_ ;
    wire \tok.n215_adj_841 ;
    wire \tok.n179_adj_842 ;
    wire \tok.n6602_cascade_ ;
    wire \tok.n6601 ;
    wire \tok.n6375 ;
    wire \tok.n847 ;
    wire \tok.n6544 ;
    wire \tok.n179_adj_657_cascade_ ;
    wire \tok.n6543 ;
    wire \tok.n464 ;
    wire \tok.n8 ;
    wire \tok.n6382 ;
    wire tail_40;
    wire tail_8;
    wire \tok.C_stk.tail_32 ;
    wire \tok.C_stk.tail_16 ;
    wire tail_24;
    wire \tok.C_stk.tail_43 ;
    wire \tok.tail_45 ;
    wire \tok.tail_44 ;
    wire \tok.tail_42 ;
    wire tail_51;
    wire tail_59;
    wire tail_48_adj_900;
    wire tail_56;
    wire C_stk_delta_1_cascade_;
    wire tail_57;
    wire \tok.tail_52 ;
    wire \tok.tail_60 ;
    wire \tok.tail_62 ;
    wire \tok.n37 ;
    wire \tok.n2559 ;
    wire \tok.tail_53 ;
    wire rd_7__N_373_cascade_;
    wire \tok.tail_61 ;
    wire tc_plus_1_1;
    wire \tok.C_stk.n6248_cascade_ ;
    wire tc_1;
    wire c_stk_r_1;
    wire \tok.C_stk.tail_1 ;
    wire tail_9;
    wire \tok.C_stk.tail_17 ;
    wire tail_25;
    wire tail_49_adj_899;
    wire \tok.C_stk.tail_33 ;
    wire tail_41;
    wire \tok.n156 ;
    wire \tok.n211_adj_741_cascade_ ;
    wire \tok.n277_cascade_ ;
    wire \tok.n265 ;
    wire \tok.n6_adj_748 ;
    wire \tok.n6331 ;
    wire \tok.n238_adj_855_cascade_ ;
    wire \tok.n4_adj_859 ;
    wire \tok.n6_adj_676 ;
    wire \tok.n298_adj_856 ;
    wire \tok.n53_cascade_ ;
    wire \tok.n992 ;
    wire \tok.n2_cascade_ ;
    wire \tok.n23 ;
    wire \tok.n174_cascade_ ;
    wire \tok.stall ;
    wire \tok.n6189 ;
    wire \tok.n6_adj_722 ;
    wire \tok.n127_adj_772 ;
    wire \tok.n10_adj_773_cascade_ ;
    wire \tok.n6146_cascade_ ;
    wire \tok.n86 ;
    wire \tok.n5_adj_715 ;
    wire \tok.n369_cascade_ ;
    wire \tok.n278 ;
    wire \tok.n233_adj_716_cascade_ ;
    wire \tok.n229 ;
    wire \tok.n6156 ;
    wire \tok.n7 ;
    wire \tok.n4_adj_648 ;
    wire \tok.n2635 ;
    wire \tok.n6653_cascade_ ;
    wire \tok.n6646_cascade_ ;
    wire \tok.n6167 ;
    wire \tok.n6645 ;
    wire \tok.n247 ;
    wire \tok.n6639 ;
    wire \tok.n280 ;
    wire \tok.n6638_cascade_ ;
    wire \tok.n6636 ;
    wire \tok.n260_adj_717 ;
    wire \tok.S_6 ;
    wire \tok.n815 ;
    wire \tok.n6510 ;
    wire \tok.n177_adj_799_cascade_ ;
    wire \tok.n252_adj_801_cascade_ ;
    wire \tok.n867 ;
    wire \tok.n233 ;
    wire \tok.n5_adj_745 ;
    wire \tok.n255_adj_793_cascade_ ;
    wire \tok.n258_adj_800 ;
    wire \tok.n6183 ;
    wire \tok.n6162_cascade_ ;
    wire \tok.n865_cascade_ ;
    wire \tok.n222_cascade_ ;
    wire \tok.n245 ;
    wire \tok.n6501 ;
    wire \tok.n186_adj_798_cascade_ ;
    wire \tok.n6496 ;
    wire \tok.n194 ;
    wire \tok.n338_adj_805_cascade_ ;
    wire \tok.n6608 ;
    wire \tok.n219 ;
    wire \tok.n190_adj_792 ;
    wire \tok.n4_adj_804 ;
    wire \tok.n174_adj_803 ;
    wire \tok.n205_adj_806 ;
    wire \tok.n177_adj_813 ;
    wire \tok.n2598_cascade_ ;
    wire \tok.n45 ;
    wire \tok.n6390 ;
    wire \tok.n821 ;
    wire \tok.n215_cascade_ ;
    wire \tok.n6547 ;
    wire \tok.n4_adj_712 ;
    wire \tok.n238 ;
    wire \tok.n6650_cascade_ ;
    wire \tok.n48 ;
    wire \tok.n211_cascade_ ;
    wire \tok.n6644 ;
    wire \tok.n260_cascade_ ;
    wire \tok.n6641 ;
    wire \tok.n266_cascade_ ;
    wire \tok.n5_adj_713 ;
    wire \tok.n256 ;
    wire \tok.n4_adj_718_cascade_ ;
    wire \tok.n221 ;
    wire \tok.A_low_1 ;
    wire \tok.n2637 ;
    wire \tok.A_low_4 ;
    wire \tok.uart.sender_6 ;
    wire \tok.uart.sender_7 ;
    wire \tok.uart.sender_8 ;
    wire \tok.uart.n950 ;
    wire \tok.n274 ;
    wire \tok.n185 ;
    wire \tok.n7410 ;
    wire reset_c;
    wire \tok.tail_50 ;
    wire \tok.tail_58 ;
    wire \tok.tc_plus_1_6 ;
    wire \tok.C_stk.n6233_cascade_ ;
    wire tc_6;
    wire \tok.c_stk_r_6 ;
    wire \tok.C_stk.tail_6 ;
    wire \tok.tail_14 ;
    wire \tok.C_stk.tail_22 ;
    wire \tok.tail_30 ;
    wire \tok.tail_54 ;
    wire \tok.C_stk.tail_38 ;
    wire \tok.tail_46 ;
    wire \tok.C_stk.n449 ;
    wire \tok.n273 ;
    wire tc_7;
    wire \tok.C_stk.n6227_cascade_ ;
    wire \tok.n15 ;
    wire \tok.c_stk_r_7 ;
    wire \tok.C_stk.tail_7 ;
    wire \tok.tail_15 ;
    wire \tok.C_stk.tail_23 ;
    wire \tok.tail_31 ;
    wire \tok.C_stk.tail_39 ;
    wire \tok.tail_47 ;
    wire rd_7__N_373;
    wire \tok.tail_55 ;
    wire C_stk_delta_1;
    wire \tok.tail_63 ;
    wire n15;
    wire \tok.tc_plus_1_7 ;
    wire \tok.S_7 ;
    wire \tok.table_wr_data_7 ;
    wire uart_rx_data_4;
    wire uart_rx_data_2;
    wire uart_rx_data_1;
    wire capture_2;
    wire \tok.A_stk_delta_1__N_4 ;
    wire \tok.A_stk_delta_1__N_4_cascade_ ;
    wire \tok.n1 ;
    wire \tok.n4_adj_702_cascade_ ;
    wire \tok.n52 ;
    wire \tok.n51_cascade_ ;
    wire \tok.n50 ;
    wire \tok.n8_adj_854 ;
    wire \tok.n174 ;
    wire \tok.n4_adj_702 ;
    wire \tok.reset_N_2 ;
    wire \tok.n256_adj_749 ;
    wire \tok.n367 ;
    wire \tok.n215_adj_750 ;
    wire \tok.depth_2 ;
    wire \tok.depth_1 ;
    wire \tok.n741 ;
    wire \tok.n806 ;
    wire \tok.depth_0 ;
    wire \tok.n6213 ;
    wire \tok.n806_cascade_ ;
    wire \tok.depth_3 ;
    wire \tok.n748 ;
    wire \tok.n47 ;
    wire \tok.n6615 ;
    wire \tok.n158_cascade_ ;
    wire \tok.n6627 ;
    wire \tok.uart_stall_N_46 ;
    wire \tok.n9 ;
    wire \tok.n10 ;
    wire \tok.n10_cascade_ ;
    wire \tok.write_flag ;
    wire \tok.n14 ;
    wire \tok.uart.n10_cascade_ ;
    wire n23_cascade_;
    wire \tok.n168_adj_710_cascade_ ;
    wire \tok.A_low_6 ;
    wire \tok.n6502 ;
    wire uart_rx_data_6;
    wire \tok.n43 ;
    wire \tok.n311 ;
    wire \tok.n190_adj_797 ;
    wire \tok.n44 ;
    wire \tok.T_2 ;
    wire \tok.T_0 ;
    wire \tok.n168_adj_690 ;
    wire \tok.n6525 ;
    wire \tok.n6526_cascade_ ;
    wire \tok.n186_adj_777_cascade_ ;
    wire \tok.n338_adj_787 ;
    wire \tok.A_low_0 ;
    wire \tok.A_low_5 ;
    wire \tok.n866_cascade_ ;
    wire \tok.n6520 ;
    wire \tok.T_5 ;
    wire \tok.n317 ;
    wire \tok.n317_cascade_ ;
    wire \tok.A_low_3 ;
    wire \tok.n168 ;
    wire \tok.n5_adj_682 ;
    wire \tok.T_4 ;
    wire \tok.n6478_cascade_ ;
    wire \tok.T_6 ;
    wire \tok.n186_adj_812_cascade_ ;
    wire \tok.T_3 ;
    wire \tok.n338_adj_819 ;
    wire \tok.T_7 ;
    wire \tok.A_low_2 ;
    wire \tok.n289 ;
    wire \tok.T_1 ;
    wire \tok.n222 ;
    wire \tok.n838 ;
    wire \tok.n863_cascade_ ;
    wire \tok.n6472 ;
    wire \tok.n9_adj_677 ;
    wire \tok.n205 ;
    wire \tok.n6477 ;
    wire capture_8;
    wire uart_rx_data_7;
    wire txtick;
    wire n23;
    wire A_low_7;
    wire sender_9;
    wire capture_3;
    wire capture_5;
    wire \tok.n891 ;
    wire \tok.uart_rx_valid ;
    wire \tok.uart.n922 ;
    wire capture_7;
    wire capture_0;
    wire capture_4;
    wire rx_data_7__N_510_cascade_;
    wire uart_rx_data_3;
    wire capture_9;
    wire capture_6;
    wire uart_rx_data_5;
    wire capture_1;
    wire rx_data_7__N_510;
    wire uart_rx_data_0;
    wire \tok.uart_tx_busy ;
    wire \tok.uart.sentbits_3 ;
    wire \tok.uart.sentbits_2 ;
    wire \tok.uart.sentbits_1 ;
    wire \tok.uart.sentbits_0 ;
    wire \tok.uart.n994 ;
    wire \tok.uart.n1013 ;
    wire rx_c;
    wire \tok.uart.n4977 ;
    wire \tok.uart.n4977_cascade_ ;
    wire bfn_13_9_0_;
    wire \tok.uart.n4819 ;
    wire \tok.uart.n4820 ;
    wire \tok.uart.bytephase_3 ;
    wire \tok.uart.n4821 ;
    wire \tok.uart.bytephase_4 ;
    wire \tok.uart.n4822 ;
    wire \tok.uart.n4823 ;
    wire \tok.uart.bytephase_5 ;
    wire n4928;
    wire \tok.uart.n6_cascade_ ;
    wire n746_cascade_;
    wire bytephase_5__N_509;
    wire n974;
    wire \tok.uart.n6211 ;
    wire \tok.uart.n2356 ;
    wire \tok.uart.n809 ;
    wire \tok.uart.n2356_cascade_ ;
    wire n746;
    wire \tok.uart.bytephase_2 ;
    wire \tok.uart.bytephase_0 ;
    wire \tok.uart.bytephase_1 ;
    wire \tok.uart.n2357 ;
    wire \tok.uart.rxclkcounter_0 ;
    wire bfn_13_11_0_;
    wire \tok.uart.rxclkcounter_1 ;
    wire \tok.uart.n4824 ;
    wire \tok.uart.rxclkcounter_2 ;
    wire \tok.uart.n4825 ;
    wire \tok.uart.rxclkcounter_3 ;
    wire \tok.uart.n4826 ;
    wire \tok.uart.rxclkcounter_4 ;
    wire \tok.uart.n4827 ;
    wire \tok.uart.rxclkcounter_5 ;
    wire \tok.uart.n4828 ;
    wire \tok.uart.n4829 ;
    wire \tok.uart.rxclkcounter_6 ;
    wire _gnd_net_;
    wire clk;
    wire \tok.uart.rxclkcounter_6__N_476 ;

    defparam \tok.vals.mem1_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .WRITE_MODE=0;
    defparam \tok.vals.mem1_physical .READ_MODE=0;
    defparam \tok.vals.mem1_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \tok.vals.mem1_physical  (
            .RDATA({\tok.table_rd_15 ,\tok.table_rd_14 ,\tok.table_rd_13 ,\tok.table_rd_12 ,\tok.table_rd_11 ,\tok.table_rd_10 ,\tok.table_rd_9 ,\tok.table_rd_8 ,\tok.table_rd_7 ,\tok.table_rd_6 ,\tok.table_rd_5 ,\tok.table_rd_4 ,\tok.table_rd_3 ,\tok.table_rd_2 ,\tok.table_rd_1 ,\tok.table_rd_0 }),
            .RADDR({dangling_wire_0,dangling_wire_1,dangling_wire_2,N__14469,N__15849,N__15402,N__14700,N__15539,N__15633,N__15465,N__14532}),
            .WADDR({dangling_wire_3,dangling_wire_4,dangling_wire_5,N__14466,N__15852,N__15399,N__14697,N__15536,N__15636,N__15468,N__14529}),
            .MASK({dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .WDATA({N__14563,N__16507,N__14590,N__16477,N__16492,N__14578,N__15319,N__13384,N__28243,N__16309,N__19966,N__16294,N__16339,N__16282,N__16324,N__14389}),
            .RCLKE(),
            .RCLK(N__38468),
            .RE(N__17518),
            .WCLKE(),
            .WCLK(N__38467),
            .WE(N__14631));
    defparam \tok.keys.mem0_physical .WRITE_MODE=0;
    defparam \tok.keys.mem0_physical .READ_MODE=0;
    defparam \tok.keys.mem0_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \tok.keys.mem0_physical  (
            .RDATA({\tok.key_rd_15 ,\tok.key_rd_14 ,\tok.key_rd_13 ,\tok.key_rd_12 ,\tok.key_rd_11 ,\tok.key_rd_10 ,\tok.key_rd_9 ,\tok.key_rd_8 ,\tok.key_rd_7 ,\tok.key_rd_6 ,\tok.key_rd_5 ,\tok.key_rd_4 ,\tok.key_rd_3 ,\tok.key_rd_2 ,\tok.key_rd_1 ,\tok.key_rd_0 }),
            .RADDR({dangling_wire_22,dangling_wire_23,dangling_wire_24,N__14479,N__15861,N__15412,N__14710,N__15550,N__15645,N__15477,N__14542}),
            .WADDR({dangling_wire_25,dangling_wire_26,dangling_wire_27,N__14478,N__15862,N__15411,N__14709,N__15549,N__15646,N__15478,N__14541}),
            .MASK({dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .WDATA({N__24196,N__32379,N__32233,N__27043,N__24001,N__29629,N__26793,N__22255,N__37442,N__30038,N__30320,N__27388,N__36532,N__33642,N__27514,N__30511}),
            .RCLKE(),
            .RCLK(N__38455),
            .RE(N__17528),
            .WCLKE(),
            .WCLK(N__38456),
            .WE(N__14632));
    defparam \tok.ram.mem2_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010001000001000000010000000100000101010001010101000101;
    defparam \tok.ram.mem2_physical .WRITE_MODE=1;
    defparam \tok.ram.mem2_physical .READ_MODE=1;
    defparam \tok.ram.mem2_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \tok.ram.mem2_physical  (
            .RDATA({dangling_wire_44,\tok.T_7 ,dangling_wire_45,\tok.T_6 ,dangling_wire_46,\tok.T_5 ,dangling_wire_47,\tok.T_4 ,dangling_wire_48,\tok.T_3 ,dangling_wire_49,\tok.T_2 ,dangling_wire_50,\tok.T_1 ,dangling_wire_51,\tok.T_0 }),
            .RADDR({dangling_wire_52,dangling_wire_53,dangling_wire_54,N__17680,N__16438,N__17623,N__19555,N__19831,N__19669,N__19813,N__19771}),
            .WADDR({dangling_wire_55,dangling_wire_56,dangling_wire_57,N__37466,N__30065,N__30342,N__27394,N__36556,N__33645,N__27561,N__30527}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,N__37468,dangling_wire_75,N__30085,dangling_wire_76,N__30318,dangling_wire_77,N__27391,dangling_wire_78,N__36553,dangling_wire_79,N__33643,dangling_wire_80,N__27551,dangling_wire_81,N__30507}),
            .RCLKE(),
            .RCLK(N__38478),
            .RE(N__17497),
            .WCLKE(),
            .WCLK(N__38479),
            .WE(N__30169));
    defparam rx_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_pad_iopad.PULLUP=1'b0;
    IO_PAD rx_pad_iopad (
            .OE(N__38690),
            .DIN(N__38689),
            .DOUT(N__38688),
            .PACKAGEPIN(rx));
    defparam rx_pad_preio.PIN_TYPE=6'b000001;
    defparam rx_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_pad_preio (
            .PADOEN(N__38690),
            .PADOUT(N__38689),
            .PADIN(N__38688),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(rx_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam reset_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam reset_pad_iopad.PULLUP=1'b0;
    IO_PAD reset_pad_iopad (
            .OE(N__38681),
            .DIN(N__38680),
            .DOUT(N__38679),
            .PACKAGEPIN(reset));
    defparam reset_pad_preio.PIN_TYPE=6'b000001;
    defparam reset_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO reset_pad_preio (
            .PADOEN(N__38681),
            .PADOUT(N__38680),
            .PADIN(N__38679),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(reset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam tx_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_pad_iopad.PULLUP=1'b0;
    IO_PAD tx_pad_iopad (
            .OE(N__38672),
            .DIN(N__38671),
            .DOUT(N__38670),
            .PACKAGEPIN(tx));
    defparam tx_pad_preio.PIN_TYPE=6'b011001;
    defparam tx_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_pad_preio (
            .PADOEN(N__38672),
            .PADOUT(N__38671),
            .PADIN(N__38670),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14953),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__9608 (
            .O(N__38653),
            .I(N__38646));
    InMux I__9607 (
            .O(N__38652),
            .I(N__38643));
    InMux I__9606 (
            .O(N__38651),
            .I(N__38636));
    InMux I__9605 (
            .O(N__38650),
            .I(N__38636));
    InMux I__9604 (
            .O(N__38649),
            .I(N__38636));
    LocalMux I__9603 (
            .O(N__38646),
            .I(\tok.uart.bytephase_1 ));
    LocalMux I__9602 (
            .O(N__38643),
            .I(\tok.uart.bytephase_1 ));
    LocalMux I__9601 (
            .O(N__38636),
            .I(\tok.uart.bytephase_1 ));
    InMux I__9600 (
            .O(N__38629),
            .I(N__38626));
    LocalMux I__9599 (
            .O(N__38626),
            .I(N__38623));
    Odrv4 I__9598 (
            .O(N__38623),
            .I(\tok.uart.n2357 ));
    InMux I__9597 (
            .O(N__38620),
            .I(N__38616));
    InMux I__9596 (
            .O(N__38619),
            .I(N__38613));
    LocalMux I__9595 (
            .O(N__38616),
            .I(\tok.uart.rxclkcounter_0 ));
    LocalMux I__9594 (
            .O(N__38613),
            .I(\tok.uart.rxclkcounter_0 ));
    InMux I__9593 (
            .O(N__38608),
            .I(bfn_13_11_0_));
    InMux I__9592 (
            .O(N__38605),
            .I(N__38601));
    InMux I__9591 (
            .O(N__38604),
            .I(N__38598));
    LocalMux I__9590 (
            .O(N__38601),
            .I(N__38595));
    LocalMux I__9589 (
            .O(N__38598),
            .I(\tok.uart.rxclkcounter_1 ));
    Odrv4 I__9588 (
            .O(N__38595),
            .I(\tok.uart.rxclkcounter_1 ));
    InMux I__9587 (
            .O(N__38590),
            .I(\tok.uart.n4824 ));
    InMux I__9586 (
            .O(N__38587),
            .I(N__38583));
    InMux I__9585 (
            .O(N__38586),
            .I(N__38580));
    LocalMux I__9584 (
            .O(N__38583),
            .I(\tok.uart.rxclkcounter_2 ));
    LocalMux I__9583 (
            .O(N__38580),
            .I(\tok.uart.rxclkcounter_2 ));
    InMux I__9582 (
            .O(N__38575),
            .I(\tok.uart.n4825 ));
    InMux I__9581 (
            .O(N__38572),
            .I(N__38568));
    InMux I__9580 (
            .O(N__38571),
            .I(N__38565));
    LocalMux I__9579 (
            .O(N__38568),
            .I(\tok.uart.rxclkcounter_3 ));
    LocalMux I__9578 (
            .O(N__38565),
            .I(\tok.uart.rxclkcounter_3 ));
    InMux I__9577 (
            .O(N__38560),
            .I(\tok.uart.n4826 ));
    CascadeMux I__9576 (
            .O(N__38557),
            .I(N__38553));
    InMux I__9575 (
            .O(N__38556),
            .I(N__38550));
    InMux I__9574 (
            .O(N__38553),
            .I(N__38547));
    LocalMux I__9573 (
            .O(N__38550),
            .I(\tok.uart.rxclkcounter_4 ));
    LocalMux I__9572 (
            .O(N__38547),
            .I(\tok.uart.rxclkcounter_4 ));
    InMux I__9571 (
            .O(N__38542),
            .I(\tok.uart.n4827 ));
    InMux I__9570 (
            .O(N__38539),
            .I(N__38535));
    InMux I__9569 (
            .O(N__38538),
            .I(N__38532));
    LocalMux I__9568 (
            .O(N__38535),
            .I(\tok.uart.rxclkcounter_5 ));
    LocalMux I__9567 (
            .O(N__38532),
            .I(\tok.uart.rxclkcounter_5 ));
    InMux I__9566 (
            .O(N__38527),
            .I(\tok.uart.n4828 ));
    InMux I__9565 (
            .O(N__38524),
            .I(\tok.uart.n4829 ));
    InMux I__9564 (
            .O(N__38521),
            .I(N__38517));
    InMux I__9563 (
            .O(N__38520),
            .I(N__38514));
    LocalMux I__9562 (
            .O(N__38517),
            .I(\tok.uart.rxclkcounter_6 ));
    LocalMux I__9561 (
            .O(N__38514),
            .I(\tok.uart.rxclkcounter_6 ));
    ClkMux I__9560 (
            .O(N__38509),
            .I(N__38257));
    ClkMux I__9559 (
            .O(N__38508),
            .I(N__38257));
    ClkMux I__9558 (
            .O(N__38507),
            .I(N__38257));
    ClkMux I__9557 (
            .O(N__38506),
            .I(N__38257));
    ClkMux I__9556 (
            .O(N__38505),
            .I(N__38257));
    ClkMux I__9555 (
            .O(N__38504),
            .I(N__38257));
    ClkMux I__9554 (
            .O(N__38503),
            .I(N__38257));
    ClkMux I__9553 (
            .O(N__38502),
            .I(N__38257));
    ClkMux I__9552 (
            .O(N__38501),
            .I(N__38257));
    ClkMux I__9551 (
            .O(N__38500),
            .I(N__38257));
    ClkMux I__9550 (
            .O(N__38499),
            .I(N__38257));
    ClkMux I__9549 (
            .O(N__38498),
            .I(N__38257));
    ClkMux I__9548 (
            .O(N__38497),
            .I(N__38257));
    ClkMux I__9547 (
            .O(N__38496),
            .I(N__38257));
    ClkMux I__9546 (
            .O(N__38495),
            .I(N__38257));
    ClkMux I__9545 (
            .O(N__38494),
            .I(N__38257));
    ClkMux I__9544 (
            .O(N__38493),
            .I(N__38257));
    ClkMux I__9543 (
            .O(N__38492),
            .I(N__38257));
    ClkMux I__9542 (
            .O(N__38491),
            .I(N__38257));
    ClkMux I__9541 (
            .O(N__38490),
            .I(N__38257));
    ClkMux I__9540 (
            .O(N__38489),
            .I(N__38257));
    ClkMux I__9539 (
            .O(N__38488),
            .I(N__38257));
    ClkMux I__9538 (
            .O(N__38487),
            .I(N__38257));
    ClkMux I__9537 (
            .O(N__38486),
            .I(N__38257));
    ClkMux I__9536 (
            .O(N__38485),
            .I(N__38257));
    ClkMux I__9535 (
            .O(N__38484),
            .I(N__38257));
    ClkMux I__9534 (
            .O(N__38483),
            .I(N__38257));
    ClkMux I__9533 (
            .O(N__38482),
            .I(N__38257));
    ClkMux I__9532 (
            .O(N__38481),
            .I(N__38257));
    ClkMux I__9531 (
            .O(N__38480),
            .I(N__38257));
    ClkMux I__9530 (
            .O(N__38479),
            .I(N__38257));
    ClkMux I__9529 (
            .O(N__38478),
            .I(N__38257));
    ClkMux I__9528 (
            .O(N__38477),
            .I(N__38257));
    ClkMux I__9527 (
            .O(N__38476),
            .I(N__38257));
    ClkMux I__9526 (
            .O(N__38475),
            .I(N__38257));
    ClkMux I__9525 (
            .O(N__38474),
            .I(N__38257));
    ClkMux I__9524 (
            .O(N__38473),
            .I(N__38257));
    ClkMux I__9523 (
            .O(N__38472),
            .I(N__38257));
    ClkMux I__9522 (
            .O(N__38471),
            .I(N__38257));
    ClkMux I__9521 (
            .O(N__38470),
            .I(N__38257));
    ClkMux I__9520 (
            .O(N__38469),
            .I(N__38257));
    ClkMux I__9519 (
            .O(N__38468),
            .I(N__38257));
    ClkMux I__9518 (
            .O(N__38467),
            .I(N__38257));
    ClkMux I__9517 (
            .O(N__38466),
            .I(N__38257));
    ClkMux I__9516 (
            .O(N__38465),
            .I(N__38257));
    ClkMux I__9515 (
            .O(N__38464),
            .I(N__38257));
    ClkMux I__9514 (
            .O(N__38463),
            .I(N__38257));
    ClkMux I__9513 (
            .O(N__38462),
            .I(N__38257));
    ClkMux I__9512 (
            .O(N__38461),
            .I(N__38257));
    ClkMux I__9511 (
            .O(N__38460),
            .I(N__38257));
    ClkMux I__9510 (
            .O(N__38459),
            .I(N__38257));
    ClkMux I__9509 (
            .O(N__38458),
            .I(N__38257));
    ClkMux I__9508 (
            .O(N__38457),
            .I(N__38257));
    ClkMux I__9507 (
            .O(N__38456),
            .I(N__38257));
    ClkMux I__9506 (
            .O(N__38455),
            .I(N__38257));
    ClkMux I__9505 (
            .O(N__38454),
            .I(N__38257));
    ClkMux I__9504 (
            .O(N__38453),
            .I(N__38257));
    ClkMux I__9503 (
            .O(N__38452),
            .I(N__38257));
    ClkMux I__9502 (
            .O(N__38451),
            .I(N__38257));
    ClkMux I__9501 (
            .O(N__38450),
            .I(N__38257));
    ClkMux I__9500 (
            .O(N__38449),
            .I(N__38257));
    ClkMux I__9499 (
            .O(N__38448),
            .I(N__38257));
    ClkMux I__9498 (
            .O(N__38447),
            .I(N__38257));
    ClkMux I__9497 (
            .O(N__38446),
            .I(N__38257));
    ClkMux I__9496 (
            .O(N__38445),
            .I(N__38257));
    ClkMux I__9495 (
            .O(N__38444),
            .I(N__38257));
    ClkMux I__9494 (
            .O(N__38443),
            .I(N__38257));
    ClkMux I__9493 (
            .O(N__38442),
            .I(N__38257));
    ClkMux I__9492 (
            .O(N__38441),
            .I(N__38257));
    ClkMux I__9491 (
            .O(N__38440),
            .I(N__38257));
    ClkMux I__9490 (
            .O(N__38439),
            .I(N__38257));
    ClkMux I__9489 (
            .O(N__38438),
            .I(N__38257));
    ClkMux I__9488 (
            .O(N__38437),
            .I(N__38257));
    ClkMux I__9487 (
            .O(N__38436),
            .I(N__38257));
    ClkMux I__9486 (
            .O(N__38435),
            .I(N__38257));
    ClkMux I__9485 (
            .O(N__38434),
            .I(N__38257));
    ClkMux I__9484 (
            .O(N__38433),
            .I(N__38257));
    ClkMux I__9483 (
            .O(N__38432),
            .I(N__38257));
    ClkMux I__9482 (
            .O(N__38431),
            .I(N__38257));
    ClkMux I__9481 (
            .O(N__38430),
            .I(N__38257));
    ClkMux I__9480 (
            .O(N__38429),
            .I(N__38257));
    ClkMux I__9479 (
            .O(N__38428),
            .I(N__38257));
    ClkMux I__9478 (
            .O(N__38427),
            .I(N__38257));
    ClkMux I__9477 (
            .O(N__38426),
            .I(N__38257));
    GlobalMux I__9476 (
            .O(N__38257),
            .I(N__38254));
    DummyBuf I__9475 (
            .O(N__38254),
            .I(clk));
    SRMux I__9474 (
            .O(N__38251),
            .I(N__38248));
    LocalMux I__9473 (
            .O(N__38248),
            .I(N__38245));
    Span4Mux_s0_h I__9472 (
            .O(N__38245),
            .I(N__38242));
    Span4Mux_h I__9471 (
            .O(N__38242),
            .I(N__38239));
    Odrv4 I__9470 (
            .O(N__38239),
            .I(\tok.uart.rxclkcounter_6__N_476 ));
    InMux I__9469 (
            .O(N__38236),
            .I(\tok.uart.n4823 ));
    InMux I__9468 (
            .O(N__38233),
            .I(N__38228));
    InMux I__9467 (
            .O(N__38232),
            .I(N__38223));
    InMux I__9466 (
            .O(N__38231),
            .I(N__38223));
    LocalMux I__9465 (
            .O(N__38228),
            .I(\tok.uart.bytephase_5 ));
    LocalMux I__9464 (
            .O(N__38223),
            .I(\tok.uart.bytephase_5 ));
    InMux I__9463 (
            .O(N__38218),
            .I(N__38209));
    InMux I__9462 (
            .O(N__38217),
            .I(N__38209));
    InMux I__9461 (
            .O(N__38216),
            .I(N__38198));
    InMux I__9460 (
            .O(N__38215),
            .I(N__38198));
    InMux I__9459 (
            .O(N__38214),
            .I(N__38198));
    LocalMux I__9458 (
            .O(N__38209),
            .I(N__38195));
    InMux I__9457 (
            .O(N__38208),
            .I(N__38192));
    InMux I__9456 (
            .O(N__38207),
            .I(N__38185));
    InMux I__9455 (
            .O(N__38206),
            .I(N__38185));
    InMux I__9454 (
            .O(N__38205),
            .I(N__38185));
    LocalMux I__9453 (
            .O(N__38198),
            .I(N__38181));
    Span4Mux_v I__9452 (
            .O(N__38195),
            .I(N__38174));
    LocalMux I__9451 (
            .O(N__38192),
            .I(N__38174));
    LocalMux I__9450 (
            .O(N__38185),
            .I(N__38174));
    InMux I__9449 (
            .O(N__38184),
            .I(N__38171));
    Odrv12 I__9448 (
            .O(N__38181),
            .I(n4928));
    Odrv4 I__9447 (
            .O(N__38174),
            .I(n4928));
    LocalMux I__9446 (
            .O(N__38171),
            .I(n4928));
    CascadeMux I__9445 (
            .O(N__38164),
            .I(\tok.uart.n6_cascade_ ));
    CascadeMux I__9444 (
            .O(N__38161),
            .I(n746_cascade_));
    SRMux I__9443 (
            .O(N__38158),
            .I(N__38154));
    InMux I__9442 (
            .O(N__38157),
            .I(N__38151));
    LocalMux I__9441 (
            .O(N__38154),
            .I(N__38148));
    LocalMux I__9440 (
            .O(N__38151),
            .I(N__38145));
    Odrv12 I__9439 (
            .O(N__38148),
            .I(bytephase_5__N_509));
    Odrv4 I__9438 (
            .O(N__38145),
            .I(bytephase_5__N_509));
    CEMux I__9437 (
            .O(N__38140),
            .I(N__38137));
    LocalMux I__9436 (
            .O(N__38137),
            .I(n974));
    InMux I__9435 (
            .O(N__38134),
            .I(N__38131));
    LocalMux I__9434 (
            .O(N__38131),
            .I(\tok.uart.n6211 ));
    InMux I__9433 (
            .O(N__38128),
            .I(N__38125));
    LocalMux I__9432 (
            .O(N__38125),
            .I(N__38122));
    Odrv4 I__9431 (
            .O(N__38122),
            .I(\tok.uart.n2356 ));
    InMux I__9430 (
            .O(N__38119),
            .I(N__38116));
    LocalMux I__9429 (
            .O(N__38116),
            .I(N__38112));
    InMux I__9428 (
            .O(N__38115),
            .I(N__38109));
    Odrv12 I__9427 (
            .O(N__38112),
            .I(\tok.uart.n809 ));
    LocalMux I__9426 (
            .O(N__38109),
            .I(\tok.uart.n809 ));
    CascadeMux I__9425 (
            .O(N__38104),
            .I(\tok.uart.n2356_cascade_ ));
    InMux I__9424 (
            .O(N__38101),
            .I(N__38095));
    InMux I__9423 (
            .O(N__38100),
            .I(N__38095));
    LocalMux I__9422 (
            .O(N__38095),
            .I(n746));
    InMux I__9421 (
            .O(N__38092),
            .I(N__38087));
    InMux I__9420 (
            .O(N__38091),
            .I(N__38082));
    InMux I__9419 (
            .O(N__38090),
            .I(N__38082));
    LocalMux I__9418 (
            .O(N__38087),
            .I(\tok.uart.bytephase_2 ));
    LocalMux I__9417 (
            .O(N__38082),
            .I(\tok.uart.bytephase_2 ));
    CascadeMux I__9416 (
            .O(N__38077),
            .I(N__38073));
    InMux I__9415 (
            .O(N__38076),
            .I(N__38068));
    InMux I__9414 (
            .O(N__38073),
            .I(N__38061));
    InMux I__9413 (
            .O(N__38072),
            .I(N__38061));
    InMux I__9412 (
            .O(N__38071),
            .I(N__38061));
    LocalMux I__9411 (
            .O(N__38068),
            .I(\tok.uart.bytephase_0 ));
    LocalMux I__9410 (
            .O(N__38061),
            .I(\tok.uart.bytephase_0 ));
    CascadeMux I__9409 (
            .O(N__38056),
            .I(N__38052));
    CascadeMux I__9408 (
            .O(N__38055),
            .I(N__38048));
    InMux I__9407 (
            .O(N__38052),
            .I(N__38035));
    InMux I__9406 (
            .O(N__38051),
            .I(N__38035));
    InMux I__9405 (
            .O(N__38048),
            .I(N__38035));
    InMux I__9404 (
            .O(N__38047),
            .I(N__38035));
    InMux I__9403 (
            .O(N__38046),
            .I(N__38035));
    LocalMux I__9402 (
            .O(N__38035),
            .I(\tok.uart.sentbits_0 ));
    CEMux I__9401 (
            .O(N__38032),
            .I(N__38029));
    LocalMux I__9400 (
            .O(N__38029),
            .I(N__38026));
    Span4Mux_s0_h I__9399 (
            .O(N__38026),
            .I(N__38023));
    Odrv4 I__9398 (
            .O(N__38023),
            .I(\tok.uart.n994 ));
    SRMux I__9397 (
            .O(N__38020),
            .I(N__38017));
    LocalMux I__9396 (
            .O(N__38017),
            .I(N__38014));
    Odrv4 I__9395 (
            .O(N__38014),
            .I(\tok.uart.n1013 ));
    CascadeMux I__9394 (
            .O(N__38011),
            .I(N__38007));
    InMux I__9393 (
            .O(N__38010),
            .I(N__38004));
    InMux I__9392 (
            .O(N__38007),
            .I(N__38001));
    LocalMux I__9391 (
            .O(N__38004),
            .I(N__37996));
    LocalMux I__9390 (
            .O(N__38001),
            .I(N__37996));
    Span4Mux_v I__9389 (
            .O(N__37996),
            .I(N__37993));
    Span4Mux_v I__9388 (
            .O(N__37993),
            .I(N__37990));
    IoSpan4Mux I__9387 (
            .O(N__37990),
            .I(N__37987));
    Odrv4 I__9386 (
            .O(N__37987),
            .I(rx_c));
    InMux I__9385 (
            .O(N__37984),
            .I(N__37981));
    LocalMux I__9384 (
            .O(N__37981),
            .I(\tok.uart.n4977 ));
    CascadeMux I__9383 (
            .O(N__37978),
            .I(\tok.uart.n4977_cascade_ ));
    InMux I__9382 (
            .O(N__37975),
            .I(bfn_13_9_0_));
    InMux I__9381 (
            .O(N__37972),
            .I(\tok.uart.n4819 ));
    InMux I__9380 (
            .O(N__37969),
            .I(\tok.uart.n4820 ));
    CascadeMux I__9379 (
            .O(N__37966),
            .I(N__37963));
    InMux I__9378 (
            .O(N__37963),
            .I(N__37956));
    InMux I__9377 (
            .O(N__37962),
            .I(N__37956));
    InMux I__9376 (
            .O(N__37961),
            .I(N__37953));
    LocalMux I__9375 (
            .O(N__37956),
            .I(N__37950));
    LocalMux I__9374 (
            .O(N__37953),
            .I(\tok.uart.bytephase_3 ));
    Odrv4 I__9373 (
            .O(N__37950),
            .I(\tok.uart.bytephase_3 ));
    InMux I__9372 (
            .O(N__37945),
            .I(\tok.uart.n4821 ));
    InMux I__9371 (
            .O(N__37942),
            .I(N__37937));
    InMux I__9370 (
            .O(N__37941),
            .I(N__37932));
    InMux I__9369 (
            .O(N__37940),
            .I(N__37932));
    LocalMux I__9368 (
            .O(N__37937),
            .I(\tok.uart.bytephase_4 ));
    LocalMux I__9367 (
            .O(N__37932),
            .I(\tok.uart.bytephase_4 ));
    InMux I__9366 (
            .O(N__37927),
            .I(\tok.uart.n4822 ));
    InMux I__9365 (
            .O(N__37924),
            .I(N__37918));
    InMux I__9364 (
            .O(N__37923),
            .I(N__37918));
    LocalMux I__9363 (
            .O(N__37918),
            .I(capture_0));
    InMux I__9362 (
            .O(N__37915),
            .I(N__37912));
    LocalMux I__9361 (
            .O(N__37912),
            .I(N__37907));
    InMux I__9360 (
            .O(N__37911),
            .I(N__37904));
    InMux I__9359 (
            .O(N__37910),
            .I(N__37901));
    Odrv4 I__9358 (
            .O(N__37907),
            .I(capture_4));
    LocalMux I__9357 (
            .O(N__37904),
            .I(capture_4));
    LocalMux I__9356 (
            .O(N__37901),
            .I(capture_4));
    CascadeMux I__9355 (
            .O(N__37894),
            .I(rx_data_7__N_510_cascade_));
    CascadeMux I__9354 (
            .O(N__37891),
            .I(N__37888));
    InMux I__9353 (
            .O(N__37888),
            .I(N__37885));
    LocalMux I__9352 (
            .O(N__37885),
            .I(N__37881));
    InMux I__9351 (
            .O(N__37884),
            .I(N__37878));
    Span4Mux_h I__9350 (
            .O(N__37881),
            .I(N__37875));
    LocalMux I__9349 (
            .O(N__37878),
            .I(uart_rx_data_3));
    Odrv4 I__9348 (
            .O(N__37875),
            .I(uart_rx_data_3));
    InMux I__9347 (
            .O(N__37870),
            .I(N__37865));
    InMux I__9346 (
            .O(N__37869),
            .I(N__37860));
    InMux I__9345 (
            .O(N__37868),
            .I(N__37860));
    LocalMux I__9344 (
            .O(N__37865),
            .I(capture_9));
    LocalMux I__9343 (
            .O(N__37860),
            .I(capture_9));
    InMux I__9342 (
            .O(N__37855),
            .I(N__37851));
    CascadeMux I__9341 (
            .O(N__37854),
            .I(N__37848));
    LocalMux I__9340 (
            .O(N__37851),
            .I(N__37844));
    InMux I__9339 (
            .O(N__37848),
            .I(N__37839));
    InMux I__9338 (
            .O(N__37847),
            .I(N__37839));
    Odrv4 I__9337 (
            .O(N__37844),
            .I(capture_6));
    LocalMux I__9336 (
            .O(N__37839),
            .I(capture_6));
    CascadeMux I__9335 (
            .O(N__37834),
            .I(N__37831));
    InMux I__9334 (
            .O(N__37831),
            .I(N__37827));
    InMux I__9333 (
            .O(N__37830),
            .I(N__37824));
    LocalMux I__9332 (
            .O(N__37827),
            .I(N__37821));
    LocalMux I__9331 (
            .O(N__37824),
            .I(uart_rx_data_5));
    Odrv4 I__9330 (
            .O(N__37821),
            .I(uart_rx_data_5));
    InMux I__9329 (
            .O(N__37816),
            .I(N__37812));
    InMux I__9328 (
            .O(N__37815),
            .I(N__37809));
    LocalMux I__9327 (
            .O(N__37812),
            .I(N__37803));
    LocalMux I__9326 (
            .O(N__37809),
            .I(N__37803));
    InMux I__9325 (
            .O(N__37808),
            .I(N__37800));
    Odrv4 I__9324 (
            .O(N__37803),
            .I(capture_1));
    LocalMux I__9323 (
            .O(N__37800),
            .I(capture_1));
    InMux I__9322 (
            .O(N__37795),
            .I(N__37792));
    LocalMux I__9321 (
            .O(N__37792),
            .I(N__37784));
    InMux I__9320 (
            .O(N__37791),
            .I(N__37781));
    InMux I__9319 (
            .O(N__37790),
            .I(N__37772));
    InMux I__9318 (
            .O(N__37789),
            .I(N__37772));
    InMux I__9317 (
            .O(N__37788),
            .I(N__37772));
    InMux I__9316 (
            .O(N__37787),
            .I(N__37769));
    Span4Mux_v I__9315 (
            .O(N__37784),
            .I(N__37764));
    LocalMux I__9314 (
            .O(N__37781),
            .I(N__37764));
    InMux I__9313 (
            .O(N__37780),
            .I(N__37759));
    InMux I__9312 (
            .O(N__37779),
            .I(N__37759));
    LocalMux I__9311 (
            .O(N__37772),
            .I(N__37754));
    LocalMux I__9310 (
            .O(N__37769),
            .I(N__37754));
    Odrv4 I__9309 (
            .O(N__37764),
            .I(rx_data_7__N_510));
    LocalMux I__9308 (
            .O(N__37759),
            .I(rx_data_7__N_510));
    Odrv4 I__9307 (
            .O(N__37754),
            .I(rx_data_7__N_510));
    CascadeMux I__9306 (
            .O(N__37747),
            .I(N__37744));
    InMux I__9305 (
            .O(N__37744),
            .I(N__37741));
    LocalMux I__9304 (
            .O(N__37741),
            .I(N__37738));
    Span4Mux_h I__9303 (
            .O(N__37738),
            .I(N__37734));
    InMux I__9302 (
            .O(N__37737),
            .I(N__37731));
    Span4Mux_h I__9301 (
            .O(N__37734),
            .I(N__37728));
    LocalMux I__9300 (
            .O(N__37731),
            .I(uart_rx_data_0));
    Odrv4 I__9299 (
            .O(N__37728),
            .I(uart_rx_data_0));
    InMux I__9298 (
            .O(N__37723),
            .I(N__37711));
    InMux I__9297 (
            .O(N__37722),
            .I(N__37711));
    InMux I__9296 (
            .O(N__37721),
            .I(N__37711));
    InMux I__9295 (
            .O(N__37720),
            .I(N__37711));
    LocalMux I__9294 (
            .O(N__37711),
            .I(\tok.uart_tx_busy ));
    InMux I__9293 (
            .O(N__37708),
            .I(N__37702));
    InMux I__9292 (
            .O(N__37707),
            .I(N__37702));
    LocalMux I__9291 (
            .O(N__37702),
            .I(\tok.uart.sentbits_3 ));
    CascadeMux I__9290 (
            .O(N__37699),
            .I(N__37694));
    InMux I__9289 (
            .O(N__37698),
            .I(N__37687));
    InMux I__9288 (
            .O(N__37697),
            .I(N__37687));
    InMux I__9287 (
            .O(N__37694),
            .I(N__37687));
    LocalMux I__9286 (
            .O(N__37687),
            .I(\tok.uart.sentbits_2 ));
    InMux I__9285 (
            .O(N__37684),
            .I(N__37672));
    InMux I__9284 (
            .O(N__37683),
            .I(N__37672));
    InMux I__9283 (
            .O(N__37682),
            .I(N__37672));
    InMux I__9282 (
            .O(N__37681),
            .I(N__37672));
    LocalMux I__9281 (
            .O(N__37672),
            .I(\tok.uart.sentbits_1 ));
    InMux I__9280 (
            .O(N__37669),
            .I(N__37665));
    InMux I__9279 (
            .O(N__37668),
            .I(N__37662));
    LocalMux I__9278 (
            .O(N__37665),
            .I(N__37658));
    LocalMux I__9277 (
            .O(N__37662),
            .I(N__37655));
    InMux I__9276 (
            .O(N__37661),
            .I(N__37652));
    Odrv12 I__9275 (
            .O(N__37658),
            .I(capture_8));
    Odrv4 I__9274 (
            .O(N__37655),
            .I(capture_8));
    LocalMux I__9273 (
            .O(N__37652),
            .I(capture_8));
    CascadeMux I__9272 (
            .O(N__37645),
            .I(N__37642));
    InMux I__9271 (
            .O(N__37642),
            .I(N__37638));
    InMux I__9270 (
            .O(N__37641),
            .I(N__37635));
    LocalMux I__9269 (
            .O(N__37638),
            .I(N__37632));
    LocalMux I__9268 (
            .O(N__37635),
            .I(uart_rx_data_7));
    Odrv4 I__9267 (
            .O(N__37632),
            .I(uart_rx_data_7));
    InMux I__9266 (
            .O(N__37627),
            .I(N__37624));
    LocalMux I__9265 (
            .O(N__37624),
            .I(N__37620));
    CascadeMux I__9264 (
            .O(N__37623),
            .I(N__37617));
    Span4Mux_s2_v I__9263 (
            .O(N__37620),
            .I(N__37613));
    InMux I__9262 (
            .O(N__37617),
            .I(N__37608));
    InMux I__9261 (
            .O(N__37616),
            .I(N__37608));
    Span4Mux_v I__9260 (
            .O(N__37613),
            .I(N__37602));
    LocalMux I__9259 (
            .O(N__37608),
            .I(N__37602));
    SRMux I__9258 (
            .O(N__37607),
            .I(N__37598));
    Span4Mux_h I__9257 (
            .O(N__37602),
            .I(N__37595));
    SRMux I__9256 (
            .O(N__37601),
            .I(N__37592));
    LocalMux I__9255 (
            .O(N__37598),
            .I(N__37588));
    Span4Mux_h I__9254 (
            .O(N__37595),
            .I(N__37585));
    LocalMux I__9253 (
            .O(N__37592),
            .I(N__37582));
    InMux I__9252 (
            .O(N__37591),
            .I(N__37579));
    Span4Mux_s2_v I__9251 (
            .O(N__37588),
            .I(N__37574));
    Span4Mux_h I__9250 (
            .O(N__37585),
            .I(N__37574));
    Odrv4 I__9249 (
            .O(N__37582),
            .I(txtick));
    LocalMux I__9248 (
            .O(N__37579),
            .I(txtick));
    Odrv4 I__9247 (
            .O(N__37574),
            .I(txtick));
    CascadeMux I__9246 (
            .O(N__37567),
            .I(N__37562));
    SRMux I__9245 (
            .O(N__37566),
            .I(N__37558));
    InMux I__9244 (
            .O(N__37565),
            .I(N__37549));
    InMux I__9243 (
            .O(N__37562),
            .I(N__37549));
    InMux I__9242 (
            .O(N__37561),
            .I(N__37549));
    LocalMux I__9241 (
            .O(N__37558),
            .I(N__37546));
    InMux I__9240 (
            .O(N__37557),
            .I(N__37541));
    InMux I__9239 (
            .O(N__37556),
            .I(N__37541));
    LocalMux I__9238 (
            .O(N__37549),
            .I(N__37537));
    Span4Mux_s2_v I__9237 (
            .O(N__37546),
            .I(N__37529));
    LocalMux I__9236 (
            .O(N__37541),
            .I(N__37529));
    InMux I__9235 (
            .O(N__37540),
            .I(N__37526));
    Span4Mux_v I__9234 (
            .O(N__37537),
            .I(N__37523));
    InMux I__9233 (
            .O(N__37536),
            .I(N__37516));
    InMux I__9232 (
            .O(N__37535),
            .I(N__37516));
    InMux I__9231 (
            .O(N__37534),
            .I(N__37516));
    Span4Mux_v I__9230 (
            .O(N__37529),
            .I(N__37512));
    LocalMux I__9229 (
            .O(N__37526),
            .I(N__37509));
    Span4Mux_h I__9228 (
            .O(N__37523),
            .I(N__37504));
    LocalMux I__9227 (
            .O(N__37516),
            .I(N__37504));
    InMux I__9226 (
            .O(N__37515),
            .I(N__37501));
    Span4Mux_h I__9225 (
            .O(N__37512),
            .I(N__37497));
    Span12Mux_h I__9224 (
            .O(N__37509),
            .I(N__37490));
    Sp12to4 I__9223 (
            .O(N__37504),
            .I(N__37490));
    LocalMux I__9222 (
            .O(N__37501),
            .I(N__37490));
    InMux I__9221 (
            .O(N__37500),
            .I(N__37487));
    Span4Mux_h I__9220 (
            .O(N__37497),
            .I(N__37484));
    Odrv12 I__9219 (
            .O(N__37490),
            .I(n23));
    LocalMux I__9218 (
            .O(N__37487),
            .I(n23));
    Odrv4 I__9217 (
            .O(N__37484),
            .I(n23));
    InMux I__9216 (
            .O(N__37477),
            .I(N__37471));
    InMux I__9215 (
            .O(N__37476),
            .I(N__37460));
    InMux I__9214 (
            .O(N__37475),
            .I(N__37460));
    InMux I__9213 (
            .O(N__37474),
            .I(N__37457));
    LocalMux I__9212 (
            .O(N__37471),
            .I(N__37452));
    InMux I__9211 (
            .O(N__37470),
            .I(N__37449));
    CascadeMux I__9210 (
            .O(N__37469),
            .I(N__37446));
    InMux I__9209 (
            .O(N__37468),
            .I(N__37439));
    InMux I__9208 (
            .O(N__37467),
            .I(N__37436));
    CascadeMux I__9207 (
            .O(N__37466),
            .I(N__37433));
    InMux I__9206 (
            .O(N__37465),
            .I(N__37430));
    LocalMux I__9205 (
            .O(N__37460),
            .I(N__37427));
    LocalMux I__9204 (
            .O(N__37457),
            .I(N__37424));
    InMux I__9203 (
            .O(N__37456),
            .I(N__37419));
    InMux I__9202 (
            .O(N__37455),
            .I(N__37419));
    Span4Mux_s0_v I__9201 (
            .O(N__37452),
            .I(N__37416));
    LocalMux I__9200 (
            .O(N__37449),
            .I(N__37413));
    InMux I__9199 (
            .O(N__37446),
            .I(N__37406));
    InMux I__9198 (
            .O(N__37445),
            .I(N__37406));
    InMux I__9197 (
            .O(N__37444),
            .I(N__37406));
    InMux I__9196 (
            .O(N__37443),
            .I(N__37403));
    InMux I__9195 (
            .O(N__37442),
            .I(N__37397));
    LocalMux I__9194 (
            .O(N__37439),
            .I(N__37394));
    LocalMux I__9193 (
            .O(N__37436),
            .I(N__37391));
    InMux I__9192 (
            .O(N__37433),
            .I(N__37388));
    LocalMux I__9191 (
            .O(N__37430),
            .I(N__37383));
    Span4Mux_s1_h I__9190 (
            .O(N__37427),
            .I(N__37380));
    Span4Mux_s3_v I__9189 (
            .O(N__37424),
            .I(N__37375));
    LocalMux I__9188 (
            .O(N__37419),
            .I(N__37375));
    Span4Mux_v I__9187 (
            .O(N__37416),
            .I(N__37372));
    Span4Mux_s1_v I__9186 (
            .O(N__37413),
            .I(N__37365));
    LocalMux I__9185 (
            .O(N__37406),
            .I(N__37365));
    LocalMux I__9184 (
            .O(N__37403),
            .I(N__37365));
    InMux I__9183 (
            .O(N__37402),
            .I(N__37360));
    InMux I__9182 (
            .O(N__37401),
            .I(N__37360));
    CascadeMux I__9181 (
            .O(N__37400),
            .I(N__37356));
    LocalMux I__9180 (
            .O(N__37397),
            .I(N__37349));
    Span4Mux_v I__9179 (
            .O(N__37394),
            .I(N__37349));
    Span4Mux_v I__9178 (
            .O(N__37391),
            .I(N__37349));
    LocalMux I__9177 (
            .O(N__37388),
            .I(N__37346));
    InMux I__9176 (
            .O(N__37387),
            .I(N__37341));
    InMux I__9175 (
            .O(N__37386),
            .I(N__37341));
    Span4Mux_s3_v I__9174 (
            .O(N__37383),
            .I(N__37334));
    Span4Mux_h I__9173 (
            .O(N__37380),
            .I(N__37334));
    Span4Mux_h I__9172 (
            .O(N__37375),
            .I(N__37334));
    Span4Mux_v I__9171 (
            .O(N__37372),
            .I(N__37329));
    Span4Mux_v I__9170 (
            .O(N__37365),
            .I(N__37329));
    LocalMux I__9169 (
            .O(N__37360),
            .I(N__37326));
    InMux I__9168 (
            .O(N__37359),
            .I(N__37321));
    InMux I__9167 (
            .O(N__37356),
            .I(N__37321));
    Span4Mux_h I__9166 (
            .O(N__37349),
            .I(N__37316));
    Span4Mux_h I__9165 (
            .O(N__37346),
            .I(N__37316));
    LocalMux I__9164 (
            .O(N__37341),
            .I(A_low_7));
    Odrv4 I__9163 (
            .O(N__37334),
            .I(A_low_7));
    Odrv4 I__9162 (
            .O(N__37329),
            .I(A_low_7));
    Odrv12 I__9161 (
            .O(N__37326),
            .I(A_low_7));
    LocalMux I__9160 (
            .O(N__37321),
            .I(A_low_7));
    Odrv4 I__9159 (
            .O(N__37316),
            .I(A_low_7));
    CascadeMux I__9158 (
            .O(N__37303),
            .I(N__37300));
    InMux I__9157 (
            .O(N__37300),
            .I(N__37296));
    InMux I__9156 (
            .O(N__37299),
            .I(N__37293));
    LocalMux I__9155 (
            .O(N__37296),
            .I(sender_9));
    LocalMux I__9154 (
            .O(N__37293),
            .I(sender_9));
    CascadeMux I__9153 (
            .O(N__37288),
            .I(N__37285));
    InMux I__9152 (
            .O(N__37285),
            .I(N__37278));
    InMux I__9151 (
            .O(N__37284),
            .I(N__37278));
    InMux I__9150 (
            .O(N__37283),
            .I(N__37275));
    LocalMux I__9149 (
            .O(N__37278),
            .I(capture_3));
    LocalMux I__9148 (
            .O(N__37275),
            .I(capture_3));
    InMux I__9147 (
            .O(N__37270),
            .I(N__37267));
    LocalMux I__9146 (
            .O(N__37267),
            .I(N__37262));
    InMux I__9145 (
            .O(N__37266),
            .I(N__37257));
    InMux I__9144 (
            .O(N__37265),
            .I(N__37257));
    Odrv4 I__9143 (
            .O(N__37262),
            .I(capture_5));
    LocalMux I__9142 (
            .O(N__37257),
            .I(capture_5));
    InMux I__9141 (
            .O(N__37252),
            .I(N__37249));
    LocalMux I__9140 (
            .O(N__37249),
            .I(N__37246));
    Span4Mux_s0_h I__9139 (
            .O(N__37246),
            .I(N__37243));
    Span4Mux_h I__9138 (
            .O(N__37243),
            .I(N__37238));
    InMux I__9137 (
            .O(N__37242),
            .I(N__37235));
    CascadeMux I__9136 (
            .O(N__37241),
            .I(N__37231));
    Span4Mux_h I__9135 (
            .O(N__37238),
            .I(N__37227));
    LocalMux I__9134 (
            .O(N__37235),
            .I(N__37224));
    InMux I__9133 (
            .O(N__37234),
            .I(N__37221));
    InMux I__9132 (
            .O(N__37231),
            .I(N__37216));
    InMux I__9131 (
            .O(N__37230),
            .I(N__37216));
    Odrv4 I__9130 (
            .O(N__37227),
            .I(\tok.n891 ));
    Odrv12 I__9129 (
            .O(N__37224),
            .I(\tok.n891 ));
    LocalMux I__9128 (
            .O(N__37221),
            .I(\tok.n891 ));
    LocalMux I__9127 (
            .O(N__37216),
            .I(\tok.n891 ));
    CascadeMux I__9126 (
            .O(N__37207),
            .I(N__37204));
    InMux I__9125 (
            .O(N__37204),
            .I(N__37195));
    InMux I__9124 (
            .O(N__37203),
            .I(N__37195));
    InMux I__9123 (
            .O(N__37202),
            .I(N__37195));
    LocalMux I__9122 (
            .O(N__37195),
            .I(N__37192));
    Span4Mux_h I__9121 (
            .O(N__37192),
            .I(N__37187));
    InMux I__9120 (
            .O(N__37191),
            .I(N__37184));
    InMux I__9119 (
            .O(N__37190),
            .I(N__37181));
    Span4Mux_h I__9118 (
            .O(N__37187),
            .I(N__37178));
    LocalMux I__9117 (
            .O(N__37184),
            .I(\tok.uart_rx_valid ));
    LocalMux I__9116 (
            .O(N__37181),
            .I(\tok.uart_rx_valid ));
    Odrv4 I__9115 (
            .O(N__37178),
            .I(\tok.uart_rx_valid ));
    CEMux I__9114 (
            .O(N__37171),
            .I(N__37168));
    LocalMux I__9113 (
            .O(N__37168),
            .I(N__37165));
    Sp12to4 I__9112 (
            .O(N__37165),
            .I(N__37162));
    Odrv12 I__9111 (
            .O(N__37162),
            .I(\tok.uart.n922 ));
    InMux I__9110 (
            .O(N__37159),
            .I(N__37156));
    LocalMux I__9109 (
            .O(N__37156),
            .I(N__37153));
    Span4Mux_v I__9108 (
            .O(N__37153),
            .I(N__37148));
    InMux I__9107 (
            .O(N__37152),
            .I(N__37143));
    InMux I__9106 (
            .O(N__37151),
            .I(N__37143));
    Odrv4 I__9105 (
            .O(N__37148),
            .I(capture_7));
    LocalMux I__9104 (
            .O(N__37143),
            .I(capture_7));
    CascadeMux I__9103 (
            .O(N__37138),
            .I(N__37131));
    InMux I__9102 (
            .O(N__37137),
            .I(N__37117));
    InMux I__9101 (
            .O(N__37136),
            .I(N__37117));
    CascadeMux I__9100 (
            .O(N__37135),
            .I(N__37114));
    InMux I__9099 (
            .O(N__37134),
            .I(N__37107));
    InMux I__9098 (
            .O(N__37131),
            .I(N__37100));
    InMux I__9097 (
            .O(N__37130),
            .I(N__37100));
    InMux I__9096 (
            .O(N__37129),
            .I(N__37100));
    CascadeMux I__9095 (
            .O(N__37128),
            .I(N__37088));
    InMux I__9094 (
            .O(N__37127),
            .I(N__37079));
    CascadeMux I__9093 (
            .O(N__37126),
            .I(N__37070));
    InMux I__9092 (
            .O(N__37125),
            .I(N__37058));
    InMux I__9091 (
            .O(N__37124),
            .I(N__37058));
    InMux I__9090 (
            .O(N__37123),
            .I(N__37053));
    InMux I__9089 (
            .O(N__37122),
            .I(N__37053));
    LocalMux I__9088 (
            .O(N__37117),
            .I(N__37050));
    InMux I__9087 (
            .O(N__37114),
            .I(N__37047));
    InMux I__9086 (
            .O(N__37113),
            .I(N__37039));
    InMux I__9085 (
            .O(N__37112),
            .I(N__37034));
    InMux I__9084 (
            .O(N__37111),
            .I(N__37034));
    InMux I__9083 (
            .O(N__37110),
            .I(N__37031));
    LocalMux I__9082 (
            .O(N__37107),
            .I(N__37026));
    LocalMux I__9081 (
            .O(N__37100),
            .I(N__37026));
    CascadeMux I__9080 (
            .O(N__37099),
            .I(N__37023));
    InMux I__9079 (
            .O(N__37098),
            .I(N__37018));
    InMux I__9078 (
            .O(N__37097),
            .I(N__37018));
    InMux I__9077 (
            .O(N__37096),
            .I(N__37011));
    InMux I__9076 (
            .O(N__37095),
            .I(N__37011));
    InMux I__9075 (
            .O(N__37094),
            .I(N__37011));
    InMux I__9074 (
            .O(N__37093),
            .I(N__37004));
    InMux I__9073 (
            .O(N__37092),
            .I(N__37004));
    InMux I__9072 (
            .O(N__37091),
            .I(N__37004));
    InMux I__9071 (
            .O(N__37088),
            .I(N__36994));
    InMux I__9070 (
            .O(N__37087),
            .I(N__36994));
    InMux I__9069 (
            .O(N__37086),
            .I(N__36994));
    InMux I__9068 (
            .O(N__37085),
            .I(N__36989));
    InMux I__9067 (
            .O(N__37084),
            .I(N__36989));
    InMux I__9066 (
            .O(N__37083),
            .I(N__36973));
    InMux I__9065 (
            .O(N__37082),
            .I(N__36973));
    LocalMux I__9064 (
            .O(N__37079),
            .I(N__36970));
    InMux I__9063 (
            .O(N__37078),
            .I(N__36959));
    InMux I__9062 (
            .O(N__37077),
            .I(N__36959));
    InMux I__9061 (
            .O(N__37076),
            .I(N__36959));
    InMux I__9060 (
            .O(N__37075),
            .I(N__36959));
    InMux I__9059 (
            .O(N__37074),
            .I(N__36959));
    InMux I__9058 (
            .O(N__37073),
            .I(N__36942));
    InMux I__9057 (
            .O(N__37070),
            .I(N__36937));
    InMux I__9056 (
            .O(N__37069),
            .I(N__36937));
    InMux I__9055 (
            .O(N__37068),
            .I(N__36932));
    InMux I__9054 (
            .O(N__37067),
            .I(N__36929));
    InMux I__9053 (
            .O(N__37066),
            .I(N__36926));
    InMux I__9052 (
            .O(N__37065),
            .I(N__36923));
    InMux I__9051 (
            .O(N__37064),
            .I(N__36918));
    InMux I__9050 (
            .O(N__37063),
            .I(N__36918));
    LocalMux I__9049 (
            .O(N__37058),
            .I(N__36909));
    LocalMux I__9048 (
            .O(N__37053),
            .I(N__36909));
    Span4Mux_h I__9047 (
            .O(N__37050),
            .I(N__36909));
    LocalMux I__9046 (
            .O(N__37047),
            .I(N__36909));
    InMux I__9045 (
            .O(N__37046),
            .I(N__36904));
    InMux I__9044 (
            .O(N__37045),
            .I(N__36904));
    InMux I__9043 (
            .O(N__37044),
            .I(N__36901));
    InMux I__9042 (
            .O(N__37043),
            .I(N__36898));
    InMux I__9041 (
            .O(N__37042),
            .I(N__36894));
    LocalMux I__9040 (
            .O(N__37039),
            .I(N__36889));
    LocalMux I__9039 (
            .O(N__37034),
            .I(N__36889));
    LocalMux I__9038 (
            .O(N__37031),
            .I(N__36884));
    Span4Mux_v I__9037 (
            .O(N__37026),
            .I(N__36884));
    InMux I__9036 (
            .O(N__37023),
            .I(N__36881));
    LocalMux I__9035 (
            .O(N__37018),
            .I(N__36874));
    LocalMux I__9034 (
            .O(N__37011),
            .I(N__36874));
    LocalMux I__9033 (
            .O(N__37004),
            .I(N__36874));
    InMux I__9032 (
            .O(N__37003),
            .I(N__36867));
    InMux I__9031 (
            .O(N__37002),
            .I(N__36867));
    InMux I__9030 (
            .O(N__37001),
            .I(N__36867));
    LocalMux I__9029 (
            .O(N__36994),
            .I(N__36862));
    LocalMux I__9028 (
            .O(N__36989),
            .I(N__36862));
    InMux I__9027 (
            .O(N__36988),
            .I(N__36853));
    InMux I__9026 (
            .O(N__36987),
            .I(N__36853));
    InMux I__9025 (
            .O(N__36986),
            .I(N__36853));
    InMux I__9024 (
            .O(N__36985),
            .I(N__36853));
    InMux I__9023 (
            .O(N__36984),
            .I(N__36845));
    InMux I__9022 (
            .O(N__36983),
            .I(N__36845));
    InMux I__9021 (
            .O(N__36982),
            .I(N__36845));
    InMux I__9020 (
            .O(N__36981),
            .I(N__36842));
    CascadeMux I__9019 (
            .O(N__36980),
            .I(N__36838));
    InMux I__9018 (
            .O(N__36979),
            .I(N__36833));
    InMux I__9017 (
            .O(N__36978),
            .I(N__36833));
    LocalMux I__9016 (
            .O(N__36973),
            .I(N__36826));
    Span4Mux_h I__9015 (
            .O(N__36970),
            .I(N__36826));
    LocalMux I__9014 (
            .O(N__36959),
            .I(N__36826));
    InMux I__9013 (
            .O(N__36958),
            .I(N__36819));
    InMux I__9012 (
            .O(N__36957),
            .I(N__36819));
    InMux I__9011 (
            .O(N__36956),
            .I(N__36819));
    InMux I__9010 (
            .O(N__36955),
            .I(N__36810));
    InMux I__9009 (
            .O(N__36954),
            .I(N__36810));
    InMux I__9008 (
            .O(N__36953),
            .I(N__36810));
    InMux I__9007 (
            .O(N__36952),
            .I(N__36810));
    InMux I__9006 (
            .O(N__36951),
            .I(N__36805));
    InMux I__9005 (
            .O(N__36950),
            .I(N__36805));
    InMux I__9004 (
            .O(N__36949),
            .I(N__36798));
    InMux I__9003 (
            .O(N__36948),
            .I(N__36798));
    InMux I__9002 (
            .O(N__36947),
            .I(N__36798));
    InMux I__9001 (
            .O(N__36946),
            .I(N__36790));
    InMux I__9000 (
            .O(N__36945),
            .I(N__36790));
    LocalMux I__8999 (
            .O(N__36942),
            .I(N__36785));
    LocalMux I__8998 (
            .O(N__36937),
            .I(N__36785));
    CascadeMux I__8997 (
            .O(N__36936),
            .I(N__36781));
    CascadeMux I__8996 (
            .O(N__36935),
            .I(N__36777));
    LocalMux I__8995 (
            .O(N__36932),
            .I(N__36774));
    LocalMux I__8994 (
            .O(N__36929),
            .I(N__36771));
    LocalMux I__8993 (
            .O(N__36926),
            .I(N__36768));
    LocalMux I__8992 (
            .O(N__36923),
            .I(N__36759));
    LocalMux I__8991 (
            .O(N__36918),
            .I(N__36759));
    Span4Mux_v I__8990 (
            .O(N__36909),
            .I(N__36759));
    LocalMux I__8989 (
            .O(N__36904),
            .I(N__36759));
    LocalMux I__8988 (
            .O(N__36901),
            .I(N__36754));
    LocalMux I__8987 (
            .O(N__36898),
            .I(N__36754));
    InMux I__8986 (
            .O(N__36897),
            .I(N__36750));
    LocalMux I__8985 (
            .O(N__36894),
            .I(N__36733));
    Span4Mux_v I__8984 (
            .O(N__36889),
            .I(N__36733));
    Span4Mux_h I__8983 (
            .O(N__36884),
            .I(N__36733));
    LocalMux I__8982 (
            .O(N__36881),
            .I(N__36733));
    Span4Mux_h I__8981 (
            .O(N__36874),
            .I(N__36733));
    LocalMux I__8980 (
            .O(N__36867),
            .I(N__36733));
    Span4Mux_v I__8979 (
            .O(N__36862),
            .I(N__36728));
    LocalMux I__8978 (
            .O(N__36853),
            .I(N__36728));
    InMux I__8977 (
            .O(N__36852),
            .I(N__36724));
    LocalMux I__8976 (
            .O(N__36845),
            .I(N__36719));
    LocalMux I__8975 (
            .O(N__36842),
            .I(N__36719));
    InMux I__8974 (
            .O(N__36841),
            .I(N__36716));
    InMux I__8973 (
            .O(N__36838),
            .I(N__36713));
    LocalMux I__8972 (
            .O(N__36833),
            .I(N__36704));
    Sp12to4 I__8971 (
            .O(N__36826),
            .I(N__36704));
    LocalMux I__8970 (
            .O(N__36819),
            .I(N__36704));
    LocalMux I__8969 (
            .O(N__36810),
            .I(N__36704));
    LocalMux I__8968 (
            .O(N__36805),
            .I(N__36699));
    LocalMux I__8967 (
            .O(N__36798),
            .I(N__36699));
    InMux I__8966 (
            .O(N__36797),
            .I(N__36694));
    InMux I__8965 (
            .O(N__36796),
            .I(N__36689));
    InMux I__8964 (
            .O(N__36795),
            .I(N__36689));
    LocalMux I__8963 (
            .O(N__36790),
            .I(N__36686));
    Span4Mux_v I__8962 (
            .O(N__36785),
            .I(N__36683));
    InMux I__8961 (
            .O(N__36784),
            .I(N__36678));
    InMux I__8960 (
            .O(N__36781),
            .I(N__36678));
    InMux I__8959 (
            .O(N__36780),
            .I(N__36673));
    InMux I__8958 (
            .O(N__36777),
            .I(N__36673));
    Span4Mux_v I__8957 (
            .O(N__36774),
            .I(N__36662));
    Span4Mux_s3_v I__8956 (
            .O(N__36771),
            .I(N__36662));
    Span4Mux_s3_v I__8955 (
            .O(N__36768),
            .I(N__36662));
    Span4Mux_s3_v I__8954 (
            .O(N__36759),
            .I(N__36662));
    Span4Mux_v I__8953 (
            .O(N__36754),
            .I(N__36662));
    InMux I__8952 (
            .O(N__36753),
            .I(N__36659));
    LocalMux I__8951 (
            .O(N__36750),
            .I(N__36656));
    InMux I__8950 (
            .O(N__36749),
            .I(N__36647));
    InMux I__8949 (
            .O(N__36748),
            .I(N__36647));
    InMux I__8948 (
            .O(N__36747),
            .I(N__36647));
    InMux I__8947 (
            .O(N__36746),
            .I(N__36647));
    Span4Mux_h I__8946 (
            .O(N__36733),
            .I(N__36644));
    Span4Mux_h I__8945 (
            .O(N__36728),
            .I(N__36641));
    CascadeMux I__8944 (
            .O(N__36727),
            .I(N__36638));
    LocalMux I__8943 (
            .O(N__36724),
            .I(N__36635));
    Span4Mux_s3_h I__8942 (
            .O(N__36719),
            .I(N__36632));
    LocalMux I__8941 (
            .O(N__36716),
            .I(N__36627));
    LocalMux I__8940 (
            .O(N__36713),
            .I(N__36627));
    Span12Mux_s3_v I__8939 (
            .O(N__36704),
            .I(N__36622));
    Span12Mux_s10_v I__8938 (
            .O(N__36699),
            .I(N__36622));
    InMux I__8937 (
            .O(N__36698),
            .I(N__36617));
    InMux I__8936 (
            .O(N__36697),
            .I(N__36617));
    LocalMux I__8935 (
            .O(N__36694),
            .I(N__36596));
    LocalMux I__8934 (
            .O(N__36689),
            .I(N__36596));
    Span12Mux_s3_v I__8933 (
            .O(N__36686),
            .I(N__36596));
    Sp12to4 I__8932 (
            .O(N__36683),
            .I(N__36596));
    LocalMux I__8931 (
            .O(N__36678),
            .I(N__36596));
    LocalMux I__8930 (
            .O(N__36673),
            .I(N__36596));
    Sp12to4 I__8929 (
            .O(N__36662),
            .I(N__36596));
    LocalMux I__8928 (
            .O(N__36659),
            .I(N__36596));
    Span12Mux_s2_h I__8927 (
            .O(N__36656),
            .I(N__36596));
    LocalMux I__8926 (
            .O(N__36647),
            .I(N__36596));
    Span4Mux_v I__8925 (
            .O(N__36644),
            .I(N__36591));
    Span4Mux_h I__8924 (
            .O(N__36641),
            .I(N__36591));
    InMux I__8923 (
            .O(N__36638),
            .I(N__36588));
    Odrv4 I__8922 (
            .O(N__36635),
            .I(\tok.T_5 ));
    Odrv4 I__8921 (
            .O(N__36632),
            .I(\tok.T_5 ));
    Odrv4 I__8920 (
            .O(N__36627),
            .I(\tok.T_5 ));
    Odrv12 I__8919 (
            .O(N__36622),
            .I(\tok.T_5 ));
    LocalMux I__8918 (
            .O(N__36617),
            .I(\tok.T_5 ));
    Odrv12 I__8917 (
            .O(N__36596),
            .I(\tok.T_5 ));
    Odrv4 I__8916 (
            .O(N__36591),
            .I(\tok.T_5 ));
    LocalMux I__8915 (
            .O(N__36588),
            .I(\tok.T_5 ));
    InMux I__8914 (
            .O(N__36571),
            .I(N__36568));
    LocalMux I__8913 (
            .O(N__36568),
            .I(N__36565));
    Span4Mux_h I__8912 (
            .O(N__36565),
            .I(N__36562));
    Odrv4 I__8911 (
            .O(N__36562),
            .I(\tok.n317 ));
    CascadeMux I__8910 (
            .O(N__36559),
            .I(\tok.n317_cascade_ ));
    CascadeMux I__8909 (
            .O(N__36556),
            .I(N__36550));
    InMux I__8908 (
            .O(N__36555),
            .I(N__36545));
    InMux I__8907 (
            .O(N__36554),
            .I(N__36542));
    InMux I__8906 (
            .O(N__36553),
            .I(N__36536));
    InMux I__8905 (
            .O(N__36550),
            .I(N__36536));
    InMux I__8904 (
            .O(N__36549),
            .I(N__36529));
    InMux I__8903 (
            .O(N__36548),
            .I(N__36525));
    LocalMux I__8902 (
            .O(N__36545),
            .I(N__36520));
    LocalMux I__8901 (
            .O(N__36542),
            .I(N__36520));
    CascadeMux I__8900 (
            .O(N__36541),
            .I(N__36517));
    LocalMux I__8899 (
            .O(N__36536),
            .I(N__36514));
    InMux I__8898 (
            .O(N__36535),
            .I(N__36510));
    CascadeMux I__8897 (
            .O(N__36534),
            .I(N__36506));
    InMux I__8896 (
            .O(N__36533),
            .I(N__36503));
    InMux I__8895 (
            .O(N__36532),
            .I(N__36500));
    LocalMux I__8894 (
            .O(N__36529),
            .I(N__36497));
    InMux I__8893 (
            .O(N__36528),
            .I(N__36494));
    LocalMux I__8892 (
            .O(N__36525),
            .I(N__36489));
    Span4Mux_h I__8891 (
            .O(N__36520),
            .I(N__36489));
    InMux I__8890 (
            .O(N__36517),
            .I(N__36486));
    Span4Mux_h I__8889 (
            .O(N__36514),
            .I(N__36483));
    InMux I__8888 (
            .O(N__36513),
            .I(N__36480));
    LocalMux I__8887 (
            .O(N__36510),
            .I(N__36476));
    InMux I__8886 (
            .O(N__36509),
            .I(N__36473));
    InMux I__8885 (
            .O(N__36506),
            .I(N__36470));
    LocalMux I__8884 (
            .O(N__36503),
            .I(N__36467));
    LocalMux I__8883 (
            .O(N__36500),
            .I(N__36464));
    Span4Mux_v I__8882 (
            .O(N__36497),
            .I(N__36461));
    LocalMux I__8881 (
            .O(N__36494),
            .I(N__36458));
    Span4Mux_s2_v I__8880 (
            .O(N__36489),
            .I(N__36446));
    LocalMux I__8879 (
            .O(N__36486),
            .I(N__36446));
    Span4Mux_s2_v I__8878 (
            .O(N__36483),
            .I(N__36446));
    LocalMux I__8877 (
            .O(N__36480),
            .I(N__36443));
    InMux I__8876 (
            .O(N__36479),
            .I(N__36440));
    Span4Mux_v I__8875 (
            .O(N__36476),
            .I(N__36435));
    LocalMux I__8874 (
            .O(N__36473),
            .I(N__36435));
    LocalMux I__8873 (
            .O(N__36470),
            .I(N__36430));
    Span4Mux_h I__8872 (
            .O(N__36467),
            .I(N__36430));
    Span4Mux_v I__8871 (
            .O(N__36464),
            .I(N__36425));
    Span4Mux_h I__8870 (
            .O(N__36461),
            .I(N__36425));
    Span4Mux_h I__8869 (
            .O(N__36458),
            .I(N__36422));
    InMux I__8868 (
            .O(N__36457),
            .I(N__36413));
    InMux I__8867 (
            .O(N__36456),
            .I(N__36413));
    InMux I__8866 (
            .O(N__36455),
            .I(N__36413));
    InMux I__8865 (
            .O(N__36454),
            .I(N__36413));
    InMux I__8864 (
            .O(N__36453),
            .I(N__36410));
    Span4Mux_v I__8863 (
            .O(N__36446),
            .I(N__36407));
    Odrv4 I__8862 (
            .O(N__36443),
            .I(\tok.A_low_3 ));
    LocalMux I__8861 (
            .O(N__36440),
            .I(\tok.A_low_3 ));
    Odrv4 I__8860 (
            .O(N__36435),
            .I(\tok.A_low_3 ));
    Odrv4 I__8859 (
            .O(N__36430),
            .I(\tok.A_low_3 ));
    Odrv4 I__8858 (
            .O(N__36425),
            .I(\tok.A_low_3 ));
    Odrv4 I__8857 (
            .O(N__36422),
            .I(\tok.A_low_3 ));
    LocalMux I__8856 (
            .O(N__36413),
            .I(\tok.A_low_3 ));
    LocalMux I__8855 (
            .O(N__36410),
            .I(\tok.A_low_3 ));
    Odrv4 I__8854 (
            .O(N__36407),
            .I(\tok.A_low_3 ));
    InMux I__8853 (
            .O(N__36388),
            .I(N__36385));
    LocalMux I__8852 (
            .O(N__36385),
            .I(N__36382));
    Span4Mux_v I__8851 (
            .O(N__36382),
            .I(N__36379));
    Odrv4 I__8850 (
            .O(N__36379),
            .I(\tok.n168 ));
    CascadeMux I__8849 (
            .O(N__36376),
            .I(N__36371));
    InMux I__8848 (
            .O(N__36375),
            .I(N__36368));
    InMux I__8847 (
            .O(N__36374),
            .I(N__36365));
    InMux I__8846 (
            .O(N__36371),
            .I(N__36361));
    LocalMux I__8845 (
            .O(N__36368),
            .I(N__36358));
    LocalMux I__8844 (
            .O(N__36365),
            .I(N__36355));
    InMux I__8843 (
            .O(N__36364),
            .I(N__36352));
    LocalMux I__8842 (
            .O(N__36361),
            .I(N__36349));
    Span4Mux_h I__8841 (
            .O(N__36358),
            .I(N__36342));
    Span4Mux_v I__8840 (
            .O(N__36355),
            .I(N__36342));
    LocalMux I__8839 (
            .O(N__36352),
            .I(N__36342));
    Span4Mux_h I__8838 (
            .O(N__36349),
            .I(N__36338));
    Span4Mux_h I__8837 (
            .O(N__36342),
            .I(N__36335));
    InMux I__8836 (
            .O(N__36341),
            .I(N__36332));
    Odrv4 I__8835 (
            .O(N__36338),
            .I(\tok.n5_adj_682 ));
    Odrv4 I__8834 (
            .O(N__36335),
            .I(\tok.n5_adj_682 ));
    LocalMux I__8833 (
            .O(N__36332),
            .I(\tok.n5_adj_682 ));
    CascadeMux I__8832 (
            .O(N__36325),
            .I(N__36312));
    InMux I__8831 (
            .O(N__36324),
            .I(N__36307));
    CascadeMux I__8830 (
            .O(N__36323),
            .I(N__36288));
    CascadeMux I__8829 (
            .O(N__36322),
            .I(N__36276));
    CascadeMux I__8828 (
            .O(N__36321),
            .I(N__36273));
    CascadeMux I__8827 (
            .O(N__36320),
            .I(N__36270));
    InMux I__8826 (
            .O(N__36319),
            .I(N__36262));
    InMux I__8825 (
            .O(N__36318),
            .I(N__36262));
    InMux I__8824 (
            .O(N__36317),
            .I(N__36262));
    InMux I__8823 (
            .O(N__36316),
            .I(N__36246));
    InMux I__8822 (
            .O(N__36315),
            .I(N__36239));
    InMux I__8821 (
            .O(N__36312),
            .I(N__36239));
    InMux I__8820 (
            .O(N__36311),
            .I(N__36239));
    CascadeMux I__8819 (
            .O(N__36310),
            .I(N__36236));
    LocalMux I__8818 (
            .O(N__36307),
            .I(N__36224));
    InMux I__8817 (
            .O(N__36306),
            .I(N__36221));
    CascadeMux I__8816 (
            .O(N__36305),
            .I(N__36216));
    CascadeMux I__8815 (
            .O(N__36304),
            .I(N__36210));
    CascadeMux I__8814 (
            .O(N__36303),
            .I(N__36207));
    InMux I__8813 (
            .O(N__36302),
            .I(N__36199));
    InMux I__8812 (
            .O(N__36301),
            .I(N__36199));
    InMux I__8811 (
            .O(N__36300),
            .I(N__36199));
    InMux I__8810 (
            .O(N__36299),
            .I(N__36196));
    InMux I__8809 (
            .O(N__36298),
            .I(N__36191));
    InMux I__8808 (
            .O(N__36297),
            .I(N__36191));
    InMux I__8807 (
            .O(N__36296),
            .I(N__36186));
    InMux I__8806 (
            .O(N__36295),
            .I(N__36186));
    CascadeMux I__8805 (
            .O(N__36294),
            .I(N__36180));
    InMux I__8804 (
            .O(N__36293),
            .I(N__36174));
    InMux I__8803 (
            .O(N__36292),
            .I(N__36169));
    InMux I__8802 (
            .O(N__36291),
            .I(N__36169));
    InMux I__8801 (
            .O(N__36288),
            .I(N__36166));
    InMux I__8800 (
            .O(N__36287),
            .I(N__36157));
    InMux I__8799 (
            .O(N__36286),
            .I(N__36157));
    InMux I__8798 (
            .O(N__36285),
            .I(N__36157));
    InMux I__8797 (
            .O(N__36284),
            .I(N__36157));
    CascadeMux I__8796 (
            .O(N__36283),
            .I(N__36139));
    InMux I__8795 (
            .O(N__36282),
            .I(N__36135));
    InMux I__8794 (
            .O(N__36281),
            .I(N__36132));
    InMux I__8793 (
            .O(N__36280),
            .I(N__36121));
    InMux I__8792 (
            .O(N__36279),
            .I(N__36121));
    InMux I__8791 (
            .O(N__36276),
            .I(N__36121));
    InMux I__8790 (
            .O(N__36273),
            .I(N__36121));
    InMux I__8789 (
            .O(N__36270),
            .I(N__36121));
    InMux I__8788 (
            .O(N__36269),
            .I(N__36118));
    LocalMux I__8787 (
            .O(N__36262),
            .I(N__36115));
    InMux I__8786 (
            .O(N__36261),
            .I(N__36108));
    InMux I__8785 (
            .O(N__36260),
            .I(N__36108));
    InMux I__8784 (
            .O(N__36259),
            .I(N__36108));
    InMux I__8783 (
            .O(N__36258),
            .I(N__36103));
    InMux I__8782 (
            .O(N__36257),
            .I(N__36103));
    CascadeMux I__8781 (
            .O(N__36256),
            .I(N__36099));
    InMux I__8780 (
            .O(N__36255),
            .I(N__36092));
    InMux I__8779 (
            .O(N__36254),
            .I(N__36092));
    InMux I__8778 (
            .O(N__36253),
            .I(N__36089));
    InMux I__8777 (
            .O(N__36252),
            .I(N__36086));
    InMux I__8776 (
            .O(N__36251),
            .I(N__36079));
    InMux I__8775 (
            .O(N__36250),
            .I(N__36079));
    InMux I__8774 (
            .O(N__36249),
            .I(N__36079));
    LocalMux I__8773 (
            .O(N__36246),
            .I(N__36074));
    LocalMux I__8772 (
            .O(N__36239),
            .I(N__36074));
    InMux I__8771 (
            .O(N__36236),
            .I(N__36065));
    InMux I__8770 (
            .O(N__36235),
            .I(N__36065));
    InMux I__8769 (
            .O(N__36234),
            .I(N__36065));
    InMux I__8768 (
            .O(N__36233),
            .I(N__36065));
    InMux I__8767 (
            .O(N__36232),
            .I(N__36062));
    CascadeMux I__8766 (
            .O(N__36231),
            .I(N__36059));
    InMux I__8765 (
            .O(N__36230),
            .I(N__36056));
    InMux I__8764 (
            .O(N__36229),
            .I(N__36053));
    CascadeMux I__8763 (
            .O(N__36228),
            .I(N__36045));
    InMux I__8762 (
            .O(N__36227),
            .I(N__36041));
    Span4Mux_h I__8761 (
            .O(N__36224),
            .I(N__36036));
    LocalMux I__8760 (
            .O(N__36221),
            .I(N__36036));
    InMux I__8759 (
            .O(N__36220),
            .I(N__36033));
    InMux I__8758 (
            .O(N__36219),
            .I(N__36024));
    InMux I__8757 (
            .O(N__36216),
            .I(N__36024));
    InMux I__8756 (
            .O(N__36215),
            .I(N__36019));
    InMux I__8755 (
            .O(N__36214),
            .I(N__36019));
    CascadeMux I__8754 (
            .O(N__36213),
            .I(N__36011));
    InMux I__8753 (
            .O(N__36210),
            .I(N__36002));
    InMux I__8752 (
            .O(N__36207),
            .I(N__36002));
    InMux I__8751 (
            .O(N__36206),
            .I(N__36002));
    LocalMux I__8750 (
            .O(N__36199),
            .I(N__35999));
    LocalMux I__8749 (
            .O(N__36196),
            .I(N__35992));
    LocalMux I__8748 (
            .O(N__36191),
            .I(N__35992));
    LocalMux I__8747 (
            .O(N__36186),
            .I(N__35992));
    InMux I__8746 (
            .O(N__36185),
            .I(N__35989));
    InMux I__8745 (
            .O(N__36184),
            .I(N__35986));
    InMux I__8744 (
            .O(N__36183),
            .I(N__35983));
    InMux I__8743 (
            .O(N__36180),
            .I(N__35976));
    InMux I__8742 (
            .O(N__36179),
            .I(N__35976));
    InMux I__8741 (
            .O(N__36178),
            .I(N__35976));
    InMux I__8740 (
            .O(N__36177),
            .I(N__35973));
    LocalMux I__8739 (
            .O(N__36174),
            .I(N__35969));
    LocalMux I__8738 (
            .O(N__36169),
            .I(N__35962));
    LocalMux I__8737 (
            .O(N__36166),
            .I(N__35962));
    LocalMux I__8736 (
            .O(N__36157),
            .I(N__35962));
    InMux I__8735 (
            .O(N__36156),
            .I(N__35953));
    InMux I__8734 (
            .O(N__36155),
            .I(N__35953));
    InMux I__8733 (
            .O(N__36154),
            .I(N__35953));
    InMux I__8732 (
            .O(N__36153),
            .I(N__35953));
    InMux I__8731 (
            .O(N__36152),
            .I(N__35944));
    InMux I__8730 (
            .O(N__36151),
            .I(N__35944));
    InMux I__8729 (
            .O(N__36150),
            .I(N__35944));
    InMux I__8728 (
            .O(N__36149),
            .I(N__35939));
    InMux I__8727 (
            .O(N__36148),
            .I(N__35939));
    InMux I__8726 (
            .O(N__36147),
            .I(N__35936));
    InMux I__8725 (
            .O(N__36146),
            .I(N__35927));
    InMux I__8724 (
            .O(N__36145),
            .I(N__35927));
    InMux I__8723 (
            .O(N__36144),
            .I(N__35927));
    InMux I__8722 (
            .O(N__36143),
            .I(N__35927));
    InMux I__8721 (
            .O(N__36142),
            .I(N__35922));
    InMux I__8720 (
            .O(N__36139),
            .I(N__35922));
    CascadeMux I__8719 (
            .O(N__36138),
            .I(N__35919));
    LocalMux I__8718 (
            .O(N__36135),
            .I(N__35915));
    LocalMux I__8717 (
            .O(N__36132),
            .I(N__35910));
    LocalMux I__8716 (
            .O(N__36121),
            .I(N__35910));
    LocalMux I__8715 (
            .O(N__36118),
            .I(N__35901));
    Span4Mux_v I__8714 (
            .O(N__36115),
            .I(N__35901));
    LocalMux I__8713 (
            .O(N__36108),
            .I(N__35901));
    LocalMux I__8712 (
            .O(N__36103),
            .I(N__35901));
    InMux I__8711 (
            .O(N__36102),
            .I(N__35896));
    InMux I__8710 (
            .O(N__36099),
            .I(N__35896));
    InMux I__8709 (
            .O(N__36098),
            .I(N__35891));
    InMux I__8708 (
            .O(N__36097),
            .I(N__35891));
    LocalMux I__8707 (
            .O(N__36092),
            .I(N__35882));
    LocalMux I__8706 (
            .O(N__36089),
            .I(N__35882));
    LocalMux I__8705 (
            .O(N__36086),
            .I(N__35882));
    LocalMux I__8704 (
            .O(N__36079),
            .I(N__35882));
    Span4Mux_s2_v I__8703 (
            .O(N__36074),
            .I(N__35875));
    LocalMux I__8702 (
            .O(N__36065),
            .I(N__35875));
    LocalMux I__8701 (
            .O(N__36062),
            .I(N__35875));
    InMux I__8700 (
            .O(N__36059),
            .I(N__35871));
    LocalMux I__8699 (
            .O(N__36056),
            .I(N__35868));
    LocalMux I__8698 (
            .O(N__36053),
            .I(N__35865));
    InMux I__8697 (
            .O(N__36052),
            .I(N__35858));
    InMux I__8696 (
            .O(N__36051),
            .I(N__35858));
    InMux I__8695 (
            .O(N__36050),
            .I(N__35858));
    InMux I__8694 (
            .O(N__36049),
            .I(N__35855));
    InMux I__8693 (
            .O(N__36048),
            .I(N__35852));
    InMux I__8692 (
            .O(N__36045),
            .I(N__35849));
    InMux I__8691 (
            .O(N__36044),
            .I(N__35846));
    LocalMux I__8690 (
            .O(N__36041),
            .I(N__35839));
    Span4Mux_h I__8689 (
            .O(N__36036),
            .I(N__35839));
    LocalMux I__8688 (
            .O(N__36033),
            .I(N__35839));
    InMux I__8687 (
            .O(N__36032),
            .I(N__35836));
    CascadeMux I__8686 (
            .O(N__36031),
            .I(N__35832));
    InMux I__8685 (
            .O(N__36030),
            .I(N__35825));
    InMux I__8684 (
            .O(N__36029),
            .I(N__35822));
    LocalMux I__8683 (
            .O(N__36024),
            .I(N__35817));
    LocalMux I__8682 (
            .O(N__36019),
            .I(N__35817));
    InMux I__8681 (
            .O(N__36018),
            .I(N__35804));
    InMux I__8680 (
            .O(N__36017),
            .I(N__35804));
    InMux I__8679 (
            .O(N__36016),
            .I(N__35804));
    InMux I__8678 (
            .O(N__36015),
            .I(N__35804));
    InMux I__8677 (
            .O(N__36014),
            .I(N__35804));
    InMux I__8676 (
            .O(N__36011),
            .I(N__35804));
    InMux I__8675 (
            .O(N__36010),
            .I(N__35799));
    InMux I__8674 (
            .O(N__36009),
            .I(N__35799));
    LocalMux I__8673 (
            .O(N__36002),
            .I(N__35792));
    Span4Mux_s3_h I__8672 (
            .O(N__35999),
            .I(N__35792));
    Span4Mux_v I__8671 (
            .O(N__35992),
            .I(N__35792));
    LocalMux I__8670 (
            .O(N__35989),
            .I(N__35783));
    LocalMux I__8669 (
            .O(N__35986),
            .I(N__35783));
    LocalMux I__8668 (
            .O(N__35983),
            .I(N__35783));
    LocalMux I__8667 (
            .O(N__35976),
            .I(N__35783));
    LocalMux I__8666 (
            .O(N__35973),
            .I(N__35780));
    InMux I__8665 (
            .O(N__35972),
            .I(N__35775));
    Span4Mux_v I__8664 (
            .O(N__35969),
            .I(N__35768));
    Span4Mux_v I__8663 (
            .O(N__35962),
            .I(N__35768));
    LocalMux I__8662 (
            .O(N__35953),
            .I(N__35768));
    InMux I__8661 (
            .O(N__35952),
            .I(N__35758));
    InMux I__8660 (
            .O(N__35951),
            .I(N__35758));
    LocalMux I__8659 (
            .O(N__35944),
            .I(N__35749));
    LocalMux I__8658 (
            .O(N__35939),
            .I(N__35749));
    LocalMux I__8657 (
            .O(N__35936),
            .I(N__35749));
    LocalMux I__8656 (
            .O(N__35927),
            .I(N__35749));
    LocalMux I__8655 (
            .O(N__35922),
            .I(N__35746));
    InMux I__8654 (
            .O(N__35919),
            .I(N__35741));
    InMux I__8653 (
            .O(N__35918),
            .I(N__35741));
    Span4Mux_s3_v I__8652 (
            .O(N__35915),
            .I(N__35734));
    Span4Mux_s3_v I__8651 (
            .O(N__35910),
            .I(N__35734));
    Span4Mux_v I__8650 (
            .O(N__35901),
            .I(N__35734));
    LocalMux I__8649 (
            .O(N__35896),
            .I(N__35725));
    LocalMux I__8648 (
            .O(N__35891),
            .I(N__35725));
    Span4Mux_v I__8647 (
            .O(N__35882),
            .I(N__35725));
    Span4Mux_v I__8646 (
            .O(N__35875),
            .I(N__35725));
    CascadeMux I__8645 (
            .O(N__35874),
            .I(N__35718));
    LocalMux I__8644 (
            .O(N__35871),
            .I(N__35712));
    Span4Mux_v I__8643 (
            .O(N__35868),
            .I(N__35707));
    Span4Mux_s3_v I__8642 (
            .O(N__35865),
            .I(N__35707));
    LocalMux I__8641 (
            .O(N__35858),
            .I(N__35704));
    LocalMux I__8640 (
            .O(N__35855),
            .I(N__35701));
    LocalMux I__8639 (
            .O(N__35852),
            .I(N__35692));
    LocalMux I__8638 (
            .O(N__35849),
            .I(N__35692));
    LocalMux I__8637 (
            .O(N__35846),
            .I(N__35692));
    Span4Mux_v I__8636 (
            .O(N__35839),
            .I(N__35692));
    LocalMux I__8635 (
            .O(N__35836),
            .I(N__35689));
    InMux I__8634 (
            .O(N__35835),
            .I(N__35676));
    InMux I__8633 (
            .O(N__35832),
            .I(N__35676));
    InMux I__8632 (
            .O(N__35831),
            .I(N__35676));
    InMux I__8631 (
            .O(N__35830),
            .I(N__35676));
    InMux I__8630 (
            .O(N__35829),
            .I(N__35676));
    InMux I__8629 (
            .O(N__35828),
            .I(N__35676));
    LocalMux I__8628 (
            .O(N__35825),
            .I(N__35671));
    LocalMux I__8627 (
            .O(N__35822),
            .I(N__35671));
    Span4Mux_h I__8626 (
            .O(N__35817),
            .I(N__35668));
    LocalMux I__8625 (
            .O(N__35804),
            .I(N__35659));
    LocalMux I__8624 (
            .O(N__35799),
            .I(N__35659));
    Span4Mux_h I__8623 (
            .O(N__35792),
            .I(N__35659));
    Span4Mux_v I__8622 (
            .O(N__35783),
            .I(N__35659));
    Span4Mux_s3_v I__8621 (
            .O(N__35780),
            .I(N__35656));
    InMux I__8620 (
            .O(N__35779),
            .I(N__35653));
    InMux I__8619 (
            .O(N__35778),
            .I(N__35650));
    LocalMux I__8618 (
            .O(N__35775),
            .I(N__35647));
    Span4Mux_s3_v I__8617 (
            .O(N__35768),
            .I(N__35644));
    InMux I__8616 (
            .O(N__35767),
            .I(N__35641));
    InMux I__8615 (
            .O(N__35766),
            .I(N__35632));
    InMux I__8614 (
            .O(N__35765),
            .I(N__35632));
    InMux I__8613 (
            .O(N__35764),
            .I(N__35632));
    InMux I__8612 (
            .O(N__35763),
            .I(N__35632));
    LocalMux I__8611 (
            .O(N__35758),
            .I(N__35629));
    Span4Mux_s3_v I__8610 (
            .O(N__35749),
            .I(N__35618));
    Span4Mux_s3_v I__8609 (
            .O(N__35746),
            .I(N__35618));
    LocalMux I__8608 (
            .O(N__35741),
            .I(N__35618));
    Span4Mux_h I__8607 (
            .O(N__35734),
            .I(N__35618));
    Span4Mux_v I__8606 (
            .O(N__35725),
            .I(N__35618));
    InMux I__8605 (
            .O(N__35724),
            .I(N__35613));
    InMux I__8604 (
            .O(N__35723),
            .I(N__35613));
    InMux I__8603 (
            .O(N__35722),
            .I(N__35607));
    InMux I__8602 (
            .O(N__35721),
            .I(N__35598));
    InMux I__8601 (
            .O(N__35718),
            .I(N__35598));
    InMux I__8600 (
            .O(N__35717),
            .I(N__35598));
    InMux I__8599 (
            .O(N__35716),
            .I(N__35598));
    InMux I__8598 (
            .O(N__35715),
            .I(N__35595));
    Span12Mux_s10_v I__8597 (
            .O(N__35712),
            .I(N__35592));
    Span4Mux_h I__8596 (
            .O(N__35707),
            .I(N__35573));
    Span4Mux_s3_v I__8595 (
            .O(N__35704),
            .I(N__35573));
    Span4Mux_v I__8594 (
            .O(N__35701),
            .I(N__35573));
    Span4Mux_v I__8593 (
            .O(N__35692),
            .I(N__35573));
    Span4Mux_s3_v I__8592 (
            .O(N__35689),
            .I(N__35573));
    LocalMux I__8591 (
            .O(N__35676),
            .I(N__35573));
    Span4Mux_s3_v I__8590 (
            .O(N__35671),
            .I(N__35573));
    Span4Mux_v I__8589 (
            .O(N__35668),
            .I(N__35573));
    Span4Mux_v I__8588 (
            .O(N__35659),
            .I(N__35573));
    Sp12to4 I__8587 (
            .O(N__35656),
            .I(N__35552));
    LocalMux I__8586 (
            .O(N__35653),
            .I(N__35552));
    LocalMux I__8585 (
            .O(N__35650),
            .I(N__35552));
    Span12Mux_s10_v I__8584 (
            .O(N__35647),
            .I(N__35552));
    Sp12to4 I__8583 (
            .O(N__35644),
            .I(N__35552));
    LocalMux I__8582 (
            .O(N__35641),
            .I(N__35552));
    LocalMux I__8581 (
            .O(N__35632),
            .I(N__35552));
    Span12Mux_s1_h I__8580 (
            .O(N__35629),
            .I(N__35552));
    Sp12to4 I__8579 (
            .O(N__35618),
            .I(N__35552));
    LocalMux I__8578 (
            .O(N__35613),
            .I(N__35552));
    InMux I__8577 (
            .O(N__35612),
            .I(N__35549));
    InMux I__8576 (
            .O(N__35611),
            .I(N__35544));
    InMux I__8575 (
            .O(N__35610),
            .I(N__35544));
    LocalMux I__8574 (
            .O(N__35607),
            .I(\tok.T_4 ));
    LocalMux I__8573 (
            .O(N__35598),
            .I(\tok.T_4 ));
    LocalMux I__8572 (
            .O(N__35595),
            .I(\tok.T_4 ));
    Odrv12 I__8571 (
            .O(N__35592),
            .I(\tok.T_4 ));
    Odrv4 I__8570 (
            .O(N__35573),
            .I(\tok.T_4 ));
    Odrv12 I__8569 (
            .O(N__35552),
            .I(\tok.T_4 ));
    LocalMux I__8568 (
            .O(N__35549),
            .I(\tok.T_4 ));
    LocalMux I__8567 (
            .O(N__35544),
            .I(\tok.T_4 ));
    CascadeMux I__8566 (
            .O(N__35527),
            .I(\tok.n6478_cascade_ ));
    CascadeMux I__8565 (
            .O(N__35524),
            .I(N__35511));
    CascadeMux I__8564 (
            .O(N__35523),
            .I(N__35497));
    InMux I__8563 (
            .O(N__35522),
            .I(N__35475));
    InMux I__8562 (
            .O(N__35521),
            .I(N__35469));
    InMux I__8561 (
            .O(N__35520),
            .I(N__35469));
    InMux I__8560 (
            .O(N__35519),
            .I(N__35460));
    InMux I__8559 (
            .O(N__35518),
            .I(N__35460));
    InMux I__8558 (
            .O(N__35517),
            .I(N__35452));
    InMux I__8557 (
            .O(N__35516),
            .I(N__35447));
    InMux I__8556 (
            .O(N__35515),
            .I(N__35447));
    InMux I__8555 (
            .O(N__35514),
            .I(N__35435));
    InMux I__8554 (
            .O(N__35511),
            .I(N__35435));
    InMux I__8553 (
            .O(N__35510),
            .I(N__35435));
    InMux I__8552 (
            .O(N__35509),
            .I(N__35432));
    InMux I__8551 (
            .O(N__35508),
            .I(N__35427));
    InMux I__8550 (
            .O(N__35507),
            .I(N__35427));
    InMux I__8549 (
            .O(N__35506),
            .I(N__35424));
    CascadeMux I__8548 (
            .O(N__35505),
            .I(N__35420));
    InMux I__8547 (
            .O(N__35504),
            .I(N__35416));
    CascadeMux I__8546 (
            .O(N__35503),
            .I(N__35412));
    InMux I__8545 (
            .O(N__35502),
            .I(N__35409));
    InMux I__8544 (
            .O(N__35501),
            .I(N__35406));
    InMux I__8543 (
            .O(N__35500),
            .I(N__35403));
    InMux I__8542 (
            .O(N__35497),
            .I(N__35398));
    InMux I__8541 (
            .O(N__35496),
            .I(N__35398));
    CascadeMux I__8540 (
            .O(N__35495),
            .I(N__35391));
    InMux I__8539 (
            .O(N__35494),
            .I(N__35367));
    InMux I__8538 (
            .O(N__35493),
            .I(N__35358));
    InMux I__8537 (
            .O(N__35492),
            .I(N__35358));
    InMux I__8536 (
            .O(N__35491),
            .I(N__35358));
    InMux I__8535 (
            .O(N__35490),
            .I(N__35358));
    InMux I__8534 (
            .O(N__35489),
            .I(N__35353));
    InMux I__8533 (
            .O(N__35488),
            .I(N__35350));
    InMux I__8532 (
            .O(N__35487),
            .I(N__35347));
    InMux I__8531 (
            .O(N__35486),
            .I(N__35342));
    InMux I__8530 (
            .O(N__35485),
            .I(N__35342));
    InMux I__8529 (
            .O(N__35484),
            .I(N__35337));
    InMux I__8528 (
            .O(N__35483),
            .I(N__35337));
    InMux I__8527 (
            .O(N__35482),
            .I(N__35332));
    InMux I__8526 (
            .O(N__35481),
            .I(N__35332));
    InMux I__8525 (
            .O(N__35480),
            .I(N__35326));
    InMux I__8524 (
            .O(N__35479),
            .I(N__35321));
    InMux I__8523 (
            .O(N__35478),
            .I(N__35321));
    LocalMux I__8522 (
            .O(N__35475),
            .I(N__35318));
    InMux I__8521 (
            .O(N__35474),
            .I(N__35315));
    LocalMux I__8520 (
            .O(N__35469),
            .I(N__35312));
    InMux I__8519 (
            .O(N__35468),
            .I(N__35305));
    InMux I__8518 (
            .O(N__35467),
            .I(N__35305));
    InMux I__8517 (
            .O(N__35466),
            .I(N__35305));
    InMux I__8516 (
            .O(N__35465),
            .I(N__35302));
    LocalMux I__8515 (
            .O(N__35460),
            .I(N__35297));
    InMux I__8514 (
            .O(N__35459),
            .I(N__35288));
    InMux I__8513 (
            .O(N__35458),
            .I(N__35288));
    InMux I__8512 (
            .O(N__35457),
            .I(N__35288));
    InMux I__8511 (
            .O(N__35456),
            .I(N__35288));
    InMux I__8510 (
            .O(N__35455),
            .I(N__35285));
    LocalMux I__8509 (
            .O(N__35452),
            .I(N__35280));
    LocalMux I__8508 (
            .O(N__35447),
            .I(N__35280));
    InMux I__8507 (
            .O(N__35446),
            .I(N__35273));
    InMux I__8506 (
            .O(N__35445),
            .I(N__35273));
    CascadeMux I__8505 (
            .O(N__35444),
            .I(N__35269));
    InMux I__8504 (
            .O(N__35443),
            .I(N__35261));
    InMux I__8503 (
            .O(N__35442),
            .I(N__35257));
    LocalMux I__8502 (
            .O(N__35435),
            .I(N__35254));
    LocalMux I__8501 (
            .O(N__35432),
            .I(N__35247));
    LocalMux I__8500 (
            .O(N__35427),
            .I(N__35247));
    LocalMux I__8499 (
            .O(N__35424),
            .I(N__35247));
    InMux I__8498 (
            .O(N__35423),
            .I(N__35242));
    InMux I__8497 (
            .O(N__35420),
            .I(N__35242));
    InMux I__8496 (
            .O(N__35419),
            .I(N__35239));
    LocalMux I__8495 (
            .O(N__35416),
            .I(N__35234));
    InMux I__8494 (
            .O(N__35415),
            .I(N__35229));
    InMux I__8493 (
            .O(N__35412),
            .I(N__35229));
    LocalMux I__8492 (
            .O(N__35409),
            .I(N__35222));
    LocalMux I__8491 (
            .O(N__35406),
            .I(N__35222));
    LocalMux I__8490 (
            .O(N__35403),
            .I(N__35222));
    LocalMux I__8489 (
            .O(N__35398),
            .I(N__35219));
    InMux I__8488 (
            .O(N__35397),
            .I(N__35214));
    InMux I__8487 (
            .O(N__35396),
            .I(N__35214));
    InMux I__8486 (
            .O(N__35395),
            .I(N__35207));
    InMux I__8485 (
            .O(N__35394),
            .I(N__35207));
    InMux I__8484 (
            .O(N__35391),
            .I(N__35207));
    InMux I__8483 (
            .O(N__35390),
            .I(N__35203));
    InMux I__8482 (
            .O(N__35389),
            .I(N__35200));
    InMux I__8481 (
            .O(N__35388),
            .I(N__35187));
    InMux I__8480 (
            .O(N__35387),
            .I(N__35187));
    InMux I__8479 (
            .O(N__35386),
            .I(N__35187));
    InMux I__8478 (
            .O(N__35385),
            .I(N__35187));
    InMux I__8477 (
            .O(N__35384),
            .I(N__35187));
    InMux I__8476 (
            .O(N__35383),
            .I(N__35180));
    InMux I__8475 (
            .O(N__35382),
            .I(N__35180));
    InMux I__8474 (
            .O(N__35381),
            .I(N__35180));
    InMux I__8473 (
            .O(N__35380),
            .I(N__35173));
    InMux I__8472 (
            .O(N__35379),
            .I(N__35173));
    InMux I__8471 (
            .O(N__35378),
            .I(N__35173));
    InMux I__8470 (
            .O(N__35377),
            .I(N__35170));
    InMux I__8469 (
            .O(N__35376),
            .I(N__35167));
    InMux I__8468 (
            .O(N__35375),
            .I(N__35164));
    InMux I__8467 (
            .O(N__35374),
            .I(N__35159));
    InMux I__8466 (
            .O(N__35373),
            .I(N__35159));
    InMux I__8465 (
            .O(N__35372),
            .I(N__35152));
    InMux I__8464 (
            .O(N__35371),
            .I(N__35152));
    InMux I__8463 (
            .O(N__35370),
            .I(N__35152));
    LocalMux I__8462 (
            .O(N__35367),
            .I(N__35147));
    LocalMux I__8461 (
            .O(N__35358),
            .I(N__35147));
    InMux I__8460 (
            .O(N__35357),
            .I(N__35142));
    InMux I__8459 (
            .O(N__35356),
            .I(N__35142));
    LocalMux I__8458 (
            .O(N__35353),
            .I(N__35137));
    LocalMux I__8457 (
            .O(N__35350),
            .I(N__35137));
    LocalMux I__8456 (
            .O(N__35347),
            .I(N__35128));
    LocalMux I__8455 (
            .O(N__35342),
            .I(N__35128));
    LocalMux I__8454 (
            .O(N__35337),
            .I(N__35128));
    LocalMux I__8453 (
            .O(N__35332),
            .I(N__35128));
    InMux I__8452 (
            .O(N__35331),
            .I(N__35124));
    InMux I__8451 (
            .O(N__35330),
            .I(N__35121));
    InMux I__8450 (
            .O(N__35329),
            .I(N__35118));
    LocalMux I__8449 (
            .O(N__35326),
            .I(N__35115));
    LocalMux I__8448 (
            .O(N__35321),
            .I(N__35110));
    Span4Mux_s2_v I__8447 (
            .O(N__35318),
            .I(N__35110));
    LocalMux I__8446 (
            .O(N__35315),
            .I(N__35103));
    Span4Mux_v I__8445 (
            .O(N__35312),
            .I(N__35103));
    LocalMux I__8444 (
            .O(N__35305),
            .I(N__35103));
    LocalMux I__8443 (
            .O(N__35302),
            .I(N__35100));
    InMux I__8442 (
            .O(N__35301),
            .I(N__35095));
    InMux I__8441 (
            .O(N__35300),
            .I(N__35095));
    Span4Mux_v I__8440 (
            .O(N__35297),
            .I(N__35090));
    LocalMux I__8439 (
            .O(N__35288),
            .I(N__35090));
    LocalMux I__8438 (
            .O(N__35285),
            .I(N__35085));
    Span4Mux_v I__8437 (
            .O(N__35280),
            .I(N__35085));
    InMux I__8436 (
            .O(N__35279),
            .I(N__35080));
    InMux I__8435 (
            .O(N__35278),
            .I(N__35080));
    LocalMux I__8434 (
            .O(N__35273),
            .I(N__35077));
    InMux I__8433 (
            .O(N__35272),
            .I(N__35070));
    InMux I__8432 (
            .O(N__35269),
            .I(N__35070));
    InMux I__8431 (
            .O(N__35268),
            .I(N__35070));
    InMux I__8430 (
            .O(N__35267),
            .I(N__35067));
    InMux I__8429 (
            .O(N__35266),
            .I(N__35064));
    InMux I__8428 (
            .O(N__35265),
            .I(N__35061));
    InMux I__8427 (
            .O(N__35264),
            .I(N__35058));
    LocalMux I__8426 (
            .O(N__35261),
            .I(N__35054));
    InMux I__8425 (
            .O(N__35260),
            .I(N__35051));
    LocalMux I__8424 (
            .O(N__35257),
            .I(N__35044));
    Span4Mux_s2_h I__8423 (
            .O(N__35254),
            .I(N__35044));
    Span4Mux_v I__8422 (
            .O(N__35247),
            .I(N__35044));
    LocalMux I__8421 (
            .O(N__35242),
            .I(N__35039));
    LocalMux I__8420 (
            .O(N__35239),
            .I(N__35039));
    InMux I__8419 (
            .O(N__35238),
            .I(N__35034));
    InMux I__8418 (
            .O(N__35237),
            .I(N__35034));
    Span4Mux_h I__8417 (
            .O(N__35234),
            .I(N__35021));
    LocalMux I__8416 (
            .O(N__35229),
            .I(N__35021));
    Span4Mux_s3_v I__8415 (
            .O(N__35222),
            .I(N__35021));
    Span4Mux_h I__8414 (
            .O(N__35219),
            .I(N__35021));
    LocalMux I__8413 (
            .O(N__35214),
            .I(N__35021));
    LocalMux I__8412 (
            .O(N__35207),
            .I(N__35021));
    InMux I__8411 (
            .O(N__35206),
            .I(N__35018));
    LocalMux I__8410 (
            .O(N__35203),
            .I(N__35015));
    LocalMux I__8409 (
            .O(N__35200),
            .I(N__35012));
    InMux I__8408 (
            .O(N__35199),
            .I(N__35009));
    InMux I__8407 (
            .O(N__35198),
            .I(N__35006));
    LocalMux I__8406 (
            .O(N__35187),
            .I(N__34999));
    LocalMux I__8405 (
            .O(N__35180),
            .I(N__34999));
    LocalMux I__8404 (
            .O(N__35173),
            .I(N__34999));
    LocalMux I__8403 (
            .O(N__35170),
            .I(N__34986));
    LocalMux I__8402 (
            .O(N__35167),
            .I(N__34986));
    LocalMux I__8401 (
            .O(N__35164),
            .I(N__34986));
    LocalMux I__8400 (
            .O(N__35159),
            .I(N__34986));
    LocalMux I__8399 (
            .O(N__35152),
            .I(N__34986));
    Span4Mux_v I__8398 (
            .O(N__35147),
            .I(N__34986));
    LocalMux I__8397 (
            .O(N__35142),
            .I(N__34979));
    Span4Mux_v I__8396 (
            .O(N__35137),
            .I(N__34979));
    Span4Mux_v I__8395 (
            .O(N__35128),
            .I(N__34979));
    InMux I__8394 (
            .O(N__35127),
            .I(N__34976));
    LocalMux I__8393 (
            .O(N__35124),
            .I(N__34971));
    LocalMux I__8392 (
            .O(N__35121),
            .I(N__34971));
    LocalMux I__8391 (
            .O(N__35118),
            .I(N__34968));
    Span4Mux_v I__8390 (
            .O(N__35115),
            .I(N__34965));
    Span4Mux_v I__8389 (
            .O(N__35110),
            .I(N__34960));
    Span4Mux_h I__8388 (
            .O(N__35103),
            .I(N__34960));
    Span4Mux_s3_v I__8387 (
            .O(N__35100),
            .I(N__34949));
    LocalMux I__8386 (
            .O(N__35095),
            .I(N__34949));
    Span4Mux_s3_v I__8385 (
            .O(N__35090),
            .I(N__34949));
    Span4Mux_v I__8384 (
            .O(N__35085),
            .I(N__34949));
    LocalMux I__8383 (
            .O(N__35080),
            .I(N__34949));
    Span4Mux_v I__8382 (
            .O(N__35077),
            .I(N__34942));
    LocalMux I__8381 (
            .O(N__35070),
            .I(N__34942));
    LocalMux I__8380 (
            .O(N__35067),
            .I(N__34942));
    LocalMux I__8379 (
            .O(N__35064),
            .I(N__34935));
    LocalMux I__8378 (
            .O(N__35061),
            .I(N__34935));
    LocalMux I__8377 (
            .O(N__35058),
            .I(N__34935));
    CascadeMux I__8376 (
            .O(N__35057),
            .I(N__34932));
    Span4Mux_h I__8375 (
            .O(N__35054),
            .I(N__34927));
    LocalMux I__8374 (
            .O(N__35051),
            .I(N__34927));
    Span4Mux_h I__8373 (
            .O(N__35044),
            .I(N__34918));
    Span4Mux_v I__8372 (
            .O(N__35039),
            .I(N__34918));
    LocalMux I__8371 (
            .O(N__35034),
            .I(N__34918));
    Span4Mux_v I__8370 (
            .O(N__35021),
            .I(N__34918));
    LocalMux I__8369 (
            .O(N__35018),
            .I(N__34910));
    Span4Mux_s2_v I__8368 (
            .O(N__35015),
            .I(N__34910));
    Span4Mux_s2_v I__8367 (
            .O(N__35012),
            .I(N__34910));
    LocalMux I__8366 (
            .O(N__35009),
            .I(N__34907));
    LocalMux I__8365 (
            .O(N__35006),
            .I(N__34896));
    Span4Mux_s2_v I__8364 (
            .O(N__34999),
            .I(N__34896));
    Span4Mux_v I__8363 (
            .O(N__34986),
            .I(N__34896));
    Span4Mux_h I__8362 (
            .O(N__34979),
            .I(N__34896));
    LocalMux I__8361 (
            .O(N__34976),
            .I(N__34896));
    Span12Mux_s10_v I__8360 (
            .O(N__34971),
            .I(N__34893));
    Span4Mux_s3_v I__8359 (
            .O(N__34968),
            .I(N__34880));
    Span4Mux_v I__8358 (
            .O(N__34965),
            .I(N__34880));
    Span4Mux_v I__8357 (
            .O(N__34960),
            .I(N__34880));
    Span4Mux_h I__8356 (
            .O(N__34949),
            .I(N__34880));
    Span4Mux_s3_v I__8355 (
            .O(N__34942),
            .I(N__34880));
    Span4Mux_s3_v I__8354 (
            .O(N__34935),
            .I(N__34880));
    InMux I__8353 (
            .O(N__34932),
            .I(N__34877));
    Span4Mux_v I__8352 (
            .O(N__34927),
            .I(N__34872));
    Span4Mux_h I__8351 (
            .O(N__34918),
            .I(N__34872));
    InMux I__8350 (
            .O(N__34917),
            .I(N__34869));
    Span4Mux_h I__8349 (
            .O(N__34910),
            .I(N__34862));
    Span4Mux_v I__8348 (
            .O(N__34907),
            .I(N__34862));
    Span4Mux_h I__8347 (
            .O(N__34896),
            .I(N__34862));
    Odrv12 I__8346 (
            .O(N__34893),
            .I(\tok.T_6 ));
    Odrv4 I__8345 (
            .O(N__34880),
            .I(\tok.T_6 ));
    LocalMux I__8344 (
            .O(N__34877),
            .I(\tok.T_6 ));
    Odrv4 I__8343 (
            .O(N__34872),
            .I(\tok.T_6 ));
    LocalMux I__8342 (
            .O(N__34869),
            .I(\tok.T_6 ));
    Odrv4 I__8341 (
            .O(N__34862),
            .I(\tok.T_6 ));
    CascadeMux I__8340 (
            .O(N__34849),
            .I(\tok.n186_adj_812_cascade_ ));
    InMux I__8339 (
            .O(N__34846),
            .I(N__34835));
    InMux I__8338 (
            .O(N__34845),
            .I(N__34832));
    InMux I__8337 (
            .O(N__34844),
            .I(N__34827));
    InMux I__8336 (
            .O(N__34843),
            .I(N__34827));
    InMux I__8335 (
            .O(N__34842),
            .I(N__34822));
    InMux I__8334 (
            .O(N__34841),
            .I(N__34822));
    CascadeMux I__8333 (
            .O(N__34840),
            .I(N__34804));
    CascadeMux I__8332 (
            .O(N__34839),
            .I(N__34787));
    CascadeMux I__8331 (
            .O(N__34838),
            .I(N__34782));
    LocalMux I__8330 (
            .O(N__34835),
            .I(N__34773));
    LocalMux I__8329 (
            .O(N__34832),
            .I(N__34773));
    LocalMux I__8328 (
            .O(N__34827),
            .I(N__34768));
    LocalMux I__8327 (
            .O(N__34822),
            .I(N__34768));
    InMux I__8326 (
            .O(N__34821),
            .I(N__34765));
    InMux I__8325 (
            .O(N__34820),
            .I(N__34755));
    InMux I__8324 (
            .O(N__34819),
            .I(N__34743));
    InMux I__8323 (
            .O(N__34818),
            .I(N__34743));
    InMux I__8322 (
            .O(N__34817),
            .I(N__34743));
    InMux I__8321 (
            .O(N__34816),
            .I(N__34736));
    InMux I__8320 (
            .O(N__34815),
            .I(N__34736));
    InMux I__8319 (
            .O(N__34814),
            .I(N__34736));
    CascadeMux I__8318 (
            .O(N__34813),
            .I(N__34733));
    InMux I__8317 (
            .O(N__34812),
            .I(N__34730));
    InMux I__8316 (
            .O(N__34811),
            .I(N__34727));
    InMux I__8315 (
            .O(N__34810),
            .I(N__34724));
    InMux I__8314 (
            .O(N__34809),
            .I(N__34717));
    InMux I__8313 (
            .O(N__34808),
            .I(N__34717));
    InMux I__8312 (
            .O(N__34807),
            .I(N__34714));
    InMux I__8311 (
            .O(N__34804),
            .I(N__34707));
    CascadeMux I__8310 (
            .O(N__34803),
            .I(N__34701));
    InMux I__8309 (
            .O(N__34802),
            .I(N__34690));
    InMux I__8308 (
            .O(N__34801),
            .I(N__34690));
    InMux I__8307 (
            .O(N__34800),
            .I(N__34690));
    InMux I__8306 (
            .O(N__34799),
            .I(N__34683));
    InMux I__8305 (
            .O(N__34798),
            .I(N__34683));
    InMux I__8304 (
            .O(N__34797),
            .I(N__34683));
    CascadeMux I__8303 (
            .O(N__34796),
            .I(N__34677));
    InMux I__8302 (
            .O(N__34795),
            .I(N__34672));
    InMux I__8301 (
            .O(N__34794),
            .I(N__34665));
    InMux I__8300 (
            .O(N__34793),
            .I(N__34665));
    InMux I__8299 (
            .O(N__34792),
            .I(N__34665));
    CascadeMux I__8298 (
            .O(N__34791),
            .I(N__34662));
    InMux I__8297 (
            .O(N__34790),
            .I(N__34657));
    InMux I__8296 (
            .O(N__34787),
            .I(N__34654));
    InMux I__8295 (
            .O(N__34786),
            .I(N__34649));
    InMux I__8294 (
            .O(N__34785),
            .I(N__34649));
    InMux I__8293 (
            .O(N__34782),
            .I(N__34644));
    InMux I__8292 (
            .O(N__34781),
            .I(N__34644));
    CascadeMux I__8291 (
            .O(N__34780),
            .I(N__34640));
    InMux I__8290 (
            .O(N__34779),
            .I(N__34637));
    InMux I__8289 (
            .O(N__34778),
            .I(N__34634));
    Span4Mux_v I__8288 (
            .O(N__34773),
            .I(N__34627));
    Span4Mux_v I__8287 (
            .O(N__34768),
            .I(N__34627));
    LocalMux I__8286 (
            .O(N__34765),
            .I(N__34627));
    InMux I__8285 (
            .O(N__34764),
            .I(N__34624));
    InMux I__8284 (
            .O(N__34763),
            .I(N__34615));
    InMux I__8283 (
            .O(N__34762),
            .I(N__34615));
    InMux I__8282 (
            .O(N__34761),
            .I(N__34615));
    InMux I__8281 (
            .O(N__34760),
            .I(N__34615));
    CascadeMux I__8280 (
            .O(N__34759),
            .I(N__34607));
    CascadeMux I__8279 (
            .O(N__34758),
            .I(N__34603));
    LocalMux I__8278 (
            .O(N__34755),
            .I(N__34600));
    InMux I__8277 (
            .O(N__34754),
            .I(N__34595));
    InMux I__8276 (
            .O(N__34753),
            .I(N__34595));
    InMux I__8275 (
            .O(N__34752),
            .I(N__34590));
    InMux I__8274 (
            .O(N__34751),
            .I(N__34590));
    InMux I__8273 (
            .O(N__34750),
            .I(N__34587));
    LocalMux I__8272 (
            .O(N__34743),
            .I(N__34582));
    LocalMux I__8271 (
            .O(N__34736),
            .I(N__34582));
    InMux I__8270 (
            .O(N__34733),
            .I(N__34579));
    LocalMux I__8269 (
            .O(N__34730),
            .I(N__34574));
    LocalMux I__8268 (
            .O(N__34727),
            .I(N__34574));
    LocalMux I__8267 (
            .O(N__34724),
            .I(N__34571));
    InMux I__8266 (
            .O(N__34723),
            .I(N__34566));
    InMux I__8265 (
            .O(N__34722),
            .I(N__34566));
    LocalMux I__8264 (
            .O(N__34717),
            .I(N__34561));
    LocalMux I__8263 (
            .O(N__34714),
            .I(N__34561));
    CascadeMux I__8262 (
            .O(N__34713),
            .I(N__34555));
    CascadeMux I__8261 (
            .O(N__34712),
            .I(N__34552));
    CascadeMux I__8260 (
            .O(N__34711),
            .I(N__34548));
    InMux I__8259 (
            .O(N__34710),
            .I(N__34544));
    LocalMux I__8258 (
            .O(N__34707),
            .I(N__34541));
    CascadeMux I__8257 (
            .O(N__34706),
            .I(N__34538));
    InMux I__8256 (
            .O(N__34705),
            .I(N__34532));
    InMux I__8255 (
            .O(N__34704),
            .I(N__34529));
    InMux I__8254 (
            .O(N__34701),
            .I(N__34524));
    InMux I__8253 (
            .O(N__34700),
            .I(N__34518));
    InMux I__8252 (
            .O(N__34699),
            .I(N__34518));
    InMux I__8251 (
            .O(N__34698),
            .I(N__34515));
    InMux I__8250 (
            .O(N__34697),
            .I(N__34511));
    LocalMux I__8249 (
            .O(N__34690),
            .I(N__34506));
    LocalMux I__8248 (
            .O(N__34683),
            .I(N__34506));
    InMux I__8247 (
            .O(N__34682),
            .I(N__34497));
    InMux I__8246 (
            .O(N__34681),
            .I(N__34497));
    InMux I__8245 (
            .O(N__34680),
            .I(N__34497));
    InMux I__8244 (
            .O(N__34677),
            .I(N__34497));
    InMux I__8243 (
            .O(N__34676),
            .I(N__34492));
    InMux I__8242 (
            .O(N__34675),
            .I(N__34492));
    LocalMux I__8241 (
            .O(N__34672),
            .I(N__34487));
    LocalMux I__8240 (
            .O(N__34665),
            .I(N__34487));
    InMux I__8239 (
            .O(N__34662),
            .I(N__34484));
    InMux I__8238 (
            .O(N__34661),
            .I(N__34476));
    InMux I__8237 (
            .O(N__34660),
            .I(N__34476));
    LocalMux I__8236 (
            .O(N__34657),
            .I(N__34467));
    LocalMux I__8235 (
            .O(N__34654),
            .I(N__34467));
    LocalMux I__8234 (
            .O(N__34649),
            .I(N__34467));
    LocalMux I__8233 (
            .O(N__34644),
            .I(N__34467));
    InMux I__8232 (
            .O(N__34643),
            .I(N__34462));
    InMux I__8231 (
            .O(N__34640),
            .I(N__34462));
    LocalMux I__8230 (
            .O(N__34637),
            .I(N__34451));
    LocalMux I__8229 (
            .O(N__34634),
            .I(N__34451));
    Span4Mux_h I__8228 (
            .O(N__34627),
            .I(N__34451));
    LocalMux I__8227 (
            .O(N__34624),
            .I(N__34451));
    LocalMux I__8226 (
            .O(N__34615),
            .I(N__34448));
    InMux I__8225 (
            .O(N__34614),
            .I(N__34443));
    InMux I__8224 (
            .O(N__34613),
            .I(N__34443));
    InMux I__8223 (
            .O(N__34612),
            .I(N__34436));
    InMux I__8222 (
            .O(N__34611),
            .I(N__34436));
    InMux I__8221 (
            .O(N__34610),
            .I(N__34436));
    InMux I__8220 (
            .O(N__34607),
            .I(N__34429));
    InMux I__8219 (
            .O(N__34606),
            .I(N__34429));
    InMux I__8218 (
            .O(N__34603),
            .I(N__34429));
    Span4Mux_h I__8217 (
            .O(N__34600),
            .I(N__34425));
    LocalMux I__8216 (
            .O(N__34595),
            .I(N__34420));
    LocalMux I__8215 (
            .O(N__34590),
            .I(N__34420));
    LocalMux I__8214 (
            .O(N__34587),
            .I(N__34415));
    Span4Mux_v I__8213 (
            .O(N__34582),
            .I(N__34415));
    LocalMux I__8212 (
            .O(N__34579),
            .I(N__34404));
    Span4Mux_v I__8211 (
            .O(N__34574),
            .I(N__34404));
    Span4Mux_s2_h I__8210 (
            .O(N__34571),
            .I(N__34404));
    LocalMux I__8209 (
            .O(N__34566),
            .I(N__34404));
    Span4Mux_s2_h I__8208 (
            .O(N__34561),
            .I(N__34404));
    CascadeMux I__8207 (
            .O(N__34560),
            .I(N__34401));
    CascadeMux I__8206 (
            .O(N__34559),
            .I(N__34398));
    InMux I__8205 (
            .O(N__34558),
            .I(N__34394));
    InMux I__8204 (
            .O(N__34555),
            .I(N__34391));
    InMux I__8203 (
            .O(N__34552),
            .I(N__34384));
    InMux I__8202 (
            .O(N__34551),
            .I(N__34384));
    InMux I__8201 (
            .O(N__34548),
            .I(N__34384));
    InMux I__8200 (
            .O(N__34547),
            .I(N__34381));
    LocalMux I__8199 (
            .O(N__34544),
            .I(N__34376));
    Span4Mux_s3_v I__8198 (
            .O(N__34541),
            .I(N__34376));
    InMux I__8197 (
            .O(N__34538),
            .I(N__34371));
    InMux I__8196 (
            .O(N__34537),
            .I(N__34371));
    InMux I__8195 (
            .O(N__34536),
            .I(N__34368));
    InMux I__8194 (
            .O(N__34535),
            .I(N__34365));
    LocalMux I__8193 (
            .O(N__34532),
            .I(N__34360));
    LocalMux I__8192 (
            .O(N__34529),
            .I(N__34360));
    InMux I__8191 (
            .O(N__34528),
            .I(N__34355));
    InMux I__8190 (
            .O(N__34527),
            .I(N__34355));
    LocalMux I__8189 (
            .O(N__34524),
            .I(N__34352));
    InMux I__8188 (
            .O(N__34523),
            .I(N__34349));
    LocalMux I__8187 (
            .O(N__34518),
            .I(N__34344));
    LocalMux I__8186 (
            .O(N__34515),
            .I(N__34344));
    InMux I__8185 (
            .O(N__34514),
            .I(N__34341));
    LocalMux I__8184 (
            .O(N__34511),
            .I(N__34334));
    Span4Mux_v I__8183 (
            .O(N__34506),
            .I(N__34334));
    LocalMux I__8182 (
            .O(N__34497),
            .I(N__34334));
    LocalMux I__8181 (
            .O(N__34492),
            .I(N__34331));
    Span4Mux_s1_v I__8180 (
            .O(N__34487),
            .I(N__34326));
    LocalMux I__8179 (
            .O(N__34484),
            .I(N__34326));
    InMux I__8178 (
            .O(N__34483),
            .I(N__34321));
    InMux I__8177 (
            .O(N__34482),
            .I(N__34321));
    InMux I__8176 (
            .O(N__34481),
            .I(N__34318));
    LocalMux I__8175 (
            .O(N__34476),
            .I(N__34311));
    Span4Mux_h I__8174 (
            .O(N__34467),
            .I(N__34311));
    LocalMux I__8173 (
            .O(N__34462),
            .I(N__34311));
    InMux I__8172 (
            .O(N__34461),
            .I(N__34308));
    InMux I__8171 (
            .O(N__34460),
            .I(N__34305));
    Span4Mux_v I__8170 (
            .O(N__34451),
            .I(N__34300));
    Span4Mux_v I__8169 (
            .O(N__34448),
            .I(N__34300));
    LocalMux I__8168 (
            .O(N__34443),
            .I(N__34293));
    LocalMux I__8167 (
            .O(N__34436),
            .I(N__34293));
    LocalMux I__8166 (
            .O(N__34429),
            .I(N__34293));
    CascadeMux I__8165 (
            .O(N__34428),
            .I(N__34290));
    Span4Mux_v I__8164 (
            .O(N__34425),
            .I(N__34281));
    Span4Mux_v I__8163 (
            .O(N__34420),
            .I(N__34281));
    Span4Mux_h I__8162 (
            .O(N__34415),
            .I(N__34281));
    Span4Mux_h I__8161 (
            .O(N__34404),
            .I(N__34281));
    InMux I__8160 (
            .O(N__34401),
            .I(N__34276));
    InMux I__8159 (
            .O(N__34398),
            .I(N__34276));
    InMux I__8158 (
            .O(N__34397),
            .I(N__34261));
    LocalMux I__8157 (
            .O(N__34394),
            .I(N__34258));
    LocalMux I__8156 (
            .O(N__34391),
            .I(N__34253));
    LocalMux I__8155 (
            .O(N__34384),
            .I(N__34253));
    LocalMux I__8154 (
            .O(N__34381),
            .I(N__34246));
    Span4Mux_v I__8153 (
            .O(N__34376),
            .I(N__34246));
    LocalMux I__8152 (
            .O(N__34371),
            .I(N__34246));
    LocalMux I__8151 (
            .O(N__34368),
            .I(N__34237));
    LocalMux I__8150 (
            .O(N__34365),
            .I(N__34237));
    Span4Mux_v I__8149 (
            .O(N__34360),
            .I(N__34237));
    LocalMux I__8148 (
            .O(N__34355),
            .I(N__34237));
    Span4Mux_v I__8147 (
            .O(N__34352),
            .I(N__34226));
    LocalMux I__8146 (
            .O(N__34349),
            .I(N__34226));
    Span4Mux_s3_h I__8145 (
            .O(N__34344),
            .I(N__34226));
    LocalMux I__8144 (
            .O(N__34341),
            .I(N__34226));
    Span4Mux_v I__8143 (
            .O(N__34334),
            .I(N__34226));
    Span4Mux_h I__8142 (
            .O(N__34331),
            .I(N__34219));
    Span4Mux_v I__8141 (
            .O(N__34326),
            .I(N__34219));
    LocalMux I__8140 (
            .O(N__34321),
            .I(N__34219));
    LocalMux I__8139 (
            .O(N__34318),
            .I(N__34212));
    Span4Mux_h I__8138 (
            .O(N__34311),
            .I(N__34212));
    LocalMux I__8137 (
            .O(N__34308),
            .I(N__34212));
    LocalMux I__8136 (
            .O(N__34305),
            .I(N__34205));
    Span4Mux_h I__8135 (
            .O(N__34300),
            .I(N__34205));
    Span4Mux_v I__8134 (
            .O(N__34293),
            .I(N__34205));
    InMux I__8133 (
            .O(N__34290),
            .I(N__34202));
    Span4Mux_h I__8132 (
            .O(N__34281),
            .I(N__34197));
    LocalMux I__8131 (
            .O(N__34276),
            .I(N__34197));
    InMux I__8130 (
            .O(N__34275),
            .I(N__34190));
    InMux I__8129 (
            .O(N__34274),
            .I(N__34190));
    InMux I__8128 (
            .O(N__34273),
            .I(N__34190));
    InMux I__8127 (
            .O(N__34272),
            .I(N__34185));
    InMux I__8126 (
            .O(N__34271),
            .I(N__34185));
    InMux I__8125 (
            .O(N__34270),
            .I(N__34176));
    InMux I__8124 (
            .O(N__34269),
            .I(N__34176));
    InMux I__8123 (
            .O(N__34268),
            .I(N__34176));
    InMux I__8122 (
            .O(N__34267),
            .I(N__34176));
    InMux I__8121 (
            .O(N__34266),
            .I(N__34169));
    InMux I__8120 (
            .O(N__34265),
            .I(N__34169));
    InMux I__8119 (
            .O(N__34264),
            .I(N__34169));
    LocalMux I__8118 (
            .O(N__34261),
            .I(N__34156));
    Span4Mux_s2_v I__8117 (
            .O(N__34258),
            .I(N__34156));
    Span4Mux_v I__8116 (
            .O(N__34253),
            .I(N__34156));
    Span4Mux_v I__8115 (
            .O(N__34246),
            .I(N__34156));
    Span4Mux_v I__8114 (
            .O(N__34237),
            .I(N__34156));
    Span4Mux_h I__8113 (
            .O(N__34226),
            .I(N__34156));
    Span4Mux_h I__8112 (
            .O(N__34219),
            .I(N__34149));
    Span4Mux_v I__8111 (
            .O(N__34212),
            .I(N__34149));
    Span4Mux_h I__8110 (
            .O(N__34205),
            .I(N__34149));
    LocalMux I__8109 (
            .O(N__34202),
            .I(N__34144));
    Span4Mux_v I__8108 (
            .O(N__34197),
            .I(N__34144));
    LocalMux I__8107 (
            .O(N__34190),
            .I(\tok.T_3 ));
    LocalMux I__8106 (
            .O(N__34185),
            .I(\tok.T_3 ));
    LocalMux I__8105 (
            .O(N__34176),
            .I(\tok.T_3 ));
    LocalMux I__8104 (
            .O(N__34169),
            .I(\tok.T_3 ));
    Odrv4 I__8103 (
            .O(N__34156),
            .I(\tok.T_3 ));
    Odrv4 I__8102 (
            .O(N__34149),
            .I(\tok.T_3 ));
    Odrv4 I__8101 (
            .O(N__34144),
            .I(\tok.T_3 ));
    InMux I__8100 (
            .O(N__34129),
            .I(N__34126));
    LocalMux I__8099 (
            .O(N__34126),
            .I(N__34123));
    Span4Mux_h I__8098 (
            .O(N__34123),
            .I(N__34120));
    Span4Mux_h I__8097 (
            .O(N__34120),
            .I(N__34117));
    Odrv4 I__8096 (
            .O(N__34117),
            .I(\tok.n338_adj_819 ));
    CascadeMux I__8095 (
            .O(N__34114),
            .I(N__34109));
    CascadeMux I__8094 (
            .O(N__34113),
            .I(N__34097));
    CascadeMux I__8093 (
            .O(N__34112),
            .I(N__34089));
    InMux I__8092 (
            .O(N__34109),
            .I(N__34084));
    InMux I__8091 (
            .O(N__34108),
            .I(N__34084));
    InMux I__8090 (
            .O(N__34107),
            .I(N__34072));
    InMux I__8089 (
            .O(N__34106),
            .I(N__34064));
    InMux I__8088 (
            .O(N__34105),
            .I(N__34064));
    CascadeMux I__8087 (
            .O(N__34104),
            .I(N__34056));
    CascadeMux I__8086 (
            .O(N__34103),
            .I(N__34049));
    CascadeMux I__8085 (
            .O(N__34102),
            .I(N__34042));
    CascadeMux I__8084 (
            .O(N__34101),
            .I(N__34037));
    CascadeMux I__8083 (
            .O(N__34100),
            .I(N__34032));
    InMux I__8082 (
            .O(N__34097),
            .I(N__34027));
    CascadeMux I__8081 (
            .O(N__34096),
            .I(N__34023));
    InMux I__8080 (
            .O(N__34095),
            .I(N__34020));
    InMux I__8079 (
            .O(N__34094),
            .I(N__34017));
    InMux I__8078 (
            .O(N__34093),
            .I(N__34012));
    InMux I__8077 (
            .O(N__34092),
            .I(N__34012));
    InMux I__8076 (
            .O(N__34089),
            .I(N__34009));
    LocalMux I__8075 (
            .O(N__34084),
            .I(N__34006));
    InMux I__8074 (
            .O(N__34083),
            .I(N__33996));
    InMux I__8073 (
            .O(N__34082),
            .I(N__33996));
    InMux I__8072 (
            .O(N__34081),
            .I(N__33996));
    CascadeMux I__8071 (
            .O(N__34080),
            .I(N__33991));
    CascadeMux I__8070 (
            .O(N__34079),
            .I(N__33988));
    InMux I__8069 (
            .O(N__34078),
            .I(N__33981));
    InMux I__8068 (
            .O(N__34077),
            .I(N__33981));
    InMux I__8067 (
            .O(N__34076),
            .I(N__33974));
    InMux I__8066 (
            .O(N__34075),
            .I(N__33974));
    LocalMux I__8065 (
            .O(N__34072),
            .I(N__33971));
    InMux I__8064 (
            .O(N__34071),
            .I(N__33968));
    InMux I__8063 (
            .O(N__34070),
            .I(N__33963));
    InMux I__8062 (
            .O(N__34069),
            .I(N__33963));
    LocalMux I__8061 (
            .O(N__34064),
            .I(N__33960));
    InMux I__8060 (
            .O(N__34063),
            .I(N__33953));
    InMux I__8059 (
            .O(N__34062),
            .I(N__33953));
    InMux I__8058 (
            .O(N__34061),
            .I(N__33953));
    CascadeMux I__8057 (
            .O(N__34060),
            .I(N__33947));
    InMux I__8056 (
            .O(N__34059),
            .I(N__33942));
    InMux I__8055 (
            .O(N__34056),
            .I(N__33937));
    InMux I__8054 (
            .O(N__34055),
            .I(N__33937));
    InMux I__8053 (
            .O(N__34054),
            .I(N__33931));
    InMux I__8052 (
            .O(N__34053),
            .I(N__33926));
    InMux I__8051 (
            .O(N__34052),
            .I(N__33926));
    InMux I__8050 (
            .O(N__34049),
            .I(N__33923));
    InMux I__8049 (
            .O(N__34048),
            .I(N__33916));
    InMux I__8048 (
            .O(N__34047),
            .I(N__33916));
    InMux I__8047 (
            .O(N__34046),
            .I(N__33916));
    InMux I__8046 (
            .O(N__34045),
            .I(N__33909));
    InMux I__8045 (
            .O(N__34042),
            .I(N__33909));
    InMux I__8044 (
            .O(N__34041),
            .I(N__33909));
    InMux I__8043 (
            .O(N__34040),
            .I(N__33906));
    InMux I__8042 (
            .O(N__34037),
            .I(N__33899));
    InMux I__8041 (
            .O(N__34036),
            .I(N__33899));
    InMux I__8040 (
            .O(N__34035),
            .I(N__33899));
    InMux I__8039 (
            .O(N__34032),
            .I(N__33892));
    InMux I__8038 (
            .O(N__34031),
            .I(N__33892));
    InMux I__8037 (
            .O(N__34030),
            .I(N__33892));
    LocalMux I__8036 (
            .O(N__34027),
            .I(N__33889));
    InMux I__8035 (
            .O(N__34026),
            .I(N__33884));
    InMux I__8034 (
            .O(N__34023),
            .I(N__33884));
    LocalMux I__8033 (
            .O(N__34020),
            .I(N__33873));
    LocalMux I__8032 (
            .O(N__34017),
            .I(N__33873));
    LocalMux I__8031 (
            .O(N__34012),
            .I(N__33873));
    LocalMux I__8030 (
            .O(N__34009),
            .I(N__33873));
    Span4Mux_v I__8029 (
            .O(N__34006),
            .I(N__33873));
    InMux I__8028 (
            .O(N__34005),
            .I(N__33868));
    InMux I__8027 (
            .O(N__34004),
            .I(N__33863));
    InMux I__8026 (
            .O(N__34003),
            .I(N__33863));
    LocalMux I__8025 (
            .O(N__33996),
            .I(N__33860));
    InMux I__8024 (
            .O(N__33995),
            .I(N__33857));
    InMux I__8023 (
            .O(N__33994),
            .I(N__33848));
    InMux I__8022 (
            .O(N__33991),
            .I(N__33848));
    InMux I__8021 (
            .O(N__33988),
            .I(N__33848));
    InMux I__8020 (
            .O(N__33987),
            .I(N__33848));
    InMux I__8019 (
            .O(N__33986),
            .I(N__33845));
    LocalMux I__8018 (
            .O(N__33981),
            .I(N__33842));
    InMux I__8017 (
            .O(N__33980),
            .I(N__33837));
    InMux I__8016 (
            .O(N__33979),
            .I(N__33837));
    LocalMux I__8015 (
            .O(N__33974),
            .I(N__33834));
    Span4Mux_v I__8014 (
            .O(N__33971),
            .I(N__33827));
    LocalMux I__8013 (
            .O(N__33968),
            .I(N__33827));
    LocalMux I__8012 (
            .O(N__33963),
            .I(N__33827));
    Span4Mux_v I__8011 (
            .O(N__33960),
            .I(N__33822));
    LocalMux I__8010 (
            .O(N__33953),
            .I(N__33822));
    InMux I__8009 (
            .O(N__33952),
            .I(N__33813));
    InMux I__8008 (
            .O(N__33951),
            .I(N__33813));
    InMux I__8007 (
            .O(N__33950),
            .I(N__33813));
    InMux I__8006 (
            .O(N__33947),
            .I(N__33813));
    InMux I__8005 (
            .O(N__33946),
            .I(N__33808));
    InMux I__8004 (
            .O(N__33945),
            .I(N__33808));
    LocalMux I__8003 (
            .O(N__33942),
            .I(N__33803));
    LocalMux I__8002 (
            .O(N__33937),
            .I(N__33803));
    InMux I__8001 (
            .O(N__33936),
            .I(N__33799));
    InMux I__8000 (
            .O(N__33935),
            .I(N__33792));
    InMux I__7999 (
            .O(N__33934),
            .I(N__33792));
    LocalMux I__7998 (
            .O(N__33931),
            .I(N__33789));
    LocalMux I__7997 (
            .O(N__33926),
            .I(N__33786));
    LocalMux I__7996 (
            .O(N__33923),
            .I(N__33779));
    LocalMux I__7995 (
            .O(N__33916),
            .I(N__33779));
    LocalMux I__7994 (
            .O(N__33909),
            .I(N__33779));
    LocalMux I__7993 (
            .O(N__33906),
            .I(N__33770));
    LocalMux I__7992 (
            .O(N__33899),
            .I(N__33770));
    LocalMux I__7991 (
            .O(N__33892),
            .I(N__33770));
    Span4Mux_v I__7990 (
            .O(N__33889),
            .I(N__33770));
    LocalMux I__7989 (
            .O(N__33884),
            .I(N__33765));
    Span4Mux_v I__7988 (
            .O(N__33873),
            .I(N__33765));
    InMux I__7987 (
            .O(N__33872),
            .I(N__33760));
    InMux I__7986 (
            .O(N__33871),
            .I(N__33760));
    LocalMux I__7985 (
            .O(N__33868),
            .I(N__33757));
    LocalMux I__7984 (
            .O(N__33863),
            .I(N__33754));
    Span4Mux_v I__7983 (
            .O(N__33860),
            .I(N__33751));
    LocalMux I__7982 (
            .O(N__33857),
            .I(N__33746));
    LocalMux I__7981 (
            .O(N__33848),
            .I(N__33746));
    LocalMux I__7980 (
            .O(N__33845),
            .I(N__33733));
    Span4Mux_s3_h I__7979 (
            .O(N__33842),
            .I(N__33733));
    LocalMux I__7978 (
            .O(N__33837),
            .I(N__33733));
    Span4Mux_v I__7977 (
            .O(N__33834),
            .I(N__33733));
    Span4Mux_s3_v I__7976 (
            .O(N__33827),
            .I(N__33733));
    Span4Mux_v I__7975 (
            .O(N__33822),
            .I(N__33733));
    LocalMux I__7974 (
            .O(N__33813),
            .I(N__33730));
    LocalMux I__7973 (
            .O(N__33808),
            .I(N__33727));
    Span4Mux_v I__7972 (
            .O(N__33803),
            .I(N__33724));
    InMux I__7971 (
            .O(N__33802),
            .I(N__33721));
    LocalMux I__7970 (
            .O(N__33799),
            .I(N__33718));
    InMux I__7969 (
            .O(N__33798),
            .I(N__33715));
    CascadeMux I__7968 (
            .O(N__33797),
            .I(N__33712));
    LocalMux I__7967 (
            .O(N__33792),
            .I(N__33696));
    Span4Mux_s2_v I__7966 (
            .O(N__33789),
            .I(N__33696));
    Span4Mux_h I__7965 (
            .O(N__33786),
            .I(N__33696));
    Span4Mux_s2_v I__7964 (
            .O(N__33779),
            .I(N__33696));
    Span4Mux_v I__7963 (
            .O(N__33770),
            .I(N__33696));
    Span4Mux_h I__7962 (
            .O(N__33765),
            .I(N__33696));
    LocalMux I__7961 (
            .O(N__33760),
            .I(N__33696));
    Span4Mux_h I__7960 (
            .O(N__33757),
            .I(N__33693));
    Span4Mux_s3_v I__7959 (
            .O(N__33754),
            .I(N__33682));
    Span4Mux_v I__7958 (
            .O(N__33751),
            .I(N__33682));
    Span4Mux_s3_v I__7957 (
            .O(N__33746),
            .I(N__33682));
    Span4Mux_h I__7956 (
            .O(N__33733),
            .I(N__33682));
    Span4Mux_s3_v I__7955 (
            .O(N__33730),
            .I(N__33682));
    Span4Mux_h I__7954 (
            .O(N__33727),
            .I(N__33675));
    Span4Mux_h I__7953 (
            .O(N__33724),
            .I(N__33675));
    LocalMux I__7952 (
            .O(N__33721),
            .I(N__33675));
    Span4Mux_s3_v I__7951 (
            .O(N__33718),
            .I(N__33670));
    LocalMux I__7950 (
            .O(N__33715),
            .I(N__33670));
    InMux I__7949 (
            .O(N__33712),
            .I(N__33667));
    InMux I__7948 (
            .O(N__33711),
            .I(N__33664));
    Span4Mux_h I__7947 (
            .O(N__33696),
            .I(N__33661));
    Odrv4 I__7946 (
            .O(N__33693),
            .I(\tok.T_7 ));
    Odrv4 I__7945 (
            .O(N__33682),
            .I(\tok.T_7 ));
    Odrv4 I__7944 (
            .O(N__33675),
            .I(\tok.T_7 ));
    Odrv4 I__7943 (
            .O(N__33670),
            .I(\tok.T_7 ));
    LocalMux I__7942 (
            .O(N__33667),
            .I(\tok.T_7 ));
    LocalMux I__7941 (
            .O(N__33664),
            .I(\tok.T_7 ));
    Odrv4 I__7940 (
            .O(N__33661),
            .I(\tok.T_7 ));
    CascadeMux I__7939 (
            .O(N__33646),
            .I(N__33639));
    CascadeMux I__7938 (
            .O(N__33645),
            .I(N__33636));
    InMux I__7937 (
            .O(N__33644),
            .I(N__33629));
    InMux I__7936 (
            .O(N__33643),
            .I(N__33626));
    InMux I__7935 (
            .O(N__33642),
            .I(N__33622));
    InMux I__7934 (
            .O(N__33639),
            .I(N__33619));
    InMux I__7933 (
            .O(N__33636),
            .I(N__33616));
    InMux I__7932 (
            .O(N__33635),
            .I(N__33611));
    InMux I__7931 (
            .O(N__33634),
            .I(N__33611));
    InMux I__7930 (
            .O(N__33633),
            .I(N__33604));
    InMux I__7929 (
            .O(N__33632),
            .I(N__33601));
    LocalMux I__7928 (
            .O(N__33629),
            .I(N__33598));
    LocalMux I__7927 (
            .O(N__33626),
            .I(N__33594));
    InMux I__7926 (
            .O(N__33625),
            .I(N__33591));
    LocalMux I__7925 (
            .O(N__33622),
            .I(N__33586));
    LocalMux I__7924 (
            .O(N__33619),
            .I(N__33586));
    LocalMux I__7923 (
            .O(N__33616),
            .I(N__33583));
    LocalMux I__7922 (
            .O(N__33611),
            .I(N__33578));
    InMux I__7921 (
            .O(N__33610),
            .I(N__33571));
    InMux I__7920 (
            .O(N__33609),
            .I(N__33571));
    InMux I__7919 (
            .O(N__33608),
            .I(N__33571));
    InMux I__7918 (
            .O(N__33607),
            .I(N__33568));
    LocalMux I__7917 (
            .O(N__33604),
            .I(N__33565));
    LocalMux I__7916 (
            .O(N__33601),
            .I(N__33558));
    Span4Mux_v I__7915 (
            .O(N__33598),
            .I(N__33555));
    InMux I__7914 (
            .O(N__33597),
            .I(N__33552));
    Span4Mux_v I__7913 (
            .O(N__33594),
            .I(N__33547));
    LocalMux I__7912 (
            .O(N__33591),
            .I(N__33547));
    Span4Mux_v I__7911 (
            .O(N__33586),
            .I(N__33542));
    Span4Mux_v I__7910 (
            .O(N__33583),
            .I(N__33542));
    InMux I__7909 (
            .O(N__33582),
            .I(N__33539));
    InMux I__7908 (
            .O(N__33581),
            .I(N__33536));
    Span4Mux_h I__7907 (
            .O(N__33578),
            .I(N__33533));
    LocalMux I__7906 (
            .O(N__33571),
            .I(N__33530));
    LocalMux I__7905 (
            .O(N__33568),
            .I(N__33525));
    Span12Mux_s5_v I__7904 (
            .O(N__33565),
            .I(N__33525));
    InMux I__7903 (
            .O(N__33564),
            .I(N__33516));
    InMux I__7902 (
            .O(N__33563),
            .I(N__33516));
    InMux I__7901 (
            .O(N__33562),
            .I(N__33516));
    InMux I__7900 (
            .O(N__33561),
            .I(N__33516));
    Span4Mux_v I__7899 (
            .O(N__33558),
            .I(N__33505));
    Span4Mux_h I__7898 (
            .O(N__33555),
            .I(N__33505));
    LocalMux I__7897 (
            .O(N__33552),
            .I(N__33505));
    Span4Mux_h I__7896 (
            .O(N__33547),
            .I(N__33505));
    Span4Mux_h I__7895 (
            .O(N__33542),
            .I(N__33505));
    LocalMux I__7894 (
            .O(N__33539),
            .I(\tok.A_low_2 ));
    LocalMux I__7893 (
            .O(N__33536),
            .I(\tok.A_low_2 ));
    Odrv4 I__7892 (
            .O(N__33533),
            .I(\tok.A_low_2 ));
    Odrv12 I__7891 (
            .O(N__33530),
            .I(\tok.A_low_2 ));
    Odrv12 I__7890 (
            .O(N__33525),
            .I(\tok.A_low_2 ));
    LocalMux I__7889 (
            .O(N__33516),
            .I(\tok.A_low_2 ));
    Odrv4 I__7888 (
            .O(N__33505),
            .I(\tok.A_low_2 ));
    InMux I__7887 (
            .O(N__33490),
            .I(N__33486));
    CascadeMux I__7886 (
            .O(N__33489),
            .I(N__33480));
    LocalMux I__7885 (
            .O(N__33486),
            .I(N__33476));
    InMux I__7884 (
            .O(N__33485),
            .I(N__33472));
    InMux I__7883 (
            .O(N__33484),
            .I(N__33468));
    CascadeMux I__7882 (
            .O(N__33483),
            .I(N__33464));
    InMux I__7881 (
            .O(N__33480),
            .I(N__33461));
    InMux I__7880 (
            .O(N__33479),
            .I(N__33458));
    Span4Mux_v I__7879 (
            .O(N__33476),
            .I(N__33455));
    InMux I__7878 (
            .O(N__33475),
            .I(N__33452));
    LocalMux I__7877 (
            .O(N__33472),
            .I(N__33449));
    InMux I__7876 (
            .O(N__33471),
            .I(N__33446));
    LocalMux I__7875 (
            .O(N__33468),
            .I(N__33442));
    InMux I__7874 (
            .O(N__33467),
            .I(N__33439));
    InMux I__7873 (
            .O(N__33464),
            .I(N__33436));
    LocalMux I__7872 (
            .O(N__33461),
            .I(N__33433));
    LocalMux I__7871 (
            .O(N__33458),
            .I(N__33421));
    Span4Mux_h I__7870 (
            .O(N__33455),
            .I(N__33421));
    LocalMux I__7869 (
            .O(N__33452),
            .I(N__33421));
    Span4Mux_v I__7868 (
            .O(N__33449),
            .I(N__33418));
    LocalMux I__7867 (
            .O(N__33446),
            .I(N__33411));
    InMux I__7866 (
            .O(N__33445),
            .I(N__33408));
    Span4Mux_s3_v I__7865 (
            .O(N__33442),
            .I(N__33405));
    LocalMux I__7864 (
            .O(N__33439),
            .I(N__33400));
    LocalMux I__7863 (
            .O(N__33436),
            .I(N__33400));
    Span4Mux_v I__7862 (
            .O(N__33433),
            .I(N__33397));
    InMux I__7861 (
            .O(N__33432),
            .I(N__33394));
    InMux I__7860 (
            .O(N__33431),
            .I(N__33391));
    InMux I__7859 (
            .O(N__33430),
            .I(N__33388));
    InMux I__7858 (
            .O(N__33429),
            .I(N__33383));
    InMux I__7857 (
            .O(N__33428),
            .I(N__33383));
    Span4Mux_v I__7856 (
            .O(N__33421),
            .I(N__33378));
    Span4Mux_v I__7855 (
            .O(N__33418),
            .I(N__33378));
    InMux I__7854 (
            .O(N__33417),
            .I(N__33373));
    InMux I__7853 (
            .O(N__33416),
            .I(N__33373));
    InMux I__7852 (
            .O(N__33415),
            .I(N__33368));
    InMux I__7851 (
            .O(N__33414),
            .I(N__33365));
    Span4Mux_s3_v I__7850 (
            .O(N__33411),
            .I(N__33362));
    LocalMux I__7849 (
            .O(N__33408),
            .I(N__33359));
    Span4Mux_s3_h I__7848 (
            .O(N__33405),
            .I(N__33352));
    Span4Mux_s3_h I__7847 (
            .O(N__33400),
            .I(N__33352));
    Span4Mux_v I__7846 (
            .O(N__33397),
            .I(N__33352));
    LocalMux I__7845 (
            .O(N__33394),
            .I(N__33347));
    LocalMux I__7844 (
            .O(N__33391),
            .I(N__33347));
    LocalMux I__7843 (
            .O(N__33388),
            .I(N__33344));
    LocalMux I__7842 (
            .O(N__33383),
            .I(N__33337));
    Sp12to4 I__7841 (
            .O(N__33378),
            .I(N__33337));
    LocalMux I__7840 (
            .O(N__33373),
            .I(N__33337));
    InMux I__7839 (
            .O(N__33372),
            .I(N__33334));
    InMux I__7838 (
            .O(N__33371),
            .I(N__33331));
    LocalMux I__7837 (
            .O(N__33368),
            .I(N__33326));
    LocalMux I__7836 (
            .O(N__33365),
            .I(N__33326));
    Span4Mux_h I__7835 (
            .O(N__33362),
            .I(N__33317));
    Span4Mux_s2_h I__7834 (
            .O(N__33359),
            .I(N__33317));
    Span4Mux_h I__7833 (
            .O(N__33352),
            .I(N__33317));
    Span4Mux_s3_v I__7832 (
            .O(N__33347),
            .I(N__33317));
    Span12Mux_s2_h I__7831 (
            .O(N__33344),
            .I(N__33312));
    Span12Mux_s11_h I__7830 (
            .O(N__33337),
            .I(N__33312));
    LocalMux I__7829 (
            .O(N__33334),
            .I(\tok.n289 ));
    LocalMux I__7828 (
            .O(N__33331),
            .I(\tok.n289 ));
    Odrv4 I__7827 (
            .O(N__33326),
            .I(\tok.n289 ));
    Odrv4 I__7826 (
            .O(N__33317),
            .I(\tok.n289 ));
    Odrv12 I__7825 (
            .O(N__33312),
            .I(\tok.n289 ));
    CascadeMux I__7824 (
            .O(N__33301),
            .I(N__33284));
    CascadeMux I__7823 (
            .O(N__33300),
            .I(N__33276));
    CascadeMux I__7822 (
            .O(N__33299),
            .I(N__33260));
    CascadeMux I__7821 (
            .O(N__33298),
            .I(N__33254));
    CascadeMux I__7820 (
            .O(N__33297),
            .I(N__33245));
    InMux I__7819 (
            .O(N__33296),
            .I(N__33241));
    InMux I__7818 (
            .O(N__33295),
            .I(N__33237));
    InMux I__7817 (
            .O(N__33294),
            .I(N__33229));
    InMux I__7816 (
            .O(N__33293),
            .I(N__33224));
    InMux I__7815 (
            .O(N__33292),
            .I(N__33224));
    InMux I__7814 (
            .O(N__33291),
            .I(N__33220));
    InMux I__7813 (
            .O(N__33290),
            .I(N__33212));
    InMux I__7812 (
            .O(N__33289),
            .I(N__33212));
    InMux I__7811 (
            .O(N__33288),
            .I(N__33209));
    InMux I__7810 (
            .O(N__33287),
            .I(N__33206));
    InMux I__7809 (
            .O(N__33284),
            .I(N__33199));
    InMux I__7808 (
            .O(N__33283),
            .I(N__33199));
    InMux I__7807 (
            .O(N__33282),
            .I(N__33199));
    CascadeMux I__7806 (
            .O(N__33281),
            .I(N__33193));
    InMux I__7805 (
            .O(N__33280),
            .I(N__33187));
    InMux I__7804 (
            .O(N__33279),
            .I(N__33176));
    InMux I__7803 (
            .O(N__33276),
            .I(N__33176));
    InMux I__7802 (
            .O(N__33275),
            .I(N__33176));
    InMux I__7801 (
            .O(N__33274),
            .I(N__33169));
    InMux I__7800 (
            .O(N__33273),
            .I(N__33169));
    InMux I__7799 (
            .O(N__33272),
            .I(N__33169));
    InMux I__7798 (
            .O(N__33271),
            .I(N__33154));
    InMux I__7797 (
            .O(N__33270),
            .I(N__33154));
    InMux I__7796 (
            .O(N__33269),
            .I(N__33154));
    InMux I__7795 (
            .O(N__33268),
            .I(N__33151));
    InMux I__7794 (
            .O(N__33267),
            .I(N__33148));
    InMux I__7793 (
            .O(N__33266),
            .I(N__33143));
    InMux I__7792 (
            .O(N__33265),
            .I(N__33143));
    InMux I__7791 (
            .O(N__33264),
            .I(N__33138));
    InMux I__7790 (
            .O(N__33263),
            .I(N__33138));
    InMux I__7789 (
            .O(N__33260),
            .I(N__33130));
    InMux I__7788 (
            .O(N__33259),
            .I(N__33130));
    InMux I__7787 (
            .O(N__33258),
            .I(N__33125));
    InMux I__7786 (
            .O(N__33257),
            .I(N__33125));
    InMux I__7785 (
            .O(N__33254),
            .I(N__33117));
    InMux I__7784 (
            .O(N__33253),
            .I(N__33117));
    InMux I__7783 (
            .O(N__33252),
            .I(N__33117));
    InMux I__7782 (
            .O(N__33251),
            .I(N__33110));
    InMux I__7781 (
            .O(N__33250),
            .I(N__33110));
    InMux I__7780 (
            .O(N__33249),
            .I(N__33110));
    InMux I__7779 (
            .O(N__33248),
            .I(N__33103));
    InMux I__7778 (
            .O(N__33245),
            .I(N__33103));
    InMux I__7777 (
            .O(N__33244),
            .I(N__33103));
    LocalMux I__7776 (
            .O(N__33241),
            .I(N__33094));
    InMux I__7775 (
            .O(N__33240),
            .I(N__33090));
    LocalMux I__7774 (
            .O(N__33237),
            .I(N__33087));
    InMux I__7773 (
            .O(N__33236),
            .I(N__33084));
    InMux I__7772 (
            .O(N__33235),
            .I(N__33079));
    InMux I__7771 (
            .O(N__33234),
            .I(N__33079));
    InMux I__7770 (
            .O(N__33233),
            .I(N__33074));
    InMux I__7769 (
            .O(N__33232),
            .I(N__33074));
    LocalMux I__7768 (
            .O(N__33229),
            .I(N__33069));
    LocalMux I__7767 (
            .O(N__33224),
            .I(N__33069));
    CascadeMux I__7766 (
            .O(N__33223),
            .I(N__33066));
    LocalMux I__7765 (
            .O(N__33220),
            .I(N__33061));
    InMux I__7764 (
            .O(N__33219),
            .I(N__33056));
    InMux I__7763 (
            .O(N__33218),
            .I(N__33056));
    InMux I__7762 (
            .O(N__33217),
            .I(N__33053));
    LocalMux I__7761 (
            .O(N__33212),
            .I(N__33044));
    LocalMux I__7760 (
            .O(N__33209),
            .I(N__33044));
    LocalMux I__7759 (
            .O(N__33206),
            .I(N__33044));
    LocalMux I__7758 (
            .O(N__33199),
            .I(N__33044));
    InMux I__7757 (
            .O(N__33198),
            .I(N__33041));
    InMux I__7756 (
            .O(N__33197),
            .I(N__33032));
    InMux I__7755 (
            .O(N__33196),
            .I(N__33032));
    InMux I__7754 (
            .O(N__33193),
            .I(N__33032));
    InMux I__7753 (
            .O(N__33192),
            .I(N__33032));
    InMux I__7752 (
            .O(N__33191),
            .I(N__33026));
    InMux I__7751 (
            .O(N__33190),
            .I(N__33026));
    LocalMux I__7750 (
            .O(N__33187),
            .I(N__33023));
    InMux I__7749 (
            .O(N__33186),
            .I(N__33015));
    InMux I__7748 (
            .O(N__33185),
            .I(N__33015));
    InMux I__7747 (
            .O(N__33184),
            .I(N__33015));
    InMux I__7746 (
            .O(N__33183),
            .I(N__33012));
    LocalMux I__7745 (
            .O(N__33176),
            .I(N__33007));
    LocalMux I__7744 (
            .O(N__33169),
            .I(N__33007));
    InMux I__7743 (
            .O(N__33168),
            .I(N__33000));
    InMux I__7742 (
            .O(N__33167),
            .I(N__33000));
    InMux I__7741 (
            .O(N__33166),
            .I(N__33000));
    InMux I__7740 (
            .O(N__33165),
            .I(N__32995));
    InMux I__7739 (
            .O(N__33164),
            .I(N__32995));
    CascadeMux I__7738 (
            .O(N__33163),
            .I(N__32992));
    InMux I__7737 (
            .O(N__33162),
            .I(N__32989));
    InMux I__7736 (
            .O(N__33161),
            .I(N__32986));
    LocalMux I__7735 (
            .O(N__33154),
            .I(N__32983));
    LocalMux I__7734 (
            .O(N__33151),
            .I(N__32978));
    LocalMux I__7733 (
            .O(N__33148),
            .I(N__32978));
    LocalMux I__7732 (
            .O(N__33143),
            .I(N__32973));
    LocalMux I__7731 (
            .O(N__33138),
            .I(N__32973));
    InMux I__7730 (
            .O(N__33137),
            .I(N__32968));
    InMux I__7729 (
            .O(N__33136),
            .I(N__32968));
    CascadeMux I__7728 (
            .O(N__33135),
            .I(N__32962));
    LocalMux I__7727 (
            .O(N__33130),
            .I(N__32950));
    LocalMux I__7726 (
            .O(N__33125),
            .I(N__32950));
    InMux I__7725 (
            .O(N__33124),
            .I(N__32947));
    LocalMux I__7724 (
            .O(N__33117),
            .I(N__32944));
    LocalMux I__7723 (
            .O(N__33110),
            .I(N__32941));
    LocalMux I__7722 (
            .O(N__33103),
            .I(N__32938));
    InMux I__7721 (
            .O(N__33102),
            .I(N__32935));
    InMux I__7720 (
            .O(N__33101),
            .I(N__32932));
    InMux I__7719 (
            .O(N__33100),
            .I(N__32929));
    InMux I__7718 (
            .O(N__33099),
            .I(N__32926));
    InMux I__7717 (
            .O(N__33098),
            .I(N__32923));
    InMux I__7716 (
            .O(N__33097),
            .I(N__32920));
    Span4Mux_s3_v I__7715 (
            .O(N__33094),
            .I(N__32917));
    InMux I__7714 (
            .O(N__33093),
            .I(N__32914));
    LocalMux I__7713 (
            .O(N__33090),
            .I(N__32907));
    Span4Mux_s3_v I__7712 (
            .O(N__33087),
            .I(N__32907));
    LocalMux I__7711 (
            .O(N__33084),
            .I(N__32907));
    LocalMux I__7710 (
            .O(N__33079),
            .I(N__32904));
    LocalMux I__7709 (
            .O(N__33074),
            .I(N__32899));
    Span4Mux_v I__7708 (
            .O(N__33069),
            .I(N__32899));
    InMux I__7707 (
            .O(N__33066),
            .I(N__32892));
    InMux I__7706 (
            .O(N__33065),
            .I(N__32892));
    InMux I__7705 (
            .O(N__33064),
            .I(N__32892));
    Span4Mux_v I__7704 (
            .O(N__33061),
            .I(N__32887));
    LocalMux I__7703 (
            .O(N__33056),
            .I(N__32887));
    LocalMux I__7702 (
            .O(N__33053),
            .I(N__32878));
    Span4Mux_v I__7701 (
            .O(N__33044),
            .I(N__32878));
    LocalMux I__7700 (
            .O(N__33041),
            .I(N__32878));
    LocalMux I__7699 (
            .O(N__33032),
            .I(N__32878));
    InMux I__7698 (
            .O(N__33031),
            .I(N__32874));
    LocalMux I__7697 (
            .O(N__33026),
            .I(N__32869));
    Span4Mux_v I__7696 (
            .O(N__33023),
            .I(N__32869));
    InMux I__7695 (
            .O(N__33022),
            .I(N__32866));
    LocalMux I__7694 (
            .O(N__33015),
            .I(N__32857));
    LocalMux I__7693 (
            .O(N__33012),
            .I(N__32857));
    Span4Mux_s3_v I__7692 (
            .O(N__33007),
            .I(N__32857));
    LocalMux I__7691 (
            .O(N__33000),
            .I(N__32857));
    LocalMux I__7690 (
            .O(N__32995),
            .I(N__32854));
    InMux I__7689 (
            .O(N__32992),
            .I(N__32848));
    LocalMux I__7688 (
            .O(N__32989),
            .I(N__32845));
    LocalMux I__7687 (
            .O(N__32986),
            .I(N__32842));
    Span4Mux_v I__7686 (
            .O(N__32983),
            .I(N__32833));
    Span4Mux_s3_v I__7685 (
            .O(N__32978),
            .I(N__32833));
    Span4Mux_h I__7684 (
            .O(N__32973),
            .I(N__32833));
    LocalMux I__7683 (
            .O(N__32968),
            .I(N__32833));
    InMux I__7682 (
            .O(N__32967),
            .I(N__32828));
    InMux I__7681 (
            .O(N__32966),
            .I(N__32828));
    InMux I__7680 (
            .O(N__32965),
            .I(N__32824));
    InMux I__7679 (
            .O(N__32962),
            .I(N__32821));
    InMux I__7678 (
            .O(N__32961),
            .I(N__32816));
    InMux I__7677 (
            .O(N__32960),
            .I(N__32816));
    InMux I__7676 (
            .O(N__32959),
            .I(N__32811));
    InMux I__7675 (
            .O(N__32958),
            .I(N__32811));
    InMux I__7674 (
            .O(N__32957),
            .I(N__32804));
    InMux I__7673 (
            .O(N__32956),
            .I(N__32804));
    InMux I__7672 (
            .O(N__32955),
            .I(N__32804));
    Span4Mux_v I__7671 (
            .O(N__32950),
            .I(N__32799));
    LocalMux I__7670 (
            .O(N__32947),
            .I(N__32799));
    Span4Mux_v I__7669 (
            .O(N__32944),
            .I(N__32790));
    Span4Mux_v I__7668 (
            .O(N__32941),
            .I(N__32790));
    Span4Mux_s2_h I__7667 (
            .O(N__32938),
            .I(N__32790));
    LocalMux I__7666 (
            .O(N__32935),
            .I(N__32790));
    LocalMux I__7665 (
            .O(N__32932),
            .I(N__32782));
    LocalMux I__7664 (
            .O(N__32929),
            .I(N__32775));
    LocalMux I__7663 (
            .O(N__32926),
            .I(N__32766));
    LocalMux I__7662 (
            .O(N__32923),
            .I(N__32766));
    LocalMux I__7661 (
            .O(N__32920),
            .I(N__32766));
    Span4Mux_v I__7660 (
            .O(N__32917),
            .I(N__32766));
    LocalMux I__7659 (
            .O(N__32914),
            .I(N__32761));
    Span4Mux_v I__7658 (
            .O(N__32907),
            .I(N__32761));
    Span4Mux_v I__7657 (
            .O(N__32904),
            .I(N__32750));
    Span4Mux_h I__7656 (
            .O(N__32899),
            .I(N__32750));
    LocalMux I__7655 (
            .O(N__32892),
            .I(N__32750));
    Span4Mux_s2_v I__7654 (
            .O(N__32887),
            .I(N__32750));
    Span4Mux_v I__7653 (
            .O(N__32878),
            .I(N__32750));
    InMux I__7652 (
            .O(N__32877),
            .I(N__32747));
    LocalMux I__7651 (
            .O(N__32874),
            .I(N__32736));
    Span4Mux_h I__7650 (
            .O(N__32869),
            .I(N__32736));
    LocalMux I__7649 (
            .O(N__32866),
            .I(N__32736));
    Span4Mux_v I__7648 (
            .O(N__32857),
            .I(N__32736));
    Span4Mux_v I__7647 (
            .O(N__32854),
            .I(N__32736));
    InMux I__7646 (
            .O(N__32853),
            .I(N__32731));
    InMux I__7645 (
            .O(N__32852),
            .I(N__32731));
    InMux I__7644 (
            .O(N__32851),
            .I(N__32728));
    LocalMux I__7643 (
            .O(N__32848),
            .I(N__32717));
    Span4Mux_h I__7642 (
            .O(N__32845),
            .I(N__32717));
    Span4Mux_s3_h I__7641 (
            .O(N__32842),
            .I(N__32717));
    Span4Mux_h I__7640 (
            .O(N__32833),
            .I(N__32717));
    LocalMux I__7639 (
            .O(N__32828),
            .I(N__32717));
    InMux I__7638 (
            .O(N__32827),
            .I(N__32714));
    LocalMux I__7637 (
            .O(N__32824),
            .I(N__32711));
    LocalMux I__7636 (
            .O(N__32821),
            .I(N__32708));
    LocalMux I__7635 (
            .O(N__32816),
            .I(N__32701));
    LocalMux I__7634 (
            .O(N__32811),
            .I(N__32701));
    LocalMux I__7633 (
            .O(N__32804),
            .I(N__32701));
    Span4Mux_s2_v I__7632 (
            .O(N__32799),
            .I(N__32696));
    Span4Mux_v I__7631 (
            .O(N__32790),
            .I(N__32696));
    InMux I__7630 (
            .O(N__32789),
            .I(N__32691));
    InMux I__7629 (
            .O(N__32788),
            .I(N__32686));
    InMux I__7628 (
            .O(N__32787),
            .I(N__32686));
    InMux I__7627 (
            .O(N__32786),
            .I(N__32683));
    InMux I__7626 (
            .O(N__32785),
            .I(N__32680));
    Span12Mux_s11_v I__7625 (
            .O(N__32782),
            .I(N__32677));
    InMux I__7624 (
            .O(N__32781),
            .I(N__32674));
    InMux I__7623 (
            .O(N__32780),
            .I(N__32667));
    InMux I__7622 (
            .O(N__32779),
            .I(N__32667));
    InMux I__7621 (
            .O(N__32778),
            .I(N__32667));
    Span4Mux_s2_v I__7620 (
            .O(N__32775),
            .I(N__32658));
    Span4Mux_v I__7619 (
            .O(N__32766),
            .I(N__32658));
    Span4Mux_v I__7618 (
            .O(N__32761),
            .I(N__32658));
    Span4Mux_h I__7617 (
            .O(N__32750),
            .I(N__32658));
    LocalMux I__7616 (
            .O(N__32747),
            .I(N__32651));
    Span4Mux_h I__7615 (
            .O(N__32736),
            .I(N__32651));
    LocalMux I__7614 (
            .O(N__32731),
            .I(N__32651));
    LocalMux I__7613 (
            .O(N__32728),
            .I(N__32644));
    Span4Mux_v I__7612 (
            .O(N__32717),
            .I(N__32644));
    LocalMux I__7611 (
            .O(N__32714),
            .I(N__32644));
    Span4Mux_s2_v I__7610 (
            .O(N__32711),
            .I(N__32635));
    Span4Mux_s2_v I__7609 (
            .O(N__32708),
            .I(N__32635));
    Span4Mux_v I__7608 (
            .O(N__32701),
            .I(N__32635));
    Span4Mux_h I__7607 (
            .O(N__32696),
            .I(N__32635));
    InMux I__7606 (
            .O(N__32695),
            .I(N__32630));
    InMux I__7605 (
            .O(N__32694),
            .I(N__32630));
    LocalMux I__7604 (
            .O(N__32691),
            .I(\tok.T_1 ));
    LocalMux I__7603 (
            .O(N__32686),
            .I(\tok.T_1 ));
    LocalMux I__7602 (
            .O(N__32683),
            .I(\tok.T_1 ));
    LocalMux I__7601 (
            .O(N__32680),
            .I(\tok.T_1 ));
    Odrv12 I__7600 (
            .O(N__32677),
            .I(\tok.T_1 ));
    LocalMux I__7599 (
            .O(N__32674),
            .I(\tok.T_1 ));
    LocalMux I__7598 (
            .O(N__32667),
            .I(\tok.T_1 ));
    Odrv4 I__7597 (
            .O(N__32658),
            .I(\tok.T_1 ));
    Odrv4 I__7596 (
            .O(N__32651),
            .I(\tok.T_1 ));
    Odrv4 I__7595 (
            .O(N__32644),
            .I(\tok.T_1 ));
    Odrv4 I__7594 (
            .O(N__32635),
            .I(\tok.T_1 ));
    LocalMux I__7593 (
            .O(N__32630),
            .I(\tok.T_1 ));
    CascadeMux I__7592 (
            .O(N__32605),
            .I(N__32602));
    InMux I__7591 (
            .O(N__32602),
            .I(N__32598));
    InMux I__7590 (
            .O(N__32601),
            .I(N__32595));
    LocalMux I__7589 (
            .O(N__32598),
            .I(N__32590));
    LocalMux I__7588 (
            .O(N__32595),
            .I(N__32587));
    CascadeMux I__7587 (
            .O(N__32594),
            .I(N__32582));
    CascadeMux I__7586 (
            .O(N__32593),
            .I(N__32578));
    Span4Mux_h I__7585 (
            .O(N__32590),
            .I(N__32573));
    Span4Mux_h I__7584 (
            .O(N__32587),
            .I(N__32573));
    InMux I__7583 (
            .O(N__32586),
            .I(N__32570));
    InMux I__7582 (
            .O(N__32585),
            .I(N__32565));
    InMux I__7581 (
            .O(N__32582),
            .I(N__32565));
    InMux I__7580 (
            .O(N__32581),
            .I(N__32560));
    InMux I__7579 (
            .O(N__32578),
            .I(N__32560));
    Odrv4 I__7578 (
            .O(N__32573),
            .I(\tok.n222 ));
    LocalMux I__7577 (
            .O(N__32570),
            .I(\tok.n222 ));
    LocalMux I__7576 (
            .O(N__32565),
            .I(\tok.n222 ));
    LocalMux I__7575 (
            .O(N__32560),
            .I(\tok.n222 ));
    InMux I__7574 (
            .O(N__32551),
            .I(N__32544));
    InMux I__7573 (
            .O(N__32550),
            .I(N__32541));
    InMux I__7572 (
            .O(N__32549),
            .I(N__32538));
    InMux I__7571 (
            .O(N__32548),
            .I(N__32535));
    InMux I__7570 (
            .O(N__32547),
            .I(N__32532));
    LocalMux I__7569 (
            .O(N__32544),
            .I(N__32529));
    LocalMux I__7568 (
            .O(N__32541),
            .I(N__32526));
    LocalMux I__7567 (
            .O(N__32538),
            .I(N__32523));
    LocalMux I__7566 (
            .O(N__32535),
            .I(N__32520));
    LocalMux I__7565 (
            .O(N__32532),
            .I(N__32517));
    Span4Mux_v I__7564 (
            .O(N__32529),
            .I(N__32514));
    Span4Mux_v I__7563 (
            .O(N__32526),
            .I(N__32509));
    Span4Mux_v I__7562 (
            .O(N__32523),
            .I(N__32509));
    Span4Mux_s2_h I__7561 (
            .O(N__32520),
            .I(N__32506));
    Span4Mux_v I__7560 (
            .O(N__32517),
            .I(N__32503));
    Span4Mux_v I__7559 (
            .O(N__32514),
            .I(N__32498));
    Span4Mux_h I__7558 (
            .O(N__32509),
            .I(N__32498));
    Span4Mux_h I__7557 (
            .O(N__32506),
            .I(N__32495));
    Span4Mux_h I__7556 (
            .O(N__32503),
            .I(N__32492));
    Odrv4 I__7555 (
            .O(N__32498),
            .I(\tok.n838 ));
    Odrv4 I__7554 (
            .O(N__32495),
            .I(\tok.n838 ));
    Odrv4 I__7553 (
            .O(N__32492),
            .I(\tok.n838 ));
    CascadeMux I__7552 (
            .O(N__32485),
            .I(\tok.n863_cascade_ ));
    InMux I__7551 (
            .O(N__32482),
            .I(N__32479));
    LocalMux I__7550 (
            .O(N__32479),
            .I(\tok.n6472 ));
    InMux I__7549 (
            .O(N__32476),
            .I(N__32473));
    LocalMux I__7548 (
            .O(N__32473),
            .I(N__32466));
    InMux I__7547 (
            .O(N__32472),
            .I(N__32461));
    InMux I__7546 (
            .O(N__32471),
            .I(N__32461));
    InMux I__7545 (
            .O(N__32470),
            .I(N__32457));
    InMux I__7544 (
            .O(N__32469),
            .I(N__32454));
    Span4Mux_v I__7543 (
            .O(N__32466),
            .I(N__32449));
    LocalMux I__7542 (
            .O(N__32461),
            .I(N__32449));
    InMux I__7541 (
            .O(N__32460),
            .I(N__32446));
    LocalMux I__7540 (
            .O(N__32457),
            .I(N__32443));
    LocalMux I__7539 (
            .O(N__32454),
            .I(N__32438));
    Span4Mux_v I__7538 (
            .O(N__32449),
            .I(N__32438));
    LocalMux I__7537 (
            .O(N__32446),
            .I(N__32435));
    Span4Mux_h I__7536 (
            .O(N__32443),
            .I(N__32426));
    Span4Mux_h I__7535 (
            .O(N__32438),
            .I(N__32426));
    Span4Mux_v I__7534 (
            .O(N__32435),
            .I(N__32426));
    InMux I__7533 (
            .O(N__32434),
            .I(N__32421));
    InMux I__7532 (
            .O(N__32433),
            .I(N__32421));
    Span4Mux_h I__7531 (
            .O(N__32426),
            .I(N__32418));
    LocalMux I__7530 (
            .O(N__32421),
            .I(N__32415));
    Span4Mux_h I__7529 (
            .O(N__32418),
            .I(N__32412));
    Odrv12 I__7528 (
            .O(N__32415),
            .I(\tok.n9_adj_677 ));
    Odrv4 I__7527 (
            .O(N__32412),
            .I(\tok.n9_adj_677 ));
    InMux I__7526 (
            .O(N__32407),
            .I(N__32404));
    LocalMux I__7525 (
            .O(N__32404),
            .I(N__32401));
    Span4Mux_v I__7524 (
            .O(N__32401),
            .I(N__32397));
    InMux I__7523 (
            .O(N__32400),
            .I(N__32394));
    Span4Mux_h I__7522 (
            .O(N__32397),
            .I(N__32391));
    LocalMux I__7521 (
            .O(N__32394),
            .I(\tok.n205 ));
    Odrv4 I__7520 (
            .O(N__32391),
            .I(\tok.n205 ));
    InMux I__7519 (
            .O(N__32386),
            .I(N__32383));
    LocalMux I__7518 (
            .O(N__32383),
            .I(\tok.n6477 ));
    InMux I__7517 (
            .O(N__32380),
            .I(N__32374));
    InMux I__7516 (
            .O(N__32379),
            .I(N__32369));
    InMux I__7515 (
            .O(N__32378),
            .I(N__32363));
    InMux I__7514 (
            .O(N__32377),
            .I(N__32363));
    LocalMux I__7513 (
            .O(N__32374),
            .I(N__32360));
    CascadeMux I__7512 (
            .O(N__32373),
            .I(N__32357));
    InMux I__7511 (
            .O(N__32372),
            .I(N__32351));
    LocalMux I__7510 (
            .O(N__32369),
            .I(N__32348));
    InMux I__7509 (
            .O(N__32368),
            .I(N__32345));
    LocalMux I__7508 (
            .O(N__32363),
            .I(N__32342));
    Span4Mux_s3_v I__7507 (
            .O(N__32360),
            .I(N__32339));
    InMux I__7506 (
            .O(N__32357),
            .I(N__32336));
    InMux I__7505 (
            .O(N__32356),
            .I(N__32331));
    InMux I__7504 (
            .O(N__32355),
            .I(N__32331));
    InMux I__7503 (
            .O(N__32354),
            .I(N__32327));
    LocalMux I__7502 (
            .O(N__32351),
            .I(N__32324));
    Span4Mux_v I__7501 (
            .O(N__32348),
            .I(N__32319));
    LocalMux I__7500 (
            .O(N__32345),
            .I(N__32319));
    Span4Mux_v I__7499 (
            .O(N__32342),
            .I(N__32316));
    Span4Mux_v I__7498 (
            .O(N__32339),
            .I(N__32313));
    LocalMux I__7497 (
            .O(N__32336),
            .I(N__32308));
    LocalMux I__7496 (
            .O(N__32331),
            .I(N__32308));
    InMux I__7495 (
            .O(N__32330),
            .I(N__32305));
    LocalMux I__7494 (
            .O(N__32327),
            .I(N__32302));
    Span4Mux_v I__7493 (
            .O(N__32324),
            .I(N__32295));
    Span4Mux_v I__7492 (
            .O(N__32319),
            .I(N__32295));
    Span4Mux_h I__7491 (
            .O(N__32316),
            .I(N__32295));
    Span4Mux_h I__7490 (
            .O(N__32313),
            .I(N__32290));
    Span4Mux_h I__7489 (
            .O(N__32308),
            .I(N__32290));
    LocalMux I__7488 (
            .O(N__32305),
            .I(\tok.n43 ));
    Odrv4 I__7487 (
            .O(N__32302),
            .I(\tok.n43 ));
    Odrv4 I__7486 (
            .O(N__32295),
            .I(\tok.n43 ));
    Odrv4 I__7485 (
            .O(N__32290),
            .I(\tok.n43 ));
    InMux I__7484 (
            .O(N__32281),
            .I(N__32278));
    LocalMux I__7483 (
            .O(N__32278),
            .I(N__32275));
    Span4Mux_h I__7482 (
            .O(N__32275),
            .I(N__32271));
    CascadeMux I__7481 (
            .O(N__32274),
            .I(N__32268));
    Span4Mux_h I__7480 (
            .O(N__32271),
            .I(N__32265));
    InMux I__7479 (
            .O(N__32268),
            .I(N__32262));
    Span4Mux_h I__7478 (
            .O(N__32265),
            .I(N__32259));
    LocalMux I__7477 (
            .O(N__32262),
            .I(N__32256));
    Odrv4 I__7476 (
            .O(N__32259),
            .I(\tok.n311 ));
    Odrv12 I__7475 (
            .O(N__32256),
            .I(\tok.n311 ));
    CascadeMux I__7474 (
            .O(N__32251),
            .I(N__32248));
    InMux I__7473 (
            .O(N__32248),
            .I(N__32244));
    InMux I__7472 (
            .O(N__32247),
            .I(N__32241));
    LocalMux I__7471 (
            .O(N__32244),
            .I(N__32236));
    LocalMux I__7470 (
            .O(N__32241),
            .I(N__32236));
    Odrv12 I__7469 (
            .O(N__32236),
            .I(\tok.n190_adj_797 ));
    InMux I__7468 (
            .O(N__32233),
            .I(N__32227));
    InMux I__7467 (
            .O(N__32232),
            .I(N__32224));
    InMux I__7466 (
            .O(N__32231),
            .I(N__32221));
    InMux I__7465 (
            .O(N__32230),
            .I(N__32217));
    LocalMux I__7464 (
            .O(N__32227),
            .I(N__32214));
    LocalMux I__7463 (
            .O(N__32224),
            .I(N__32211));
    LocalMux I__7462 (
            .O(N__32221),
            .I(N__32207));
    InMux I__7461 (
            .O(N__32220),
            .I(N__32204));
    LocalMux I__7460 (
            .O(N__32217),
            .I(N__32201));
    Span4Mux_h I__7459 (
            .O(N__32214),
            .I(N__32197));
    Span4Mux_v I__7458 (
            .O(N__32211),
            .I(N__32194));
    InMux I__7457 (
            .O(N__32210),
            .I(N__32191));
    Span4Mux_h I__7456 (
            .O(N__32207),
            .I(N__32183));
    LocalMux I__7455 (
            .O(N__32204),
            .I(N__32183));
    Span4Mux_h I__7454 (
            .O(N__32201),
            .I(N__32180));
    InMux I__7453 (
            .O(N__32200),
            .I(N__32177));
    Span4Mux_v I__7452 (
            .O(N__32197),
            .I(N__32170));
    Span4Mux_v I__7451 (
            .O(N__32194),
            .I(N__32170));
    LocalMux I__7450 (
            .O(N__32191),
            .I(N__32170));
    InMux I__7449 (
            .O(N__32190),
            .I(N__32164));
    InMux I__7448 (
            .O(N__32189),
            .I(N__32164));
    InMux I__7447 (
            .O(N__32188),
            .I(N__32161));
    Span4Mux_h I__7446 (
            .O(N__32183),
            .I(N__32154));
    Span4Mux_h I__7445 (
            .O(N__32180),
            .I(N__32154));
    LocalMux I__7444 (
            .O(N__32177),
            .I(N__32154));
    Span4Mux_h I__7443 (
            .O(N__32170),
            .I(N__32151));
    InMux I__7442 (
            .O(N__32169),
            .I(N__32148));
    LocalMux I__7441 (
            .O(N__32164),
            .I(N__32145));
    LocalMux I__7440 (
            .O(N__32161),
            .I(\tok.n44 ));
    Odrv4 I__7439 (
            .O(N__32154),
            .I(\tok.n44 ));
    Odrv4 I__7438 (
            .O(N__32151),
            .I(\tok.n44 ));
    LocalMux I__7437 (
            .O(N__32148),
            .I(\tok.n44 ));
    Odrv12 I__7436 (
            .O(N__32145),
            .I(\tok.n44 ));
    CascadeMux I__7435 (
            .O(N__32134),
            .I(N__32128));
    InMux I__7434 (
            .O(N__32133),
            .I(N__32101));
    InMux I__7433 (
            .O(N__32132),
            .I(N__32101));
    CascadeMux I__7432 (
            .O(N__32131),
            .I(N__32088));
    InMux I__7431 (
            .O(N__32128),
            .I(N__32084));
    InMux I__7430 (
            .O(N__32127),
            .I(N__32081));
    CascadeMux I__7429 (
            .O(N__32126),
            .I(N__32072));
    InMux I__7428 (
            .O(N__32125),
            .I(N__32066));
    InMux I__7427 (
            .O(N__32124),
            .I(N__32066));
    InMux I__7426 (
            .O(N__32123),
            .I(N__32060));
    InMux I__7425 (
            .O(N__32122),
            .I(N__32056));
    InMux I__7424 (
            .O(N__32121),
            .I(N__32053));
    InMux I__7423 (
            .O(N__32120),
            .I(N__32046));
    InMux I__7422 (
            .O(N__32119),
            .I(N__32046));
    InMux I__7421 (
            .O(N__32118),
            .I(N__32046));
    CascadeMux I__7420 (
            .O(N__32117),
            .I(N__32038));
    CascadeMux I__7419 (
            .O(N__32116),
            .I(N__32035));
    InMux I__7418 (
            .O(N__32115),
            .I(N__32030));
    InMux I__7417 (
            .O(N__32114),
            .I(N__32025));
    InMux I__7416 (
            .O(N__32113),
            .I(N__32025));
    CascadeMux I__7415 (
            .O(N__32112),
            .I(N__32015));
    InMux I__7414 (
            .O(N__32111),
            .I(N__32012));
    InMux I__7413 (
            .O(N__32110),
            .I(N__32005));
    InMux I__7412 (
            .O(N__32109),
            .I(N__32005));
    InMux I__7411 (
            .O(N__32108),
            .I(N__32005));
    InMux I__7410 (
            .O(N__32107),
            .I(N__32002));
    InMux I__7409 (
            .O(N__32106),
            .I(N__31999));
    LocalMux I__7408 (
            .O(N__32101),
            .I(N__31996));
    InMux I__7407 (
            .O(N__32100),
            .I(N__31989));
    InMux I__7406 (
            .O(N__32099),
            .I(N__31989));
    InMux I__7405 (
            .O(N__32098),
            .I(N__31989));
    InMux I__7404 (
            .O(N__32097),
            .I(N__31982));
    InMux I__7403 (
            .O(N__32096),
            .I(N__31982));
    InMux I__7402 (
            .O(N__32095),
            .I(N__31982));
    CascadeMux I__7401 (
            .O(N__32094),
            .I(N__31975));
    InMux I__7400 (
            .O(N__32093),
            .I(N__31968));
    InMux I__7399 (
            .O(N__32092),
            .I(N__31968));
    InMux I__7398 (
            .O(N__32091),
            .I(N__31961));
    InMux I__7397 (
            .O(N__32088),
            .I(N__31961));
    InMux I__7396 (
            .O(N__32087),
            .I(N__31961));
    LocalMux I__7395 (
            .O(N__32084),
            .I(N__31950));
    LocalMux I__7394 (
            .O(N__32081),
            .I(N__31950));
    InMux I__7393 (
            .O(N__32080),
            .I(N__31945));
    InMux I__7392 (
            .O(N__32079),
            .I(N__31945));
    InMux I__7391 (
            .O(N__32078),
            .I(N__31928));
    InMux I__7390 (
            .O(N__32077),
            .I(N__31923));
    InMux I__7389 (
            .O(N__32076),
            .I(N__31923));
    CascadeMux I__7388 (
            .O(N__32075),
            .I(N__31909));
    InMux I__7387 (
            .O(N__32072),
            .I(N__31902));
    InMux I__7386 (
            .O(N__32071),
            .I(N__31899));
    LocalMux I__7385 (
            .O(N__32066),
            .I(N__31893));
    InMux I__7384 (
            .O(N__32065),
            .I(N__31886));
    InMux I__7383 (
            .O(N__32064),
            .I(N__31886));
    InMux I__7382 (
            .O(N__32063),
            .I(N__31886));
    LocalMux I__7381 (
            .O(N__32060),
            .I(N__31881));
    InMux I__7380 (
            .O(N__32059),
            .I(N__31872));
    LocalMux I__7379 (
            .O(N__32056),
            .I(N__31865));
    LocalMux I__7378 (
            .O(N__32053),
            .I(N__31865));
    LocalMux I__7377 (
            .O(N__32046),
            .I(N__31865));
    InMux I__7376 (
            .O(N__32045),
            .I(N__31858));
    InMux I__7375 (
            .O(N__32044),
            .I(N__31858));
    InMux I__7374 (
            .O(N__32043),
            .I(N__31858));
    InMux I__7373 (
            .O(N__32042),
            .I(N__31855));
    InMux I__7372 (
            .O(N__32041),
            .I(N__31844));
    InMux I__7371 (
            .O(N__32038),
            .I(N__31844));
    InMux I__7370 (
            .O(N__32035),
            .I(N__31844));
    InMux I__7369 (
            .O(N__32034),
            .I(N__31844));
    InMux I__7368 (
            .O(N__32033),
            .I(N__31844));
    LocalMux I__7367 (
            .O(N__32030),
            .I(N__31839));
    LocalMux I__7366 (
            .O(N__32025),
            .I(N__31839));
    InMux I__7365 (
            .O(N__32024),
            .I(N__31834));
    InMux I__7364 (
            .O(N__32023),
            .I(N__31834));
    InMux I__7363 (
            .O(N__32022),
            .I(N__31829));
    InMux I__7362 (
            .O(N__32021),
            .I(N__31829));
    InMux I__7361 (
            .O(N__32020),
            .I(N__31823));
    InMux I__7360 (
            .O(N__32019),
            .I(N__31818));
    InMux I__7359 (
            .O(N__32018),
            .I(N__31818));
    InMux I__7358 (
            .O(N__32015),
            .I(N__31815));
    LocalMux I__7357 (
            .O(N__32012),
            .I(N__31810));
    LocalMux I__7356 (
            .O(N__32005),
            .I(N__31810));
    LocalMux I__7355 (
            .O(N__32002),
            .I(N__31801));
    LocalMux I__7354 (
            .O(N__31999),
            .I(N__31801));
    Span4Mux_s2_h I__7353 (
            .O(N__31996),
            .I(N__31801));
    LocalMux I__7352 (
            .O(N__31989),
            .I(N__31801));
    LocalMux I__7351 (
            .O(N__31982),
            .I(N__31798));
    InMux I__7350 (
            .O(N__31981),
            .I(N__31789));
    InMux I__7349 (
            .O(N__31980),
            .I(N__31789));
    InMux I__7348 (
            .O(N__31979),
            .I(N__31789));
    InMux I__7347 (
            .O(N__31978),
            .I(N__31789));
    InMux I__7346 (
            .O(N__31975),
            .I(N__31782));
    InMux I__7345 (
            .O(N__31974),
            .I(N__31782));
    InMux I__7344 (
            .O(N__31973),
            .I(N__31782));
    LocalMux I__7343 (
            .O(N__31968),
            .I(N__31779));
    LocalMux I__7342 (
            .O(N__31961),
            .I(N__31776));
    InMux I__7341 (
            .O(N__31960),
            .I(N__31769));
    InMux I__7340 (
            .O(N__31959),
            .I(N__31769));
    InMux I__7339 (
            .O(N__31958),
            .I(N__31769));
    CascadeMux I__7338 (
            .O(N__31957),
            .I(N__31766));
    InMux I__7337 (
            .O(N__31956),
            .I(N__31762));
    InMux I__7336 (
            .O(N__31955),
            .I(N__31759));
    Span4Mux_s2_h I__7335 (
            .O(N__31950),
            .I(N__31756));
    LocalMux I__7334 (
            .O(N__31945),
            .I(N__31753));
    InMux I__7333 (
            .O(N__31944),
            .I(N__31746));
    InMux I__7332 (
            .O(N__31943),
            .I(N__31746));
    InMux I__7331 (
            .O(N__31942),
            .I(N__31746));
    InMux I__7330 (
            .O(N__31941),
            .I(N__31738));
    InMux I__7329 (
            .O(N__31940),
            .I(N__31738));
    InMux I__7328 (
            .O(N__31939),
            .I(N__31735));
    InMux I__7327 (
            .O(N__31938),
            .I(N__31730));
    InMux I__7326 (
            .O(N__31937),
            .I(N__31730));
    InMux I__7325 (
            .O(N__31936),
            .I(N__31725));
    InMux I__7324 (
            .O(N__31935),
            .I(N__31725));
    InMux I__7323 (
            .O(N__31934),
            .I(N__31720));
    InMux I__7322 (
            .O(N__31933),
            .I(N__31720));
    InMux I__7321 (
            .O(N__31932),
            .I(N__31715));
    InMux I__7320 (
            .O(N__31931),
            .I(N__31715));
    LocalMux I__7319 (
            .O(N__31928),
            .I(N__31712));
    LocalMux I__7318 (
            .O(N__31923),
            .I(N__31709));
    InMux I__7317 (
            .O(N__31922),
            .I(N__31704));
    InMux I__7316 (
            .O(N__31921),
            .I(N__31704));
    InMux I__7315 (
            .O(N__31920),
            .I(N__31699));
    InMux I__7314 (
            .O(N__31919),
            .I(N__31699));
    InMux I__7313 (
            .O(N__31918),
            .I(N__31694));
    InMux I__7312 (
            .O(N__31917),
            .I(N__31694));
    InMux I__7311 (
            .O(N__31916),
            .I(N__31691));
    InMux I__7310 (
            .O(N__31915),
            .I(N__31682));
    InMux I__7309 (
            .O(N__31914),
            .I(N__31682));
    InMux I__7308 (
            .O(N__31913),
            .I(N__31682));
    InMux I__7307 (
            .O(N__31912),
            .I(N__31682));
    InMux I__7306 (
            .O(N__31909),
            .I(N__31679));
    InMux I__7305 (
            .O(N__31908),
            .I(N__31676));
    InMux I__7304 (
            .O(N__31907),
            .I(N__31673));
    InMux I__7303 (
            .O(N__31906),
            .I(N__31666));
    InMux I__7302 (
            .O(N__31905),
            .I(N__31666));
    LocalMux I__7301 (
            .O(N__31902),
            .I(N__31661));
    LocalMux I__7300 (
            .O(N__31899),
            .I(N__31661));
    InMux I__7299 (
            .O(N__31898),
            .I(N__31658));
    InMux I__7298 (
            .O(N__31897),
            .I(N__31653));
    InMux I__7297 (
            .O(N__31896),
            .I(N__31653));
    Span4Mux_v I__7296 (
            .O(N__31893),
            .I(N__31650));
    LocalMux I__7295 (
            .O(N__31886),
            .I(N__31647));
    InMux I__7294 (
            .O(N__31885),
            .I(N__31642));
    InMux I__7293 (
            .O(N__31884),
            .I(N__31642));
    Span4Mux_v I__7292 (
            .O(N__31881),
            .I(N__31639));
    InMux I__7291 (
            .O(N__31880),
            .I(N__31634));
    InMux I__7290 (
            .O(N__31879),
            .I(N__31634));
    InMux I__7289 (
            .O(N__31878),
            .I(N__31625));
    InMux I__7288 (
            .O(N__31877),
            .I(N__31625));
    InMux I__7287 (
            .O(N__31876),
            .I(N__31625));
    InMux I__7286 (
            .O(N__31875),
            .I(N__31625));
    LocalMux I__7285 (
            .O(N__31872),
            .I(N__31618));
    Span4Mux_h I__7284 (
            .O(N__31865),
            .I(N__31618));
    LocalMux I__7283 (
            .O(N__31858),
            .I(N__31618));
    LocalMux I__7282 (
            .O(N__31855),
            .I(N__31611));
    LocalMux I__7281 (
            .O(N__31844),
            .I(N__31611));
    Span4Mux_s2_h I__7280 (
            .O(N__31839),
            .I(N__31611));
    LocalMux I__7279 (
            .O(N__31834),
            .I(N__31606));
    LocalMux I__7278 (
            .O(N__31829),
            .I(N__31606));
    InMux I__7277 (
            .O(N__31828),
            .I(N__31601));
    InMux I__7276 (
            .O(N__31827),
            .I(N__31601));
    InMux I__7275 (
            .O(N__31826),
            .I(N__31598));
    LocalMux I__7274 (
            .O(N__31823),
            .I(N__31593));
    LocalMux I__7273 (
            .O(N__31818),
            .I(N__31593));
    LocalMux I__7272 (
            .O(N__31815),
            .I(N__31582));
    Span4Mux_h I__7271 (
            .O(N__31810),
            .I(N__31582));
    Span4Mux_h I__7270 (
            .O(N__31801),
            .I(N__31582));
    Span4Mux_v I__7269 (
            .O(N__31798),
            .I(N__31582));
    LocalMux I__7268 (
            .O(N__31789),
            .I(N__31582));
    LocalMux I__7267 (
            .O(N__31782),
            .I(N__31573));
    Span4Mux_v I__7266 (
            .O(N__31779),
            .I(N__31573));
    Span4Mux_s2_h I__7265 (
            .O(N__31776),
            .I(N__31573));
    LocalMux I__7264 (
            .O(N__31769),
            .I(N__31573));
    InMux I__7263 (
            .O(N__31766),
            .I(N__31569));
    InMux I__7262 (
            .O(N__31765),
            .I(N__31566));
    LocalMux I__7261 (
            .O(N__31762),
            .I(N__31555));
    LocalMux I__7260 (
            .O(N__31759),
            .I(N__31555));
    Span4Mux_v I__7259 (
            .O(N__31756),
            .I(N__31555));
    Span4Mux_s3_v I__7258 (
            .O(N__31753),
            .I(N__31555));
    LocalMux I__7257 (
            .O(N__31746),
            .I(N__31555));
    InMux I__7256 (
            .O(N__31745),
            .I(N__31550));
    InMux I__7255 (
            .O(N__31744),
            .I(N__31550));
    InMux I__7254 (
            .O(N__31743),
            .I(N__31542));
    LocalMux I__7253 (
            .O(N__31738),
            .I(N__31539));
    LocalMux I__7252 (
            .O(N__31735),
            .I(N__31535));
    LocalMux I__7251 (
            .O(N__31730),
            .I(N__31528));
    LocalMux I__7250 (
            .O(N__31725),
            .I(N__31528));
    LocalMux I__7249 (
            .O(N__31720),
            .I(N__31528));
    LocalMux I__7248 (
            .O(N__31715),
            .I(N__31525));
    Span4Mux_s3_h I__7247 (
            .O(N__31712),
            .I(N__31520));
    Span4Mux_v I__7246 (
            .O(N__31709),
            .I(N__31520));
    LocalMux I__7245 (
            .O(N__31704),
            .I(N__31513));
    LocalMux I__7244 (
            .O(N__31699),
            .I(N__31513));
    LocalMux I__7243 (
            .O(N__31694),
            .I(N__31513));
    LocalMux I__7242 (
            .O(N__31691),
            .I(N__31510));
    LocalMux I__7241 (
            .O(N__31682),
            .I(N__31507));
    LocalMux I__7240 (
            .O(N__31679),
            .I(N__31504));
    LocalMux I__7239 (
            .O(N__31676),
            .I(N__31499));
    LocalMux I__7238 (
            .O(N__31673),
            .I(N__31499));
    InMux I__7237 (
            .O(N__31672),
            .I(N__31494));
    InMux I__7236 (
            .O(N__31671),
            .I(N__31494));
    LocalMux I__7235 (
            .O(N__31666),
            .I(N__31487));
    Span4Mux_v I__7234 (
            .O(N__31661),
            .I(N__31487));
    LocalMux I__7233 (
            .O(N__31658),
            .I(N__31487));
    LocalMux I__7232 (
            .O(N__31653),
            .I(N__31476));
    Span4Mux_v I__7231 (
            .O(N__31650),
            .I(N__31476));
    Span4Mux_s2_v I__7230 (
            .O(N__31647),
            .I(N__31476));
    LocalMux I__7229 (
            .O(N__31642),
            .I(N__31476));
    Span4Mux_v I__7228 (
            .O(N__31639),
            .I(N__31476));
    LocalMux I__7227 (
            .O(N__31634),
            .I(N__31471));
    LocalMux I__7226 (
            .O(N__31625),
            .I(N__31471));
    Span4Mux_v I__7225 (
            .O(N__31618),
            .I(N__31463));
    Span4Mux_h I__7224 (
            .O(N__31611),
            .I(N__31463));
    Span4Mux_h I__7223 (
            .O(N__31606),
            .I(N__31458));
    LocalMux I__7222 (
            .O(N__31601),
            .I(N__31458));
    LocalMux I__7221 (
            .O(N__31598),
            .I(N__31455));
    Span4Mux_v I__7220 (
            .O(N__31593),
            .I(N__31448));
    Span4Mux_v I__7219 (
            .O(N__31582),
            .I(N__31448));
    Span4Mux_h I__7218 (
            .O(N__31573),
            .I(N__31448));
    InMux I__7217 (
            .O(N__31572),
            .I(N__31445));
    LocalMux I__7216 (
            .O(N__31569),
            .I(N__31436));
    LocalMux I__7215 (
            .O(N__31566),
            .I(N__31436));
    Sp12to4 I__7214 (
            .O(N__31555),
            .I(N__31436));
    LocalMux I__7213 (
            .O(N__31550),
            .I(N__31436));
    InMux I__7212 (
            .O(N__31549),
            .I(N__31431));
    InMux I__7211 (
            .O(N__31548),
            .I(N__31431));
    InMux I__7210 (
            .O(N__31547),
            .I(N__31428));
    InMux I__7209 (
            .O(N__31546),
            .I(N__31423));
    InMux I__7208 (
            .O(N__31545),
            .I(N__31423));
    LocalMux I__7207 (
            .O(N__31542),
            .I(N__31420));
    Span4Mux_v I__7206 (
            .O(N__31539),
            .I(N__31417));
    InMux I__7205 (
            .O(N__31538),
            .I(N__31414));
    Span12Mux_s3_h I__7204 (
            .O(N__31535),
            .I(N__31409));
    Span12Mux_s10_h I__7203 (
            .O(N__31528),
            .I(N__31409));
    Span4Mux_v I__7202 (
            .O(N__31525),
            .I(N__31398));
    Span4Mux_h I__7201 (
            .O(N__31520),
            .I(N__31398));
    Span4Mux_v I__7200 (
            .O(N__31513),
            .I(N__31398));
    Span4Mux_s2_v I__7199 (
            .O(N__31510),
            .I(N__31398));
    Span4Mux_v I__7198 (
            .O(N__31507),
            .I(N__31398));
    Span4Mux_v I__7197 (
            .O(N__31504),
            .I(N__31389));
    Span4Mux_v I__7196 (
            .O(N__31499),
            .I(N__31389));
    LocalMux I__7195 (
            .O(N__31494),
            .I(N__31389));
    Span4Mux_h I__7194 (
            .O(N__31487),
            .I(N__31389));
    Sp12to4 I__7193 (
            .O(N__31476),
            .I(N__31384));
    Span12Mux_s11_v I__7192 (
            .O(N__31471),
            .I(N__31384));
    InMux I__7191 (
            .O(N__31470),
            .I(N__31377));
    InMux I__7190 (
            .O(N__31469),
            .I(N__31377));
    InMux I__7189 (
            .O(N__31468),
            .I(N__31377));
    Span4Mux_h I__7188 (
            .O(N__31463),
            .I(N__31372));
    Span4Mux_v I__7187 (
            .O(N__31458),
            .I(N__31372));
    Span4Mux_v I__7186 (
            .O(N__31455),
            .I(N__31365));
    Span4Mux_h I__7185 (
            .O(N__31448),
            .I(N__31365));
    LocalMux I__7184 (
            .O(N__31445),
            .I(N__31365));
    Span12Mux_s10_h I__7183 (
            .O(N__31436),
            .I(N__31362));
    LocalMux I__7182 (
            .O(N__31431),
            .I(\tok.T_2 ));
    LocalMux I__7181 (
            .O(N__31428),
            .I(\tok.T_2 ));
    LocalMux I__7180 (
            .O(N__31423),
            .I(\tok.T_2 ));
    Odrv4 I__7179 (
            .O(N__31420),
            .I(\tok.T_2 ));
    Odrv4 I__7178 (
            .O(N__31417),
            .I(\tok.T_2 ));
    LocalMux I__7177 (
            .O(N__31414),
            .I(\tok.T_2 ));
    Odrv12 I__7176 (
            .O(N__31409),
            .I(\tok.T_2 ));
    Odrv4 I__7175 (
            .O(N__31398),
            .I(\tok.T_2 ));
    Odrv4 I__7174 (
            .O(N__31389),
            .I(\tok.T_2 ));
    Odrv12 I__7173 (
            .O(N__31384),
            .I(\tok.T_2 ));
    LocalMux I__7172 (
            .O(N__31377),
            .I(\tok.T_2 ));
    Odrv4 I__7171 (
            .O(N__31372),
            .I(\tok.T_2 ));
    Odrv4 I__7170 (
            .O(N__31365),
            .I(\tok.T_2 ));
    Odrv12 I__7169 (
            .O(N__31362),
            .I(\tok.T_2 ));
    InMux I__7168 (
            .O(N__31333),
            .I(N__31291));
    InMux I__7167 (
            .O(N__31332),
            .I(N__31291));
    InMux I__7166 (
            .O(N__31331),
            .I(N__31286));
    InMux I__7165 (
            .O(N__31330),
            .I(N__31286));
    InMux I__7164 (
            .O(N__31329),
            .I(N__31276));
    InMux I__7163 (
            .O(N__31328),
            .I(N__31276));
    InMux I__7162 (
            .O(N__31327),
            .I(N__31276));
    InMux I__7161 (
            .O(N__31326),
            .I(N__31276));
    InMux I__7160 (
            .O(N__31325),
            .I(N__31271));
    InMux I__7159 (
            .O(N__31324),
            .I(N__31271));
    InMux I__7158 (
            .O(N__31323),
            .I(N__31262));
    InMux I__7157 (
            .O(N__31322),
            .I(N__31262));
    InMux I__7156 (
            .O(N__31321),
            .I(N__31262));
    InMux I__7155 (
            .O(N__31320),
            .I(N__31262));
    InMux I__7154 (
            .O(N__31319),
            .I(N__31253));
    InMux I__7153 (
            .O(N__31318),
            .I(N__31253));
    InMux I__7152 (
            .O(N__31317),
            .I(N__31253));
    InMux I__7151 (
            .O(N__31316),
            .I(N__31253));
    InMux I__7150 (
            .O(N__31315),
            .I(N__31244));
    InMux I__7149 (
            .O(N__31314),
            .I(N__31244));
    InMux I__7148 (
            .O(N__31313),
            .I(N__31241));
    InMux I__7147 (
            .O(N__31312),
            .I(N__31232));
    CascadeMux I__7146 (
            .O(N__31311),
            .I(N__31217));
    InMux I__7145 (
            .O(N__31310),
            .I(N__31203));
    InMux I__7144 (
            .O(N__31309),
            .I(N__31196));
    InMux I__7143 (
            .O(N__31308),
            .I(N__31196));
    InMux I__7142 (
            .O(N__31307),
            .I(N__31196));
    InMux I__7141 (
            .O(N__31306),
            .I(N__31189));
    InMux I__7140 (
            .O(N__31305),
            .I(N__31189));
    InMux I__7139 (
            .O(N__31304),
            .I(N__31189));
    InMux I__7138 (
            .O(N__31303),
            .I(N__31182));
    InMux I__7137 (
            .O(N__31302),
            .I(N__31182));
    InMux I__7136 (
            .O(N__31301),
            .I(N__31175));
    InMux I__7135 (
            .O(N__31300),
            .I(N__31175));
    InMux I__7134 (
            .O(N__31299),
            .I(N__31175));
    InMux I__7133 (
            .O(N__31298),
            .I(N__31168));
    InMux I__7132 (
            .O(N__31297),
            .I(N__31168));
    InMux I__7131 (
            .O(N__31296),
            .I(N__31156));
    LocalMux I__7130 (
            .O(N__31291),
            .I(N__31151));
    LocalMux I__7129 (
            .O(N__31286),
            .I(N__31151));
    InMux I__7128 (
            .O(N__31285),
            .I(N__31148));
    LocalMux I__7127 (
            .O(N__31276),
            .I(N__31145));
    LocalMux I__7126 (
            .O(N__31271),
            .I(N__31138));
    LocalMux I__7125 (
            .O(N__31262),
            .I(N__31138));
    LocalMux I__7124 (
            .O(N__31253),
            .I(N__31138));
    InMux I__7123 (
            .O(N__31252),
            .I(N__31131));
    InMux I__7122 (
            .O(N__31251),
            .I(N__31131));
    InMux I__7121 (
            .O(N__31250),
            .I(N__31131));
    InMux I__7120 (
            .O(N__31249),
            .I(N__31127));
    LocalMux I__7119 (
            .O(N__31244),
            .I(N__31122));
    LocalMux I__7118 (
            .O(N__31241),
            .I(N__31122));
    InMux I__7117 (
            .O(N__31240),
            .I(N__31113));
    InMux I__7116 (
            .O(N__31239),
            .I(N__31113));
    InMux I__7115 (
            .O(N__31238),
            .I(N__31113));
    InMux I__7114 (
            .O(N__31237),
            .I(N__31113));
    InMux I__7113 (
            .O(N__31236),
            .I(N__31105));
    InMux I__7112 (
            .O(N__31235),
            .I(N__31105));
    LocalMux I__7111 (
            .O(N__31232),
            .I(N__31102));
    InMux I__7110 (
            .O(N__31231),
            .I(N__31097));
    InMux I__7109 (
            .O(N__31230),
            .I(N__31097));
    InMux I__7108 (
            .O(N__31229),
            .I(N__31083));
    InMux I__7107 (
            .O(N__31228),
            .I(N__31080));
    InMux I__7106 (
            .O(N__31227),
            .I(N__31073));
    InMux I__7105 (
            .O(N__31226),
            .I(N__31073));
    InMux I__7104 (
            .O(N__31225),
            .I(N__31073));
    InMux I__7103 (
            .O(N__31224),
            .I(N__31065));
    InMux I__7102 (
            .O(N__31223),
            .I(N__31058));
    InMux I__7101 (
            .O(N__31222),
            .I(N__31058));
    InMux I__7100 (
            .O(N__31221),
            .I(N__31058));
    InMux I__7099 (
            .O(N__31220),
            .I(N__31051));
    InMux I__7098 (
            .O(N__31217),
            .I(N__31051));
    InMux I__7097 (
            .O(N__31216),
            .I(N__31051));
    CascadeMux I__7096 (
            .O(N__31215),
            .I(N__31045));
    CascadeMux I__7095 (
            .O(N__31214),
            .I(N__31042));
    InMux I__7094 (
            .O(N__31213),
            .I(N__31036));
    InMux I__7093 (
            .O(N__31212),
            .I(N__31036));
    InMux I__7092 (
            .O(N__31211),
            .I(N__31031));
    InMux I__7091 (
            .O(N__31210),
            .I(N__31031));
    InMux I__7090 (
            .O(N__31209),
            .I(N__31022));
    InMux I__7089 (
            .O(N__31208),
            .I(N__31022));
    InMux I__7088 (
            .O(N__31207),
            .I(N__31022));
    InMux I__7087 (
            .O(N__31206),
            .I(N__31022));
    LocalMux I__7086 (
            .O(N__31203),
            .I(N__31019));
    LocalMux I__7085 (
            .O(N__31196),
            .I(N__31016));
    LocalMux I__7084 (
            .O(N__31189),
            .I(N__31013));
    InMux I__7083 (
            .O(N__31188),
            .I(N__31008));
    InMux I__7082 (
            .O(N__31187),
            .I(N__31008));
    LocalMux I__7081 (
            .O(N__31182),
            .I(N__31003));
    LocalMux I__7080 (
            .O(N__31175),
            .I(N__31003));
    InMux I__7079 (
            .O(N__31174),
            .I(N__30998));
    InMux I__7078 (
            .O(N__31173),
            .I(N__30998));
    LocalMux I__7077 (
            .O(N__31168),
            .I(N__30995));
    InMux I__7076 (
            .O(N__31167),
            .I(N__30986));
    InMux I__7075 (
            .O(N__31166),
            .I(N__30986));
    InMux I__7074 (
            .O(N__31165),
            .I(N__30986));
    InMux I__7073 (
            .O(N__31164),
            .I(N__30986));
    InMux I__7072 (
            .O(N__31163),
            .I(N__30975));
    InMux I__7071 (
            .O(N__31162),
            .I(N__30975));
    InMux I__7070 (
            .O(N__31161),
            .I(N__30975));
    InMux I__7069 (
            .O(N__31160),
            .I(N__30975));
    InMux I__7068 (
            .O(N__31159),
            .I(N__30975));
    LocalMux I__7067 (
            .O(N__31156),
            .I(N__30967));
    Span4Mux_s3_v I__7066 (
            .O(N__31151),
            .I(N__30956));
    LocalMux I__7065 (
            .O(N__31148),
            .I(N__30956));
    Span4Mux_h I__7064 (
            .O(N__31145),
            .I(N__30956));
    Span4Mux_h I__7063 (
            .O(N__31138),
            .I(N__30956));
    LocalMux I__7062 (
            .O(N__31131),
            .I(N__30956));
    InMux I__7061 (
            .O(N__31130),
            .I(N__30951));
    LocalMux I__7060 (
            .O(N__31127),
            .I(N__30948));
    Span4Mux_s3_h I__7059 (
            .O(N__31122),
            .I(N__30943));
    LocalMux I__7058 (
            .O(N__31113),
            .I(N__30943));
    InMux I__7057 (
            .O(N__31112),
            .I(N__30940));
    CascadeMux I__7056 (
            .O(N__31111),
            .I(N__30934));
    InMux I__7055 (
            .O(N__31110),
            .I(N__30931));
    LocalMux I__7054 (
            .O(N__31105),
            .I(N__30926));
    Span4Mux_v I__7053 (
            .O(N__31102),
            .I(N__30926));
    LocalMux I__7052 (
            .O(N__31097),
            .I(N__30923));
    InMux I__7051 (
            .O(N__31096),
            .I(N__30916));
    InMux I__7050 (
            .O(N__31095),
            .I(N__30916));
    InMux I__7049 (
            .O(N__31094),
            .I(N__30916));
    InMux I__7048 (
            .O(N__31093),
            .I(N__30913));
    InMux I__7047 (
            .O(N__31092),
            .I(N__30908));
    InMux I__7046 (
            .O(N__31091),
            .I(N__30908));
    InMux I__7045 (
            .O(N__31090),
            .I(N__30901));
    InMux I__7044 (
            .O(N__31089),
            .I(N__30901));
    InMux I__7043 (
            .O(N__31088),
            .I(N__30898));
    InMux I__7042 (
            .O(N__31087),
            .I(N__30893));
    InMux I__7041 (
            .O(N__31086),
            .I(N__30893));
    LocalMux I__7040 (
            .O(N__31083),
            .I(N__30886));
    LocalMux I__7039 (
            .O(N__31080),
            .I(N__30886));
    LocalMux I__7038 (
            .O(N__31073),
            .I(N__30886));
    InMux I__7037 (
            .O(N__31072),
            .I(N__30881));
    InMux I__7036 (
            .O(N__31071),
            .I(N__30881));
    InMux I__7035 (
            .O(N__31070),
            .I(N__30874));
    InMux I__7034 (
            .O(N__31069),
            .I(N__30874));
    InMux I__7033 (
            .O(N__31068),
            .I(N__30874));
    LocalMux I__7032 (
            .O(N__31065),
            .I(N__30867));
    LocalMux I__7031 (
            .O(N__31058),
            .I(N__30867));
    LocalMux I__7030 (
            .O(N__31051),
            .I(N__30867));
    InMux I__7029 (
            .O(N__31050),
            .I(N__30860));
    InMux I__7028 (
            .O(N__31049),
            .I(N__30860));
    InMux I__7027 (
            .O(N__31048),
            .I(N__30860));
    InMux I__7026 (
            .O(N__31045),
            .I(N__30854));
    InMux I__7025 (
            .O(N__31042),
            .I(N__30851));
    InMux I__7024 (
            .O(N__31041),
            .I(N__30848));
    LocalMux I__7023 (
            .O(N__31036),
            .I(N__30843));
    LocalMux I__7022 (
            .O(N__31031),
            .I(N__30843));
    LocalMux I__7021 (
            .O(N__31022),
            .I(N__30832));
    Span4Mux_v I__7020 (
            .O(N__31019),
            .I(N__30832));
    Span4Mux_v I__7019 (
            .O(N__31016),
            .I(N__30832));
    Span4Mux_s1_h I__7018 (
            .O(N__31013),
            .I(N__30832));
    LocalMux I__7017 (
            .O(N__31008),
            .I(N__30832));
    Span4Mux_h I__7016 (
            .O(N__31003),
            .I(N__30821));
    LocalMux I__7015 (
            .O(N__30998),
            .I(N__30821));
    Span4Mux_v I__7014 (
            .O(N__30995),
            .I(N__30821));
    LocalMux I__7013 (
            .O(N__30986),
            .I(N__30821));
    LocalMux I__7012 (
            .O(N__30975),
            .I(N__30821));
    CascadeMux I__7011 (
            .O(N__30974),
            .I(N__30818));
    InMux I__7010 (
            .O(N__30973),
            .I(N__30815));
    InMux I__7009 (
            .O(N__30972),
            .I(N__30808));
    InMux I__7008 (
            .O(N__30971),
            .I(N__30808));
    InMux I__7007 (
            .O(N__30970),
            .I(N__30808));
    Span4Mux_s3_v I__7006 (
            .O(N__30967),
            .I(N__30803));
    Span4Mux_h I__7005 (
            .O(N__30956),
            .I(N__30803));
    InMux I__7004 (
            .O(N__30955),
            .I(N__30798));
    InMux I__7003 (
            .O(N__30954),
            .I(N__30798));
    LocalMux I__7002 (
            .O(N__30951),
            .I(N__30789));
    Span4Mux_v I__7001 (
            .O(N__30948),
            .I(N__30789));
    Span4Mux_h I__7000 (
            .O(N__30943),
            .I(N__30789));
    LocalMux I__6999 (
            .O(N__30940),
            .I(N__30789));
    InMux I__6998 (
            .O(N__30939),
            .I(N__30778));
    InMux I__6997 (
            .O(N__30938),
            .I(N__30778));
    InMux I__6996 (
            .O(N__30937),
            .I(N__30778));
    InMux I__6995 (
            .O(N__30934),
            .I(N__30775));
    LocalMux I__6994 (
            .O(N__30931),
            .I(N__30764));
    Span4Mux_h I__6993 (
            .O(N__30926),
            .I(N__30764));
    Span4Mux_v I__6992 (
            .O(N__30923),
            .I(N__30764));
    LocalMux I__6991 (
            .O(N__30916),
            .I(N__30764));
    LocalMux I__6990 (
            .O(N__30913),
            .I(N__30764));
    LocalMux I__6989 (
            .O(N__30908),
            .I(N__30761));
    InMux I__6988 (
            .O(N__30907),
            .I(N__30756));
    InMux I__6987 (
            .O(N__30906),
            .I(N__30756));
    LocalMux I__6986 (
            .O(N__30901),
            .I(N__30747));
    LocalMux I__6985 (
            .O(N__30898),
            .I(N__30747));
    LocalMux I__6984 (
            .O(N__30893),
            .I(N__30747));
    Span4Mux_v I__6983 (
            .O(N__30886),
            .I(N__30747));
    LocalMux I__6982 (
            .O(N__30881),
            .I(N__30738));
    LocalMux I__6981 (
            .O(N__30874),
            .I(N__30738));
    Span4Mux_v I__6980 (
            .O(N__30867),
            .I(N__30738));
    LocalMux I__6979 (
            .O(N__30860),
            .I(N__30738));
    InMux I__6978 (
            .O(N__30859),
            .I(N__30733));
    InMux I__6977 (
            .O(N__30858),
            .I(N__30733));
    CascadeMux I__6976 (
            .O(N__30857),
            .I(N__30730));
    LocalMux I__6975 (
            .O(N__30854),
            .I(N__30722));
    LocalMux I__6974 (
            .O(N__30851),
            .I(N__30722));
    LocalMux I__6973 (
            .O(N__30848),
            .I(N__30711));
    Span4Mux_v I__6972 (
            .O(N__30843),
            .I(N__30704));
    Span4Mux_h I__6971 (
            .O(N__30832),
            .I(N__30704));
    Span4Mux_v I__6970 (
            .O(N__30821),
            .I(N__30704));
    InMux I__6969 (
            .O(N__30818),
            .I(N__30701));
    LocalMux I__6968 (
            .O(N__30815),
            .I(N__30694));
    LocalMux I__6967 (
            .O(N__30808),
            .I(N__30694));
    Span4Mux_v I__6966 (
            .O(N__30803),
            .I(N__30694));
    LocalMux I__6965 (
            .O(N__30798),
            .I(N__30689));
    Span4Mux_v I__6964 (
            .O(N__30789),
            .I(N__30689));
    InMux I__6963 (
            .O(N__30788),
            .I(N__30682));
    InMux I__6962 (
            .O(N__30787),
            .I(N__30682));
    InMux I__6961 (
            .O(N__30786),
            .I(N__30682));
    InMux I__6960 (
            .O(N__30785),
            .I(N__30679));
    LocalMux I__6959 (
            .O(N__30778),
            .I(N__30676));
    LocalMux I__6958 (
            .O(N__30775),
            .I(N__30673));
    Span4Mux_h I__6957 (
            .O(N__30764),
            .I(N__30668));
    Span4Mux_s3_h I__6956 (
            .O(N__30761),
            .I(N__30668));
    LocalMux I__6955 (
            .O(N__30756),
            .I(N__30659));
    Span4Mux_h I__6954 (
            .O(N__30747),
            .I(N__30659));
    Span4Mux_v I__6953 (
            .O(N__30738),
            .I(N__30659));
    LocalMux I__6952 (
            .O(N__30733),
            .I(N__30659));
    InMux I__6951 (
            .O(N__30730),
            .I(N__30656));
    InMux I__6950 (
            .O(N__30729),
            .I(N__30649));
    InMux I__6949 (
            .O(N__30728),
            .I(N__30649));
    InMux I__6948 (
            .O(N__30727),
            .I(N__30649));
    Span4Mux_s3_h I__6947 (
            .O(N__30722),
            .I(N__30646));
    InMux I__6946 (
            .O(N__30721),
            .I(N__30641));
    InMux I__6945 (
            .O(N__30720),
            .I(N__30641));
    InMux I__6944 (
            .O(N__30719),
            .I(N__30636));
    InMux I__6943 (
            .O(N__30718),
            .I(N__30636));
    InMux I__6942 (
            .O(N__30717),
            .I(N__30629));
    InMux I__6941 (
            .O(N__30716),
            .I(N__30629));
    InMux I__6940 (
            .O(N__30715),
            .I(N__30629));
    InMux I__6939 (
            .O(N__30714),
            .I(N__30626));
    Span4Mux_v I__6938 (
            .O(N__30711),
            .I(N__30621));
    Span4Mux_h I__6937 (
            .O(N__30704),
            .I(N__30621));
    LocalMux I__6936 (
            .O(N__30701),
            .I(N__30614));
    Span4Mux_v I__6935 (
            .O(N__30694),
            .I(N__30614));
    Span4Mux_h I__6934 (
            .O(N__30689),
            .I(N__30614));
    LocalMux I__6933 (
            .O(N__30682),
            .I(N__30607));
    LocalMux I__6932 (
            .O(N__30679),
            .I(N__30607));
    Span12Mux_s11_v I__6931 (
            .O(N__30676),
            .I(N__30607));
    Span4Mux_v I__6930 (
            .O(N__30673),
            .I(N__30598));
    Span4Mux_v I__6929 (
            .O(N__30668),
            .I(N__30598));
    Span4Mux_h I__6928 (
            .O(N__30659),
            .I(N__30598));
    LocalMux I__6927 (
            .O(N__30656),
            .I(N__30598));
    LocalMux I__6926 (
            .O(N__30649),
            .I(\tok.T_0 ));
    Odrv4 I__6925 (
            .O(N__30646),
            .I(\tok.T_0 ));
    LocalMux I__6924 (
            .O(N__30641),
            .I(\tok.T_0 ));
    LocalMux I__6923 (
            .O(N__30636),
            .I(\tok.T_0 ));
    LocalMux I__6922 (
            .O(N__30629),
            .I(\tok.T_0 ));
    LocalMux I__6921 (
            .O(N__30626),
            .I(\tok.T_0 ));
    Odrv4 I__6920 (
            .O(N__30621),
            .I(\tok.T_0 ));
    Odrv4 I__6919 (
            .O(N__30614),
            .I(\tok.T_0 ));
    Odrv12 I__6918 (
            .O(N__30607),
            .I(\tok.T_0 ));
    Odrv4 I__6917 (
            .O(N__30598),
            .I(\tok.T_0 ));
    CascadeMux I__6916 (
            .O(N__30577),
            .I(N__30574));
    InMux I__6915 (
            .O(N__30574),
            .I(N__30571));
    LocalMux I__6914 (
            .O(N__30571),
            .I(\tok.n168_adj_690 ));
    InMux I__6913 (
            .O(N__30568),
            .I(N__30565));
    LocalMux I__6912 (
            .O(N__30565),
            .I(N__30562));
    Span4Mux_s3_h I__6911 (
            .O(N__30562),
            .I(N__30559));
    Span4Mux_h I__6910 (
            .O(N__30559),
            .I(N__30556));
    Odrv4 I__6909 (
            .O(N__30556),
            .I(\tok.n6525 ));
    CascadeMux I__6908 (
            .O(N__30553),
            .I(\tok.n6526_cascade_ ));
    CascadeMux I__6907 (
            .O(N__30550),
            .I(\tok.n186_adj_777_cascade_ ));
    CascadeMux I__6906 (
            .O(N__30547),
            .I(N__30544));
    InMux I__6905 (
            .O(N__30544),
            .I(N__30541));
    LocalMux I__6904 (
            .O(N__30541),
            .I(N__30538));
    Odrv12 I__6903 (
            .O(N__30538),
            .I(\tok.n338_adj_787 ));
    CascadeMux I__6902 (
            .O(N__30535),
            .I(N__30528));
    CascadeMux I__6901 (
            .O(N__30534),
            .I(N__30521));
    InMux I__6900 (
            .O(N__30533),
            .I(N__30518));
    InMux I__6899 (
            .O(N__30532),
            .I(N__30515));
    InMux I__6898 (
            .O(N__30531),
            .I(N__30512));
    InMux I__6897 (
            .O(N__30528),
            .I(N__30504));
    CascadeMux I__6896 (
            .O(N__30527),
            .I(N__30500));
    InMux I__6895 (
            .O(N__30526),
            .I(N__30496));
    InMux I__6894 (
            .O(N__30525),
            .I(N__30493));
    InMux I__6893 (
            .O(N__30524),
            .I(N__30488));
    InMux I__6892 (
            .O(N__30521),
            .I(N__30488));
    LocalMux I__6891 (
            .O(N__30518),
            .I(N__30482));
    LocalMux I__6890 (
            .O(N__30515),
            .I(N__30482));
    LocalMux I__6889 (
            .O(N__30512),
            .I(N__30479));
    InMux I__6888 (
            .O(N__30511),
            .I(N__30475));
    InMux I__6887 (
            .O(N__30510),
            .I(N__30470));
    InMux I__6886 (
            .O(N__30509),
            .I(N__30470));
    CascadeMux I__6885 (
            .O(N__30508),
            .I(N__30467));
    InMux I__6884 (
            .O(N__30507),
            .I(N__30464));
    LocalMux I__6883 (
            .O(N__30504),
            .I(N__30461));
    InMux I__6882 (
            .O(N__30503),
            .I(N__30458));
    InMux I__6881 (
            .O(N__30500),
            .I(N__30455));
    CascadeMux I__6880 (
            .O(N__30499),
            .I(N__30452));
    LocalMux I__6879 (
            .O(N__30496),
            .I(N__30449));
    LocalMux I__6878 (
            .O(N__30493),
            .I(N__30446));
    LocalMux I__6877 (
            .O(N__30488),
            .I(N__30443));
    InMux I__6876 (
            .O(N__30487),
            .I(N__30440));
    Span4Mux_s3_v I__6875 (
            .O(N__30482),
            .I(N__30435));
    Span4Mux_h I__6874 (
            .O(N__30479),
            .I(N__30435));
    InMux I__6873 (
            .O(N__30478),
            .I(N__30432));
    LocalMux I__6872 (
            .O(N__30475),
            .I(N__30429));
    LocalMux I__6871 (
            .O(N__30470),
            .I(N__30426));
    InMux I__6870 (
            .O(N__30467),
            .I(N__30423));
    LocalMux I__6869 (
            .O(N__30464),
            .I(N__30414));
    Span4Mux_v I__6868 (
            .O(N__30461),
            .I(N__30414));
    LocalMux I__6867 (
            .O(N__30458),
            .I(N__30414));
    LocalMux I__6866 (
            .O(N__30455),
            .I(N__30414));
    InMux I__6865 (
            .O(N__30452),
            .I(N__30411));
    Span4Mux_v I__6864 (
            .O(N__30449),
            .I(N__30407));
    Span4Mux_v I__6863 (
            .O(N__30446),
            .I(N__30404));
    Span4Mux_s3_v I__6862 (
            .O(N__30443),
            .I(N__30395));
    LocalMux I__6861 (
            .O(N__30440),
            .I(N__30395));
    Span4Mux_h I__6860 (
            .O(N__30435),
            .I(N__30395));
    LocalMux I__6859 (
            .O(N__30432),
            .I(N__30395));
    Span4Mux_v I__6858 (
            .O(N__30429),
            .I(N__30382));
    Span4Mux_v I__6857 (
            .O(N__30426),
            .I(N__30382));
    LocalMux I__6856 (
            .O(N__30423),
            .I(N__30382));
    Span4Mux_v I__6855 (
            .O(N__30414),
            .I(N__30382));
    LocalMux I__6854 (
            .O(N__30411),
            .I(N__30379));
    InMux I__6853 (
            .O(N__30410),
            .I(N__30376));
    Span4Mux_h I__6852 (
            .O(N__30407),
            .I(N__30369));
    Span4Mux_h I__6851 (
            .O(N__30404),
            .I(N__30369));
    Span4Mux_v I__6850 (
            .O(N__30395),
            .I(N__30369));
    InMux I__6849 (
            .O(N__30394),
            .I(N__30360));
    InMux I__6848 (
            .O(N__30393),
            .I(N__30360));
    InMux I__6847 (
            .O(N__30392),
            .I(N__30360));
    InMux I__6846 (
            .O(N__30391),
            .I(N__30360));
    Span4Mux_h I__6845 (
            .O(N__30382),
            .I(N__30357));
    Odrv12 I__6844 (
            .O(N__30379),
            .I(\tok.A_low_0 ));
    LocalMux I__6843 (
            .O(N__30376),
            .I(\tok.A_low_0 ));
    Odrv4 I__6842 (
            .O(N__30369),
            .I(\tok.A_low_0 ));
    LocalMux I__6841 (
            .O(N__30360),
            .I(\tok.A_low_0 ));
    Odrv4 I__6840 (
            .O(N__30357),
            .I(\tok.A_low_0 ));
    InMux I__6839 (
            .O(N__30346),
            .I(N__30339));
    CascadeMux I__6838 (
            .O(N__30345),
            .I(N__30336));
    InMux I__6837 (
            .O(N__30344),
            .I(N__30333));
    InMux I__6836 (
            .O(N__30343),
            .I(N__30330));
    CascadeMux I__6835 (
            .O(N__30342),
            .I(N__30315));
    LocalMux I__6834 (
            .O(N__30339),
            .I(N__30309));
    InMux I__6833 (
            .O(N__30336),
            .I(N__30306));
    LocalMux I__6832 (
            .O(N__30333),
            .I(N__30303));
    LocalMux I__6831 (
            .O(N__30330),
            .I(N__30300));
    InMux I__6830 (
            .O(N__30329),
            .I(N__30293));
    InMux I__6829 (
            .O(N__30328),
            .I(N__30293));
    InMux I__6828 (
            .O(N__30327),
            .I(N__30293));
    InMux I__6827 (
            .O(N__30326),
            .I(N__30286));
    InMux I__6826 (
            .O(N__30325),
            .I(N__30286));
    InMux I__6825 (
            .O(N__30324),
            .I(N__30286));
    InMux I__6824 (
            .O(N__30323),
            .I(N__30283));
    InMux I__6823 (
            .O(N__30322),
            .I(N__30280));
    InMux I__6822 (
            .O(N__30321),
            .I(N__30277));
    InMux I__6821 (
            .O(N__30320),
            .I(N__30274));
    InMux I__6820 (
            .O(N__30319),
            .I(N__30271));
    InMux I__6819 (
            .O(N__30318),
            .I(N__30268));
    InMux I__6818 (
            .O(N__30315),
            .I(N__30265));
    InMux I__6817 (
            .O(N__30314),
            .I(N__30260));
    InMux I__6816 (
            .O(N__30313),
            .I(N__30260));
    CascadeMux I__6815 (
            .O(N__30312),
            .I(N__30255));
    Span4Mux_s2_h I__6814 (
            .O(N__30309),
            .I(N__30250));
    LocalMux I__6813 (
            .O(N__30306),
            .I(N__30250));
    Span4Mux_s3_h I__6812 (
            .O(N__30303),
            .I(N__30247));
    Span4Mux_s3_h I__6811 (
            .O(N__30300),
            .I(N__30240));
    LocalMux I__6810 (
            .O(N__30293),
            .I(N__30240));
    LocalMux I__6809 (
            .O(N__30286),
            .I(N__30240));
    LocalMux I__6808 (
            .O(N__30283),
            .I(N__30237));
    LocalMux I__6807 (
            .O(N__30280),
            .I(N__30232));
    LocalMux I__6806 (
            .O(N__30277),
            .I(N__30232));
    LocalMux I__6805 (
            .O(N__30274),
            .I(N__30227));
    LocalMux I__6804 (
            .O(N__30271),
            .I(N__30227));
    LocalMux I__6803 (
            .O(N__30268),
            .I(N__30222));
    LocalMux I__6802 (
            .O(N__30265),
            .I(N__30222));
    LocalMux I__6801 (
            .O(N__30260),
            .I(N__30219));
    InMux I__6800 (
            .O(N__30259),
            .I(N__30214));
    InMux I__6799 (
            .O(N__30258),
            .I(N__30214));
    InMux I__6798 (
            .O(N__30255),
            .I(N__30211));
    Span4Mux_h I__6797 (
            .O(N__30250),
            .I(N__30206));
    Span4Mux_h I__6796 (
            .O(N__30247),
            .I(N__30206));
    Span4Mux_h I__6795 (
            .O(N__30240),
            .I(N__30203));
    Span4Mux_v I__6794 (
            .O(N__30237),
            .I(N__30194));
    Span4Mux_h I__6793 (
            .O(N__30232),
            .I(N__30194));
    Span4Mux_v I__6792 (
            .O(N__30227),
            .I(N__30194));
    Span4Mux_v I__6791 (
            .O(N__30222),
            .I(N__30194));
    Odrv12 I__6790 (
            .O(N__30219),
            .I(\tok.A_low_5 ));
    LocalMux I__6789 (
            .O(N__30214),
            .I(\tok.A_low_5 ));
    LocalMux I__6788 (
            .O(N__30211),
            .I(\tok.A_low_5 ));
    Odrv4 I__6787 (
            .O(N__30206),
            .I(\tok.A_low_5 ));
    Odrv4 I__6786 (
            .O(N__30203),
            .I(\tok.A_low_5 ));
    Odrv4 I__6785 (
            .O(N__30194),
            .I(\tok.A_low_5 ));
    CascadeMux I__6784 (
            .O(N__30181),
            .I(\tok.n866_cascade_ ));
    InMux I__6783 (
            .O(N__30178),
            .I(N__30175));
    LocalMux I__6782 (
            .O(N__30175),
            .I(\tok.n6520 ));
    CascadeMux I__6781 (
            .O(N__30172),
            .I(\tok.n10_cascade_ ));
    SRMux I__6780 (
            .O(N__30169),
            .I(N__30166));
    LocalMux I__6779 (
            .O(N__30166),
            .I(N__30163));
    Span4Mux_h I__6778 (
            .O(N__30163),
            .I(N__30160));
    Span4Mux_h I__6777 (
            .O(N__30160),
            .I(N__30157));
    Span4Mux_s2_v I__6776 (
            .O(N__30157),
            .I(N__30154));
    Span4Mux_v I__6775 (
            .O(N__30154),
            .I(N__30151));
    Odrv4 I__6774 (
            .O(N__30151),
            .I(\tok.write_flag ));
    InMux I__6773 (
            .O(N__30148),
            .I(N__30135));
    InMux I__6772 (
            .O(N__30147),
            .I(N__30135));
    InMux I__6771 (
            .O(N__30146),
            .I(N__30135));
    InMux I__6770 (
            .O(N__30145),
            .I(N__30131));
    InMux I__6769 (
            .O(N__30144),
            .I(N__30124));
    InMux I__6768 (
            .O(N__30143),
            .I(N__30124));
    InMux I__6767 (
            .O(N__30142),
            .I(N__30124));
    LocalMux I__6766 (
            .O(N__30135),
            .I(N__30121));
    InMux I__6765 (
            .O(N__30134),
            .I(N__30118));
    LocalMux I__6764 (
            .O(N__30131),
            .I(N__30113));
    LocalMux I__6763 (
            .O(N__30124),
            .I(N__30113));
    Span4Mux_v I__6762 (
            .O(N__30121),
            .I(N__30110));
    LocalMux I__6761 (
            .O(N__30118),
            .I(N__30105));
    Span4Mux_h I__6760 (
            .O(N__30113),
            .I(N__30105));
    Sp12to4 I__6759 (
            .O(N__30110),
            .I(N__30102));
    Span4Mux_v I__6758 (
            .O(N__30105),
            .I(N__30099));
    Odrv12 I__6757 (
            .O(N__30102),
            .I(\tok.n14 ));
    Odrv4 I__6756 (
            .O(N__30099),
            .I(\tok.n14 ));
    CascadeMux I__6755 (
            .O(N__30094),
            .I(\tok.uart.n10_cascade_ ));
    CascadeMux I__6754 (
            .O(N__30091),
            .I(n23_cascade_));
    CascadeMux I__6753 (
            .O(N__30088),
            .I(\tok.n168_adj_710_cascade_ ));
    InMux I__6752 (
            .O(N__30085),
            .I(N__30080));
    InMux I__6751 (
            .O(N__30084),
            .I(N__30075));
    InMux I__6750 (
            .O(N__30083),
            .I(N__30075));
    LocalMux I__6749 (
            .O(N__30080),
            .I(N__30067));
    LocalMux I__6748 (
            .O(N__30075),
            .I(N__30067));
    CascadeMux I__6747 (
            .O(N__30074),
            .I(N__30059));
    InMux I__6746 (
            .O(N__30073),
            .I(N__30055));
    InMux I__6745 (
            .O(N__30072),
            .I(N__30050));
    Span4Mux_h I__6744 (
            .O(N__30067),
            .I(N__30047));
    CascadeMux I__6743 (
            .O(N__30066),
            .I(N__30044));
    CascadeMux I__6742 (
            .O(N__30065),
            .I(N__30039));
    InMux I__6741 (
            .O(N__30064),
            .I(N__30035));
    InMux I__6740 (
            .O(N__30063),
            .I(N__30032));
    InMux I__6739 (
            .O(N__30062),
            .I(N__30029));
    InMux I__6738 (
            .O(N__30059),
            .I(N__30023));
    InMux I__6737 (
            .O(N__30058),
            .I(N__30020));
    LocalMux I__6736 (
            .O(N__30055),
            .I(N__30017));
    InMux I__6735 (
            .O(N__30054),
            .I(N__30014));
    CascadeMux I__6734 (
            .O(N__30053),
            .I(N__30011));
    LocalMux I__6733 (
            .O(N__30050),
            .I(N__30005));
    IoSpan4Mux I__6732 (
            .O(N__30047),
            .I(N__30005));
    InMux I__6731 (
            .O(N__30044),
            .I(N__30000));
    InMux I__6730 (
            .O(N__30043),
            .I(N__30000));
    InMux I__6729 (
            .O(N__30042),
            .I(N__29997));
    InMux I__6728 (
            .O(N__30039),
            .I(N__29994));
    InMux I__6727 (
            .O(N__30038),
            .I(N__29991));
    LocalMux I__6726 (
            .O(N__30035),
            .I(N__29988));
    LocalMux I__6725 (
            .O(N__30032),
            .I(N__29985));
    LocalMux I__6724 (
            .O(N__30029),
            .I(N__29982));
    InMux I__6723 (
            .O(N__30028),
            .I(N__29977));
    InMux I__6722 (
            .O(N__30027),
            .I(N__29977));
    InMux I__6721 (
            .O(N__30026),
            .I(N__29974));
    LocalMux I__6720 (
            .O(N__30023),
            .I(N__29971));
    LocalMux I__6719 (
            .O(N__30020),
            .I(N__29968));
    Span4Mux_s3_v I__6718 (
            .O(N__30017),
            .I(N__29963));
    LocalMux I__6717 (
            .O(N__30014),
            .I(N__29963));
    InMux I__6716 (
            .O(N__30011),
            .I(N__29960));
    InMux I__6715 (
            .O(N__30010),
            .I(N__29957));
    Span4Mux_s2_v I__6714 (
            .O(N__30005),
            .I(N__29948));
    LocalMux I__6713 (
            .O(N__30000),
            .I(N__29948));
    LocalMux I__6712 (
            .O(N__29997),
            .I(N__29948));
    LocalMux I__6711 (
            .O(N__29994),
            .I(N__29948));
    LocalMux I__6710 (
            .O(N__29991),
            .I(N__29945));
    Span4Mux_v I__6709 (
            .O(N__29988),
            .I(N__29942));
    Span4Mux_v I__6708 (
            .O(N__29985),
            .I(N__29939));
    Span4Mux_v I__6707 (
            .O(N__29982),
            .I(N__29932));
    LocalMux I__6706 (
            .O(N__29977),
            .I(N__29932));
    LocalMux I__6705 (
            .O(N__29974),
            .I(N__29932));
    Span4Mux_s2_v I__6704 (
            .O(N__29971),
            .I(N__29926));
    Span4Mux_h I__6703 (
            .O(N__29968),
            .I(N__29926));
    Span4Mux_v I__6702 (
            .O(N__29963),
            .I(N__29917));
    LocalMux I__6701 (
            .O(N__29960),
            .I(N__29917));
    LocalMux I__6700 (
            .O(N__29957),
            .I(N__29917));
    Span4Mux_v I__6699 (
            .O(N__29948),
            .I(N__29917));
    Span12Mux_s8_v I__6698 (
            .O(N__29945),
            .I(N__29912));
    Sp12to4 I__6697 (
            .O(N__29942),
            .I(N__29912));
    Span4Mux_v I__6696 (
            .O(N__29939),
            .I(N__29907));
    Span4Mux_v I__6695 (
            .O(N__29932),
            .I(N__29907));
    InMux I__6694 (
            .O(N__29931),
            .I(N__29904));
    Span4Mux_v I__6693 (
            .O(N__29926),
            .I(N__29899));
    Span4Mux_h I__6692 (
            .O(N__29917),
            .I(N__29899));
    Odrv12 I__6691 (
            .O(N__29912),
            .I(\tok.A_low_6 ));
    Odrv4 I__6690 (
            .O(N__29907),
            .I(\tok.A_low_6 ));
    LocalMux I__6689 (
            .O(N__29904),
            .I(\tok.A_low_6 ));
    Odrv4 I__6688 (
            .O(N__29899),
            .I(\tok.A_low_6 ));
    InMux I__6687 (
            .O(N__29890),
            .I(N__29887));
    LocalMux I__6686 (
            .O(N__29887),
            .I(\tok.n6502 ));
    InMux I__6685 (
            .O(N__29884),
            .I(N__29878));
    InMux I__6684 (
            .O(N__29883),
            .I(N__29878));
    LocalMux I__6683 (
            .O(N__29878),
            .I(uart_rx_data_6));
    InMux I__6682 (
            .O(N__29875),
            .I(N__29865));
    InMux I__6681 (
            .O(N__29874),
            .I(N__29865));
    InMux I__6680 (
            .O(N__29873),
            .I(N__29856));
    InMux I__6679 (
            .O(N__29872),
            .I(N__29856));
    InMux I__6678 (
            .O(N__29871),
            .I(N__29856));
    InMux I__6677 (
            .O(N__29870),
            .I(N__29856));
    LocalMux I__6676 (
            .O(N__29865),
            .I(\tok.depth_1 ));
    LocalMux I__6675 (
            .O(N__29856),
            .I(\tok.depth_1 ));
    CascadeMux I__6674 (
            .O(N__29851),
            .I(N__29848));
    InMux I__6673 (
            .O(N__29848),
            .I(N__29842));
    InMux I__6672 (
            .O(N__29847),
            .I(N__29842));
    LocalMux I__6671 (
            .O(N__29842),
            .I(\tok.n741 ));
    CascadeMux I__6670 (
            .O(N__29839),
            .I(N__29835));
    CascadeMux I__6669 (
            .O(N__29838),
            .I(N__29832));
    InMux I__6668 (
            .O(N__29835),
            .I(N__29827));
    InMux I__6667 (
            .O(N__29832),
            .I(N__29827));
    LocalMux I__6666 (
            .O(N__29827),
            .I(N__29824));
    Span4Mux_h I__6665 (
            .O(N__29824),
            .I(N__29821));
    Odrv4 I__6664 (
            .O(N__29821),
            .I(\tok.n806 ));
    CascadeMux I__6663 (
            .O(N__29818),
            .I(N__29815));
    InMux I__6662 (
            .O(N__29815),
            .I(N__29806));
    InMux I__6661 (
            .O(N__29814),
            .I(N__29806));
    InMux I__6660 (
            .O(N__29813),
            .I(N__29803));
    CascadeMux I__6659 (
            .O(N__29812),
            .I(N__29799));
    CascadeMux I__6658 (
            .O(N__29811),
            .I(N__29795));
    LocalMux I__6657 (
            .O(N__29806),
            .I(N__29789));
    LocalMux I__6656 (
            .O(N__29803),
            .I(N__29789));
    InMux I__6655 (
            .O(N__29802),
            .I(N__29784));
    InMux I__6654 (
            .O(N__29799),
            .I(N__29784));
    InMux I__6653 (
            .O(N__29798),
            .I(N__29777));
    InMux I__6652 (
            .O(N__29795),
            .I(N__29777));
    InMux I__6651 (
            .O(N__29794),
            .I(N__29777));
    Odrv4 I__6650 (
            .O(N__29789),
            .I(\tok.depth_0 ));
    LocalMux I__6649 (
            .O(N__29784),
            .I(\tok.depth_0 ));
    LocalMux I__6648 (
            .O(N__29777),
            .I(\tok.depth_0 ));
    InMux I__6647 (
            .O(N__29770),
            .I(N__29767));
    LocalMux I__6646 (
            .O(N__29767),
            .I(\tok.n6213 ));
    CascadeMux I__6645 (
            .O(N__29764),
            .I(\tok.n806_cascade_ ));
    CascadeMux I__6644 (
            .O(N__29761),
            .I(N__29754));
    CascadeMux I__6643 (
            .O(N__29760),
            .I(N__29750));
    InMux I__6642 (
            .O(N__29759),
            .I(N__29747));
    InMux I__6641 (
            .O(N__29758),
            .I(N__29744));
    InMux I__6640 (
            .O(N__29757),
            .I(N__29741));
    InMux I__6639 (
            .O(N__29754),
            .I(N__29734));
    InMux I__6638 (
            .O(N__29753),
            .I(N__29734));
    InMux I__6637 (
            .O(N__29750),
            .I(N__29734));
    LocalMux I__6636 (
            .O(N__29747),
            .I(\tok.depth_3 ));
    LocalMux I__6635 (
            .O(N__29744),
            .I(\tok.depth_3 ));
    LocalMux I__6634 (
            .O(N__29741),
            .I(\tok.depth_3 ));
    LocalMux I__6633 (
            .O(N__29734),
            .I(\tok.depth_3 ));
    CascadeMux I__6632 (
            .O(N__29725),
            .I(N__29720));
    CascadeMux I__6631 (
            .O(N__29724),
            .I(N__29715));
    CascadeMux I__6630 (
            .O(N__29723),
            .I(N__29712));
    InMux I__6629 (
            .O(N__29720),
            .I(N__29707));
    InMux I__6628 (
            .O(N__29719),
            .I(N__29703));
    InMux I__6627 (
            .O(N__29718),
            .I(N__29700));
    InMux I__6626 (
            .O(N__29715),
            .I(N__29697));
    InMux I__6625 (
            .O(N__29712),
            .I(N__29694));
    InMux I__6624 (
            .O(N__29711),
            .I(N__29691));
    InMux I__6623 (
            .O(N__29710),
            .I(N__29688));
    LocalMux I__6622 (
            .O(N__29707),
            .I(N__29685));
    InMux I__6621 (
            .O(N__29706),
            .I(N__29682));
    LocalMux I__6620 (
            .O(N__29703),
            .I(N__29677));
    LocalMux I__6619 (
            .O(N__29700),
            .I(N__29677));
    LocalMux I__6618 (
            .O(N__29697),
            .I(N__29674));
    LocalMux I__6617 (
            .O(N__29694),
            .I(N__29671));
    LocalMux I__6616 (
            .O(N__29691),
            .I(N__29668));
    LocalMux I__6615 (
            .O(N__29688),
            .I(N__29661));
    Span4Mux_h I__6614 (
            .O(N__29685),
            .I(N__29661));
    LocalMux I__6613 (
            .O(N__29682),
            .I(N__29661));
    Span4Mux_v I__6612 (
            .O(N__29677),
            .I(N__29658));
    Span4Mux_v I__6611 (
            .O(N__29674),
            .I(N__29653));
    Span4Mux_v I__6610 (
            .O(N__29671),
            .I(N__29653));
    Span4Mux_h I__6609 (
            .O(N__29668),
            .I(N__29650));
    Span4Mux_h I__6608 (
            .O(N__29661),
            .I(N__29647));
    Span4Mux_h I__6607 (
            .O(N__29658),
            .I(N__29644));
    Span4Mux_h I__6606 (
            .O(N__29653),
            .I(N__29641));
    Span4Mux_v I__6605 (
            .O(N__29650),
            .I(N__29634));
    Span4Mux_v I__6604 (
            .O(N__29647),
            .I(N__29634));
    Span4Mux_h I__6603 (
            .O(N__29644),
            .I(N__29634));
    Odrv4 I__6602 (
            .O(N__29641),
            .I(\tok.n748 ));
    Odrv4 I__6601 (
            .O(N__29634),
            .I(\tok.n748 ));
    InMux I__6600 (
            .O(N__29629),
            .I(N__29623));
    InMux I__6599 (
            .O(N__29628),
            .I(N__29614));
    InMux I__6598 (
            .O(N__29627),
            .I(N__29611));
    InMux I__6597 (
            .O(N__29626),
            .I(N__29608));
    LocalMux I__6596 (
            .O(N__29623),
            .I(N__29605));
    InMux I__6595 (
            .O(N__29622),
            .I(N__29600));
    InMux I__6594 (
            .O(N__29621),
            .I(N__29600));
    InMux I__6593 (
            .O(N__29620),
            .I(N__29597));
    InMux I__6592 (
            .O(N__29619),
            .I(N__29592));
    InMux I__6591 (
            .O(N__29618),
            .I(N__29587));
    InMux I__6590 (
            .O(N__29617),
            .I(N__29587));
    LocalMux I__6589 (
            .O(N__29614),
            .I(N__29584));
    LocalMux I__6588 (
            .O(N__29611),
            .I(N__29581));
    LocalMux I__6587 (
            .O(N__29608),
            .I(N__29578));
    Span4Mux_v I__6586 (
            .O(N__29605),
            .I(N__29572));
    LocalMux I__6585 (
            .O(N__29600),
            .I(N__29572));
    LocalMux I__6584 (
            .O(N__29597),
            .I(N__29569));
    CascadeMux I__6583 (
            .O(N__29596),
            .I(N__29566));
    InMux I__6582 (
            .O(N__29595),
            .I(N__29563));
    LocalMux I__6581 (
            .O(N__29592),
            .I(N__29559));
    LocalMux I__6580 (
            .O(N__29587),
            .I(N__29556));
    Span4Mux_h I__6579 (
            .O(N__29584),
            .I(N__29553));
    Span4Mux_h I__6578 (
            .O(N__29581),
            .I(N__29550));
    Span4Mux_v I__6577 (
            .O(N__29578),
            .I(N__29544));
    InMux I__6576 (
            .O(N__29577),
            .I(N__29541));
    Span4Mux_v I__6575 (
            .O(N__29572),
            .I(N__29536));
    Span4Mux_s3_h I__6574 (
            .O(N__29569),
            .I(N__29536));
    InMux I__6573 (
            .O(N__29566),
            .I(N__29533));
    LocalMux I__6572 (
            .O(N__29563),
            .I(N__29530));
    CascadeMux I__6571 (
            .O(N__29562),
            .I(N__29526));
    Span4Mux_v I__6570 (
            .O(N__29559),
            .I(N__29521));
    Span4Mux_v I__6569 (
            .O(N__29556),
            .I(N__29521));
    Span4Mux_v I__6568 (
            .O(N__29553),
            .I(N__29516));
    Span4Mux_h I__6567 (
            .O(N__29550),
            .I(N__29516));
    InMux I__6566 (
            .O(N__29549),
            .I(N__29509));
    InMux I__6565 (
            .O(N__29548),
            .I(N__29509));
    InMux I__6564 (
            .O(N__29547),
            .I(N__29509));
    Span4Mux_h I__6563 (
            .O(N__29544),
            .I(N__29504));
    LocalMux I__6562 (
            .O(N__29541),
            .I(N__29504));
    Span4Mux_h I__6561 (
            .O(N__29536),
            .I(N__29501));
    LocalMux I__6560 (
            .O(N__29533),
            .I(N__29496));
    Span12Mux_s7_h I__6559 (
            .O(N__29530),
            .I(N__29496));
    InMux I__6558 (
            .O(N__29529),
            .I(N__29491));
    InMux I__6557 (
            .O(N__29526),
            .I(N__29491));
    Odrv4 I__6556 (
            .O(N__29521),
            .I(\tok.n47 ));
    Odrv4 I__6555 (
            .O(N__29516),
            .I(\tok.n47 ));
    LocalMux I__6554 (
            .O(N__29509),
            .I(\tok.n47 ));
    Odrv4 I__6553 (
            .O(N__29504),
            .I(\tok.n47 ));
    Odrv4 I__6552 (
            .O(N__29501),
            .I(\tok.n47 ));
    Odrv12 I__6551 (
            .O(N__29496),
            .I(\tok.n47 ));
    LocalMux I__6550 (
            .O(N__29491),
            .I(\tok.n47 ));
    CascadeMux I__6549 (
            .O(N__29476),
            .I(N__29473));
    InMux I__6548 (
            .O(N__29473),
            .I(N__29470));
    LocalMux I__6547 (
            .O(N__29470),
            .I(N__29467));
    Span12Mux_s9_h I__6546 (
            .O(N__29467),
            .I(N__29464));
    Odrv12 I__6545 (
            .O(N__29464),
            .I(\tok.n6615 ));
    CascadeMux I__6544 (
            .O(N__29461),
            .I(\tok.n158_cascade_ ));
    InMux I__6543 (
            .O(N__29458),
            .I(N__29455));
    LocalMux I__6542 (
            .O(N__29455),
            .I(N__29452));
    Odrv4 I__6541 (
            .O(N__29452),
            .I(\tok.n6627 ));
    InMux I__6540 (
            .O(N__29449),
            .I(N__29440));
    InMux I__6539 (
            .O(N__29448),
            .I(N__29440));
    InMux I__6538 (
            .O(N__29447),
            .I(N__29440));
    LocalMux I__6537 (
            .O(N__29440),
            .I(N__29437));
    Span4Mux_h I__6536 (
            .O(N__29437),
            .I(N__29434));
    Span4Mux_h I__6535 (
            .O(N__29434),
            .I(N__29431));
    Odrv4 I__6534 (
            .O(N__29431),
            .I(\tok.uart_stall_N_46 ));
    InMux I__6533 (
            .O(N__29428),
            .I(N__29425));
    LocalMux I__6532 (
            .O(N__29425),
            .I(\tok.n9 ));
    CascadeMux I__6531 (
            .O(N__29422),
            .I(N__29419));
    InMux I__6530 (
            .O(N__29419),
            .I(N__29416));
    LocalMux I__6529 (
            .O(N__29416),
            .I(\tok.n10 ));
    InMux I__6528 (
            .O(N__29413),
            .I(N__29409));
    CascadeMux I__6527 (
            .O(N__29412),
            .I(N__29405));
    LocalMux I__6526 (
            .O(N__29409),
            .I(N__29402));
    InMux I__6525 (
            .O(N__29408),
            .I(N__29397));
    InMux I__6524 (
            .O(N__29405),
            .I(N__29392));
    Span12Mux_h I__6523 (
            .O(N__29402),
            .I(N__29389));
    InMux I__6522 (
            .O(N__29401),
            .I(N__29384));
    InMux I__6521 (
            .O(N__29400),
            .I(N__29384));
    LocalMux I__6520 (
            .O(N__29397),
            .I(N__29381));
    InMux I__6519 (
            .O(N__29396),
            .I(N__29376));
    InMux I__6518 (
            .O(N__29395),
            .I(N__29376));
    LocalMux I__6517 (
            .O(N__29392),
            .I(N__29373));
    Odrv12 I__6516 (
            .O(N__29389),
            .I(\tok.A_stk_delta_1__N_4 ));
    LocalMux I__6515 (
            .O(N__29384),
            .I(\tok.A_stk_delta_1__N_4 ));
    Odrv4 I__6514 (
            .O(N__29381),
            .I(\tok.A_stk_delta_1__N_4 ));
    LocalMux I__6513 (
            .O(N__29376),
            .I(\tok.A_stk_delta_1__N_4 ));
    Odrv4 I__6512 (
            .O(N__29373),
            .I(\tok.A_stk_delta_1__N_4 ));
    CascadeMux I__6511 (
            .O(N__29362),
            .I(\tok.A_stk_delta_1__N_4_cascade_ ));
    CascadeMux I__6510 (
            .O(N__29359),
            .I(N__29356));
    InMux I__6509 (
            .O(N__29356),
            .I(N__29347));
    InMux I__6508 (
            .O(N__29355),
            .I(N__29347));
    InMux I__6507 (
            .O(N__29354),
            .I(N__29347));
    LocalMux I__6506 (
            .O(N__29347),
            .I(N__29341));
    InMux I__6505 (
            .O(N__29346),
            .I(N__29334));
    InMux I__6504 (
            .O(N__29345),
            .I(N__29334));
    InMux I__6503 (
            .O(N__29344),
            .I(N__29334));
    Span4Mux_s1_h I__6502 (
            .O(N__29341),
            .I(N__29331));
    LocalMux I__6501 (
            .O(N__29334),
            .I(N__29328));
    Odrv4 I__6500 (
            .O(N__29331),
            .I(\tok.n1 ));
    Odrv12 I__6499 (
            .O(N__29328),
            .I(\tok.n1 ));
    CascadeMux I__6498 (
            .O(N__29323),
            .I(\tok.n4_adj_702_cascade_ ));
    InMux I__6497 (
            .O(N__29320),
            .I(N__29317));
    LocalMux I__6496 (
            .O(N__29317),
            .I(\tok.n52 ));
    CascadeMux I__6495 (
            .O(N__29314),
            .I(\tok.n51_cascade_ ));
    InMux I__6494 (
            .O(N__29311),
            .I(N__29308));
    LocalMux I__6493 (
            .O(N__29308),
            .I(\tok.n50 ));
    InMux I__6492 (
            .O(N__29305),
            .I(N__29302));
    LocalMux I__6491 (
            .O(N__29302),
            .I(\tok.n8_adj_854 ));
    InMux I__6490 (
            .O(N__29299),
            .I(N__29290));
    InMux I__6489 (
            .O(N__29298),
            .I(N__29290));
    InMux I__6488 (
            .O(N__29297),
            .I(N__29290));
    LocalMux I__6487 (
            .O(N__29290),
            .I(\tok.n174 ));
    InMux I__6486 (
            .O(N__29287),
            .I(N__29282));
    InMux I__6485 (
            .O(N__29286),
            .I(N__29277));
    InMux I__6484 (
            .O(N__29285),
            .I(N__29277));
    LocalMux I__6483 (
            .O(N__29282),
            .I(\tok.n4_adj_702 ));
    LocalMux I__6482 (
            .O(N__29277),
            .I(\tok.n4_adj_702 ));
    SRMux I__6481 (
            .O(N__29272),
            .I(N__29266));
    SRMux I__6480 (
            .O(N__29271),
            .I(N__29263));
    SRMux I__6479 (
            .O(N__29270),
            .I(N__29256));
    SRMux I__6478 (
            .O(N__29269),
            .I(N__29251));
    LocalMux I__6477 (
            .O(N__29266),
            .I(N__29246));
    LocalMux I__6476 (
            .O(N__29263),
            .I(N__29246));
    SRMux I__6475 (
            .O(N__29262),
            .I(N__29243));
    SRMux I__6474 (
            .O(N__29261),
            .I(N__29238));
    SRMux I__6473 (
            .O(N__29260),
            .I(N__29234));
    SRMux I__6472 (
            .O(N__29259),
            .I(N__29231));
    LocalMux I__6471 (
            .O(N__29256),
            .I(N__29227));
    SRMux I__6470 (
            .O(N__29255),
            .I(N__29224));
    SRMux I__6469 (
            .O(N__29254),
            .I(N__29221));
    LocalMux I__6468 (
            .O(N__29251),
            .I(N__29217));
    Span4Mux_s1_v I__6467 (
            .O(N__29246),
            .I(N__29211));
    LocalMux I__6466 (
            .O(N__29243),
            .I(N__29211));
    SRMux I__6465 (
            .O(N__29242),
            .I(N__29208));
    SRMux I__6464 (
            .O(N__29241),
            .I(N__29205));
    LocalMux I__6463 (
            .O(N__29238),
            .I(N__29201));
    SRMux I__6462 (
            .O(N__29237),
            .I(N__29198));
    LocalMux I__6461 (
            .O(N__29234),
            .I(N__29195));
    LocalMux I__6460 (
            .O(N__29231),
            .I(N__29192));
    SRMux I__6459 (
            .O(N__29230),
            .I(N__29189));
    Span4Mux_v I__6458 (
            .O(N__29227),
            .I(N__29184));
    LocalMux I__6457 (
            .O(N__29224),
            .I(N__29184));
    LocalMux I__6456 (
            .O(N__29221),
            .I(N__29181));
    SRMux I__6455 (
            .O(N__29220),
            .I(N__29176));
    Span4Mux_v I__6454 (
            .O(N__29217),
            .I(N__29173));
    SRMux I__6453 (
            .O(N__29216),
            .I(N__29170));
    Span4Mux_v I__6452 (
            .O(N__29211),
            .I(N__29163));
    LocalMux I__6451 (
            .O(N__29208),
            .I(N__29163));
    LocalMux I__6450 (
            .O(N__29205),
            .I(N__29160));
    SRMux I__6449 (
            .O(N__29204),
            .I(N__29157));
    Span4Mux_v I__6448 (
            .O(N__29201),
            .I(N__29152));
    LocalMux I__6447 (
            .O(N__29198),
            .I(N__29152));
    Span4Mux_h I__6446 (
            .O(N__29195),
            .I(N__29149));
    Span4Mux_v I__6445 (
            .O(N__29192),
            .I(N__29144));
    LocalMux I__6444 (
            .O(N__29189),
            .I(N__29144));
    Span4Mux_v I__6443 (
            .O(N__29184),
            .I(N__29141));
    Span4Mux_v I__6442 (
            .O(N__29181),
            .I(N__29138));
    SRMux I__6441 (
            .O(N__29180),
            .I(N__29135));
    SRMux I__6440 (
            .O(N__29179),
            .I(N__29132));
    LocalMux I__6439 (
            .O(N__29176),
            .I(N__29129));
    Span4Mux_v I__6438 (
            .O(N__29173),
            .I(N__29124));
    LocalMux I__6437 (
            .O(N__29170),
            .I(N__29124));
    SRMux I__6436 (
            .O(N__29169),
            .I(N__29121));
    SRMux I__6435 (
            .O(N__29168),
            .I(N__29118));
    Span4Mux_v I__6434 (
            .O(N__29163),
            .I(N__29113));
    Span4Mux_h I__6433 (
            .O(N__29160),
            .I(N__29108));
    LocalMux I__6432 (
            .O(N__29157),
            .I(N__29108));
    Span4Mux_h I__6431 (
            .O(N__29152),
            .I(N__29105));
    Span4Mux_v I__6430 (
            .O(N__29149),
            .I(N__29100));
    Span4Mux_h I__6429 (
            .O(N__29144),
            .I(N__29100));
    IoSpan4Mux I__6428 (
            .O(N__29141),
            .I(N__29097));
    Span4Mux_h I__6427 (
            .O(N__29138),
            .I(N__29092));
    LocalMux I__6426 (
            .O(N__29135),
            .I(N__29092));
    LocalMux I__6425 (
            .O(N__29132),
            .I(N__29089));
    Span4Mux_v I__6424 (
            .O(N__29129),
            .I(N__29086));
    Span4Mux_v I__6423 (
            .O(N__29124),
            .I(N__29081));
    LocalMux I__6422 (
            .O(N__29121),
            .I(N__29081));
    LocalMux I__6421 (
            .O(N__29118),
            .I(N__29078));
    SRMux I__6420 (
            .O(N__29117),
            .I(N__29075));
    SRMux I__6419 (
            .O(N__29116),
            .I(N__29072));
    Span4Mux_h I__6418 (
            .O(N__29113),
            .I(N__29067));
    Span4Mux_v I__6417 (
            .O(N__29108),
            .I(N__29067));
    Span4Mux_h I__6416 (
            .O(N__29105),
            .I(N__29062));
    Span4Mux_h I__6415 (
            .O(N__29100),
            .I(N__29062));
    Span4Mux_s0_v I__6414 (
            .O(N__29097),
            .I(N__29057));
    Span4Mux_v I__6413 (
            .O(N__29092),
            .I(N__29057));
    Span4Mux_v I__6412 (
            .O(N__29089),
            .I(N__29054));
    Span4Mux_h I__6411 (
            .O(N__29086),
            .I(N__29049));
    Span4Mux_h I__6410 (
            .O(N__29081),
            .I(N__29049));
    Span4Mux_h I__6409 (
            .O(N__29078),
            .I(N__29046));
    LocalMux I__6408 (
            .O(N__29075),
            .I(N__29043));
    LocalMux I__6407 (
            .O(N__29072),
            .I(N__29040));
    Span4Mux_v I__6406 (
            .O(N__29067),
            .I(N__29037));
    Span4Mux_v I__6405 (
            .O(N__29062),
            .I(N__29034));
    Span4Mux_h I__6404 (
            .O(N__29057),
            .I(N__29029));
    Span4Mux_h I__6403 (
            .O(N__29054),
            .I(N__29029));
    Span4Mux_h I__6402 (
            .O(N__29049),
            .I(N__29024));
    Span4Mux_v I__6401 (
            .O(N__29046),
            .I(N__29024));
    Span12Mux_h I__6400 (
            .O(N__29043),
            .I(N__29019));
    Sp12to4 I__6399 (
            .O(N__29040),
            .I(N__29019));
    Odrv4 I__6398 (
            .O(N__29037),
            .I(\tok.reset_N_2 ));
    Odrv4 I__6397 (
            .O(N__29034),
            .I(\tok.reset_N_2 ));
    Odrv4 I__6396 (
            .O(N__29029),
            .I(\tok.reset_N_2 ));
    Odrv4 I__6395 (
            .O(N__29024),
            .I(\tok.reset_N_2 ));
    Odrv12 I__6394 (
            .O(N__29019),
            .I(\tok.reset_N_2 ));
    InMux I__6393 (
            .O(N__29008),
            .I(N__29005));
    LocalMux I__6392 (
            .O(N__29005),
            .I(N__29002));
    Odrv4 I__6391 (
            .O(N__29002),
            .I(\tok.n256_adj_749 ));
    InMux I__6390 (
            .O(N__28999),
            .I(N__28996));
    LocalMux I__6389 (
            .O(N__28996),
            .I(\tok.n367 ));
    InMux I__6388 (
            .O(N__28993),
            .I(N__28990));
    LocalMux I__6387 (
            .O(N__28990),
            .I(N__28987));
    Span12Mux_s8_h I__6386 (
            .O(N__28987),
            .I(N__28984));
    Odrv12 I__6385 (
            .O(N__28984),
            .I(\tok.n215_adj_750 ));
    CascadeMux I__6384 (
            .O(N__28981),
            .I(N__28974));
    InMux I__6383 (
            .O(N__28980),
            .I(N__28966));
    InMux I__6382 (
            .O(N__28979),
            .I(N__28966));
    InMux I__6381 (
            .O(N__28978),
            .I(N__28959));
    InMux I__6380 (
            .O(N__28977),
            .I(N__28959));
    InMux I__6379 (
            .O(N__28974),
            .I(N__28959));
    InMux I__6378 (
            .O(N__28973),
            .I(N__28956));
    InMux I__6377 (
            .O(N__28972),
            .I(N__28953));
    InMux I__6376 (
            .O(N__28971),
            .I(N__28950));
    LocalMux I__6375 (
            .O(N__28966),
            .I(\tok.depth_2 ));
    LocalMux I__6374 (
            .O(N__28959),
            .I(\tok.depth_2 ));
    LocalMux I__6373 (
            .O(N__28956),
            .I(\tok.depth_2 ));
    LocalMux I__6372 (
            .O(N__28953),
            .I(\tok.depth_2 ));
    LocalMux I__6371 (
            .O(N__28950),
            .I(\tok.depth_2 ));
    InMux I__6370 (
            .O(N__28939),
            .I(N__28936));
    LocalMux I__6369 (
            .O(N__28936),
            .I(N__28932));
    InMux I__6368 (
            .O(N__28935),
            .I(N__28929));
    Span4Mux_h I__6367 (
            .O(N__28932),
            .I(N__28926));
    LocalMux I__6366 (
            .O(N__28929),
            .I(\tok.tail_47 ));
    Odrv4 I__6365 (
            .O(N__28926),
            .I(\tok.tail_47 ));
    CEMux I__6364 (
            .O(N__28921),
            .I(N__28914));
    CEMux I__6363 (
            .O(N__28920),
            .I(N__28911));
    CEMux I__6362 (
            .O(N__28919),
            .I(N__28906));
    CEMux I__6361 (
            .O(N__28918),
            .I(N__28902));
    CEMux I__6360 (
            .O(N__28917),
            .I(N__28899));
    LocalMux I__6359 (
            .O(N__28914),
            .I(N__28896));
    LocalMux I__6358 (
            .O(N__28911),
            .I(N__28893));
    CEMux I__6357 (
            .O(N__28910),
            .I(N__28890));
    CEMux I__6356 (
            .O(N__28909),
            .I(N__28886));
    LocalMux I__6355 (
            .O(N__28906),
            .I(N__28883));
    CEMux I__6354 (
            .O(N__28905),
            .I(N__28880));
    LocalMux I__6353 (
            .O(N__28902),
            .I(N__28877));
    LocalMux I__6352 (
            .O(N__28899),
            .I(N__28874));
    Span4Mux_h I__6351 (
            .O(N__28896),
            .I(N__28866));
    Span4Mux_s2_v I__6350 (
            .O(N__28893),
            .I(N__28866));
    LocalMux I__6349 (
            .O(N__28890),
            .I(N__28866));
    CEMux I__6348 (
            .O(N__28889),
            .I(N__28863));
    LocalMux I__6347 (
            .O(N__28886),
            .I(N__28859));
    Span4Mux_s2_v I__6346 (
            .O(N__28883),
            .I(N__28856));
    LocalMux I__6345 (
            .O(N__28880),
            .I(N__28853));
    Span4Mux_s2_v I__6344 (
            .O(N__28877),
            .I(N__28850));
    Span4Mux_v I__6343 (
            .O(N__28874),
            .I(N__28847));
    CEMux I__6342 (
            .O(N__28873),
            .I(N__28844));
    Span4Mux_s2_h I__6341 (
            .O(N__28866),
            .I(N__28839));
    LocalMux I__6340 (
            .O(N__28863),
            .I(N__28839));
    InMux I__6339 (
            .O(N__28862),
            .I(N__28836));
    Span4Mux_s2_v I__6338 (
            .O(N__28859),
            .I(N__28827));
    Span4Mux_h I__6337 (
            .O(N__28856),
            .I(N__28822));
    Span4Mux_s2_v I__6336 (
            .O(N__28853),
            .I(N__28822));
    Span4Mux_h I__6335 (
            .O(N__28850),
            .I(N__28817));
    Span4Mux_s0_h I__6334 (
            .O(N__28847),
            .I(N__28817));
    LocalMux I__6333 (
            .O(N__28844),
            .I(N__28812));
    Sp12to4 I__6332 (
            .O(N__28839),
            .I(N__28812));
    LocalMux I__6331 (
            .O(N__28836),
            .I(N__28809));
    InMux I__6330 (
            .O(N__28835),
            .I(N__28806));
    InMux I__6329 (
            .O(N__28834),
            .I(N__28795));
    InMux I__6328 (
            .O(N__28833),
            .I(N__28795));
    InMux I__6327 (
            .O(N__28832),
            .I(N__28795));
    InMux I__6326 (
            .O(N__28831),
            .I(N__28795));
    InMux I__6325 (
            .O(N__28830),
            .I(N__28795));
    Odrv4 I__6324 (
            .O(N__28827),
            .I(rd_7__N_373));
    Odrv4 I__6323 (
            .O(N__28822),
            .I(rd_7__N_373));
    Odrv4 I__6322 (
            .O(N__28817),
            .I(rd_7__N_373));
    Odrv12 I__6321 (
            .O(N__28812),
            .I(rd_7__N_373));
    Odrv4 I__6320 (
            .O(N__28809),
            .I(rd_7__N_373));
    LocalMux I__6319 (
            .O(N__28806),
            .I(rd_7__N_373));
    LocalMux I__6318 (
            .O(N__28795),
            .I(rd_7__N_373));
    CascadeMux I__6317 (
            .O(N__28780),
            .I(N__28777));
    InMux I__6316 (
            .O(N__28777),
            .I(N__28773));
    InMux I__6315 (
            .O(N__28776),
            .I(N__28770));
    LocalMux I__6314 (
            .O(N__28773),
            .I(N__28767));
    LocalMux I__6313 (
            .O(N__28770),
            .I(N__28764));
    Span4Mux_s2_h I__6312 (
            .O(N__28767),
            .I(N__28761));
    Span4Mux_s1_h I__6311 (
            .O(N__28764),
            .I(N__28758));
    Odrv4 I__6310 (
            .O(N__28761),
            .I(\tok.tail_55 ));
    Odrv4 I__6309 (
            .O(N__28758),
            .I(\tok.tail_55 ));
    InMux I__6308 (
            .O(N__28753),
            .I(N__28720));
    InMux I__6307 (
            .O(N__28752),
            .I(N__28720));
    InMux I__6306 (
            .O(N__28751),
            .I(N__28720));
    InMux I__6305 (
            .O(N__28750),
            .I(N__28720));
    InMux I__6304 (
            .O(N__28749),
            .I(N__28720));
    InMux I__6303 (
            .O(N__28748),
            .I(N__28720));
    InMux I__6302 (
            .O(N__28747),
            .I(N__28707));
    InMux I__6301 (
            .O(N__28746),
            .I(N__28707));
    InMux I__6300 (
            .O(N__28745),
            .I(N__28707));
    InMux I__6299 (
            .O(N__28744),
            .I(N__28707));
    InMux I__6298 (
            .O(N__28743),
            .I(N__28707));
    InMux I__6297 (
            .O(N__28742),
            .I(N__28707));
    InMux I__6296 (
            .O(N__28741),
            .I(N__28694));
    InMux I__6295 (
            .O(N__28740),
            .I(N__28694));
    InMux I__6294 (
            .O(N__28739),
            .I(N__28694));
    InMux I__6293 (
            .O(N__28738),
            .I(N__28694));
    InMux I__6292 (
            .O(N__28737),
            .I(N__28694));
    InMux I__6291 (
            .O(N__28736),
            .I(N__28694));
    InMux I__6290 (
            .O(N__28735),
            .I(N__28686));
    InMux I__6289 (
            .O(N__28734),
            .I(N__28681));
    InMux I__6288 (
            .O(N__28733),
            .I(N__28681));
    LocalMux I__6287 (
            .O(N__28720),
            .I(N__28671));
    LocalMux I__6286 (
            .O(N__28707),
            .I(N__28666));
    LocalMux I__6285 (
            .O(N__28694),
            .I(N__28666));
    InMux I__6284 (
            .O(N__28693),
            .I(N__28649));
    InMux I__6283 (
            .O(N__28692),
            .I(N__28649));
    InMux I__6282 (
            .O(N__28691),
            .I(N__28649));
    InMux I__6281 (
            .O(N__28690),
            .I(N__28649));
    InMux I__6280 (
            .O(N__28689),
            .I(N__28649));
    LocalMux I__6279 (
            .O(N__28686),
            .I(N__28646));
    LocalMux I__6278 (
            .O(N__28681),
            .I(N__28643));
    InMux I__6277 (
            .O(N__28680),
            .I(N__28630));
    InMux I__6276 (
            .O(N__28679),
            .I(N__28630));
    InMux I__6275 (
            .O(N__28678),
            .I(N__28630));
    InMux I__6274 (
            .O(N__28677),
            .I(N__28630));
    InMux I__6273 (
            .O(N__28676),
            .I(N__28630));
    InMux I__6272 (
            .O(N__28675),
            .I(N__28630));
    InMux I__6271 (
            .O(N__28674),
            .I(N__28603));
    Span4Mux_s2_v I__6270 (
            .O(N__28671),
            .I(N__28600));
    Span4Mux_h I__6269 (
            .O(N__28666),
            .I(N__28597));
    InMux I__6268 (
            .O(N__28665),
            .I(N__28584));
    InMux I__6267 (
            .O(N__28664),
            .I(N__28584));
    InMux I__6266 (
            .O(N__28663),
            .I(N__28584));
    InMux I__6265 (
            .O(N__28662),
            .I(N__28584));
    InMux I__6264 (
            .O(N__28661),
            .I(N__28584));
    InMux I__6263 (
            .O(N__28660),
            .I(N__28584));
    LocalMux I__6262 (
            .O(N__28649),
            .I(N__28581));
    Span4Mux_v I__6261 (
            .O(N__28646),
            .I(N__28574));
    Span4Mux_s2_v I__6260 (
            .O(N__28643),
            .I(N__28574));
    LocalMux I__6259 (
            .O(N__28630),
            .I(N__28574));
    InMux I__6258 (
            .O(N__28629),
            .I(N__28559));
    InMux I__6257 (
            .O(N__28628),
            .I(N__28559));
    InMux I__6256 (
            .O(N__28627),
            .I(N__28559));
    InMux I__6255 (
            .O(N__28626),
            .I(N__28559));
    InMux I__6254 (
            .O(N__28625),
            .I(N__28559));
    InMux I__6253 (
            .O(N__28624),
            .I(N__28559));
    InMux I__6252 (
            .O(N__28623),
            .I(N__28559));
    InMux I__6251 (
            .O(N__28622),
            .I(N__28546));
    InMux I__6250 (
            .O(N__28621),
            .I(N__28546));
    InMux I__6249 (
            .O(N__28620),
            .I(N__28546));
    InMux I__6248 (
            .O(N__28619),
            .I(N__28546));
    InMux I__6247 (
            .O(N__28618),
            .I(N__28546));
    InMux I__6246 (
            .O(N__28617),
            .I(N__28546));
    InMux I__6245 (
            .O(N__28616),
            .I(N__28533));
    InMux I__6244 (
            .O(N__28615),
            .I(N__28533));
    InMux I__6243 (
            .O(N__28614),
            .I(N__28533));
    InMux I__6242 (
            .O(N__28613),
            .I(N__28533));
    InMux I__6241 (
            .O(N__28612),
            .I(N__28533));
    InMux I__6240 (
            .O(N__28611),
            .I(N__28533));
    InMux I__6239 (
            .O(N__28610),
            .I(N__28522));
    InMux I__6238 (
            .O(N__28609),
            .I(N__28522));
    InMux I__6237 (
            .O(N__28608),
            .I(N__28522));
    InMux I__6236 (
            .O(N__28607),
            .I(N__28522));
    InMux I__6235 (
            .O(N__28606),
            .I(N__28522));
    LocalMux I__6234 (
            .O(N__28603),
            .I(C_stk_delta_1));
    Odrv4 I__6233 (
            .O(N__28600),
            .I(C_stk_delta_1));
    Odrv4 I__6232 (
            .O(N__28597),
            .I(C_stk_delta_1));
    LocalMux I__6231 (
            .O(N__28584),
            .I(C_stk_delta_1));
    Odrv4 I__6230 (
            .O(N__28581),
            .I(C_stk_delta_1));
    Odrv4 I__6229 (
            .O(N__28574),
            .I(C_stk_delta_1));
    LocalMux I__6228 (
            .O(N__28559),
            .I(C_stk_delta_1));
    LocalMux I__6227 (
            .O(N__28546),
            .I(C_stk_delta_1));
    LocalMux I__6226 (
            .O(N__28533),
            .I(C_stk_delta_1));
    LocalMux I__6225 (
            .O(N__28522),
            .I(C_stk_delta_1));
    InMux I__6224 (
            .O(N__28501),
            .I(N__28498));
    LocalMux I__6223 (
            .O(N__28498),
            .I(N__28495));
    Span4Mux_s1_v I__6222 (
            .O(N__28495),
            .I(N__28491));
    InMux I__6221 (
            .O(N__28494),
            .I(N__28488));
    Odrv4 I__6220 (
            .O(N__28491),
            .I(\tok.tail_63 ));
    LocalMux I__6219 (
            .O(N__28488),
            .I(\tok.tail_63 ));
    InMux I__6218 (
            .O(N__28483),
            .I(N__28480));
    LocalMux I__6217 (
            .O(N__28480),
            .I(N__28469));
    InMux I__6216 (
            .O(N__28479),
            .I(N__28458));
    InMux I__6215 (
            .O(N__28478),
            .I(N__28458));
    InMux I__6214 (
            .O(N__28477),
            .I(N__28458));
    InMux I__6213 (
            .O(N__28476),
            .I(N__28458));
    InMux I__6212 (
            .O(N__28475),
            .I(N__28458));
    InMux I__6211 (
            .O(N__28474),
            .I(N__28455));
    CascadeMux I__6210 (
            .O(N__28473),
            .I(N__28452));
    InMux I__6209 (
            .O(N__28472),
            .I(N__28444));
    Span4Mux_h I__6208 (
            .O(N__28469),
            .I(N__28441));
    LocalMux I__6207 (
            .O(N__28458),
            .I(N__28438));
    LocalMux I__6206 (
            .O(N__28455),
            .I(N__28435));
    InMux I__6205 (
            .O(N__28452),
            .I(N__28426));
    InMux I__6204 (
            .O(N__28451),
            .I(N__28426));
    InMux I__6203 (
            .O(N__28450),
            .I(N__28426));
    InMux I__6202 (
            .O(N__28449),
            .I(N__28426));
    InMux I__6201 (
            .O(N__28448),
            .I(N__28419));
    InMux I__6200 (
            .O(N__28447),
            .I(N__28419));
    LocalMux I__6199 (
            .O(N__28444),
            .I(N__28416));
    Sp12to4 I__6198 (
            .O(N__28441),
            .I(N__28413));
    Span4Mux_s3_v I__6197 (
            .O(N__28438),
            .I(N__28410));
    Span4Mux_v I__6196 (
            .O(N__28435),
            .I(N__28405));
    LocalMux I__6195 (
            .O(N__28426),
            .I(N__28405));
    InMux I__6194 (
            .O(N__28425),
            .I(N__28402));
    InMux I__6193 (
            .O(N__28424),
            .I(N__28399));
    LocalMux I__6192 (
            .O(N__28419),
            .I(N__28396));
    Odrv12 I__6191 (
            .O(N__28416),
            .I(n15));
    Odrv12 I__6190 (
            .O(N__28413),
            .I(n15));
    Odrv4 I__6189 (
            .O(N__28410),
            .I(n15));
    Odrv4 I__6188 (
            .O(N__28405),
            .I(n15));
    LocalMux I__6187 (
            .O(N__28402),
            .I(n15));
    LocalMux I__6186 (
            .O(N__28399),
            .I(n15));
    Odrv4 I__6185 (
            .O(N__28396),
            .I(n15));
    InMux I__6184 (
            .O(N__28381),
            .I(N__28377));
    InMux I__6183 (
            .O(N__28380),
            .I(N__28374));
    LocalMux I__6182 (
            .O(N__28377),
            .I(N__28370));
    LocalMux I__6181 (
            .O(N__28374),
            .I(N__28367));
    CascadeMux I__6180 (
            .O(N__28373),
            .I(N__28364));
    Span4Mux_s3_h I__6179 (
            .O(N__28370),
            .I(N__28360));
    Span4Mux_s2_h I__6178 (
            .O(N__28367),
            .I(N__28357));
    InMux I__6177 (
            .O(N__28364),
            .I(N__28352));
    InMux I__6176 (
            .O(N__28363),
            .I(N__28352));
    Span4Mux_h I__6175 (
            .O(N__28360),
            .I(N__28349));
    Span4Mux_h I__6174 (
            .O(N__28357),
            .I(N__28344));
    LocalMux I__6173 (
            .O(N__28352),
            .I(N__28344));
    Odrv4 I__6172 (
            .O(N__28349),
            .I(\tok.tc_plus_1_7 ));
    Odrv4 I__6171 (
            .O(N__28344),
            .I(\tok.tc_plus_1_7 ));
    InMux I__6170 (
            .O(N__28339),
            .I(N__28335));
    InMux I__6169 (
            .O(N__28338),
            .I(N__28331));
    LocalMux I__6168 (
            .O(N__28335),
            .I(N__28325));
    InMux I__6167 (
            .O(N__28334),
            .I(N__28322));
    LocalMux I__6166 (
            .O(N__28331),
            .I(N__28319));
    CascadeMux I__6165 (
            .O(N__28330),
            .I(N__28316));
    InMux I__6164 (
            .O(N__28329),
            .I(N__28313));
    InMux I__6163 (
            .O(N__28328),
            .I(N__28310));
    Span4Mux_v I__6162 (
            .O(N__28325),
            .I(N__28307));
    LocalMux I__6161 (
            .O(N__28322),
            .I(N__28302));
    Span4Mux_h I__6160 (
            .O(N__28319),
            .I(N__28302));
    InMux I__6159 (
            .O(N__28316),
            .I(N__28299));
    LocalMux I__6158 (
            .O(N__28313),
            .I(N__28294));
    LocalMux I__6157 (
            .O(N__28310),
            .I(N__28291));
    Span4Mux_h I__6156 (
            .O(N__28307),
            .I(N__28286));
    Span4Mux_v I__6155 (
            .O(N__28302),
            .I(N__28286));
    LocalMux I__6154 (
            .O(N__28299),
            .I(N__28283));
    InMux I__6153 (
            .O(N__28298),
            .I(N__28280));
    InMux I__6152 (
            .O(N__28297),
            .I(N__28277));
    Span4Mux_v I__6151 (
            .O(N__28294),
            .I(N__28274));
    Span4Mux_v I__6150 (
            .O(N__28291),
            .I(N__28271));
    Span4Mux_h I__6149 (
            .O(N__28286),
            .I(N__28266));
    Span4Mux_v I__6148 (
            .O(N__28283),
            .I(N__28266));
    LocalMux I__6147 (
            .O(N__28280),
            .I(N__28263));
    LocalMux I__6146 (
            .O(N__28277),
            .I(N__28258));
    Span4Mux_v I__6145 (
            .O(N__28274),
            .I(N__28258));
    Span4Mux_v I__6144 (
            .O(N__28271),
            .I(N__28253));
    Span4Mux_v I__6143 (
            .O(N__28266),
            .I(N__28253));
    Span12Mux_v I__6142 (
            .O(N__28263),
            .I(N__28250));
    Odrv4 I__6141 (
            .O(N__28258),
            .I(\tok.S_7 ));
    Odrv4 I__6140 (
            .O(N__28253),
            .I(\tok.S_7 ));
    Odrv12 I__6139 (
            .O(N__28250),
            .I(\tok.S_7 ));
    InMux I__6138 (
            .O(N__28243),
            .I(N__28240));
    LocalMux I__6137 (
            .O(N__28240),
            .I(N__28237));
    Span4Mux_v I__6136 (
            .O(N__28237),
            .I(N__28234));
    Sp12to4 I__6135 (
            .O(N__28234),
            .I(N__28231));
    Span12Mux_h I__6134 (
            .O(N__28231),
            .I(N__28228));
    Odrv12 I__6133 (
            .O(N__28228),
            .I(\tok.table_wr_data_7 ));
    InMux I__6132 (
            .O(N__28225),
            .I(N__28222));
    LocalMux I__6131 (
            .O(N__28222),
            .I(N__28218));
    InMux I__6130 (
            .O(N__28221),
            .I(N__28215));
    Span4Mux_h I__6129 (
            .O(N__28218),
            .I(N__28212));
    LocalMux I__6128 (
            .O(N__28215),
            .I(uart_rx_data_4));
    Odrv4 I__6127 (
            .O(N__28212),
            .I(uart_rx_data_4));
    InMux I__6126 (
            .O(N__28207),
            .I(N__28204));
    LocalMux I__6125 (
            .O(N__28204),
            .I(N__28200));
    InMux I__6124 (
            .O(N__28203),
            .I(N__28197));
    Span4Mux_h I__6123 (
            .O(N__28200),
            .I(N__28194));
    LocalMux I__6122 (
            .O(N__28197),
            .I(uart_rx_data_2));
    Odrv4 I__6121 (
            .O(N__28194),
            .I(uart_rx_data_2));
    InMux I__6120 (
            .O(N__28189),
            .I(N__28185));
    InMux I__6119 (
            .O(N__28188),
            .I(N__28182));
    LocalMux I__6118 (
            .O(N__28185),
            .I(N__28179));
    LocalMux I__6117 (
            .O(N__28182),
            .I(uart_rx_data_1));
    Odrv4 I__6116 (
            .O(N__28179),
            .I(uart_rx_data_1));
    InMux I__6115 (
            .O(N__28174),
            .I(N__28169));
    InMux I__6114 (
            .O(N__28173),
            .I(N__28164));
    InMux I__6113 (
            .O(N__28172),
            .I(N__28164));
    LocalMux I__6112 (
            .O(N__28169),
            .I(capture_2));
    LocalMux I__6111 (
            .O(N__28164),
            .I(capture_2));
    CascadeMux I__6110 (
            .O(N__28159),
            .I(N__28155));
    InMux I__6109 (
            .O(N__28158),
            .I(N__28152));
    InMux I__6108 (
            .O(N__28155),
            .I(N__28149));
    LocalMux I__6107 (
            .O(N__28152),
            .I(\tok.tail_54 ));
    LocalMux I__6106 (
            .O(N__28149),
            .I(\tok.tail_54 ));
    InMux I__6105 (
            .O(N__28144),
            .I(N__28138));
    InMux I__6104 (
            .O(N__28143),
            .I(N__28138));
    LocalMux I__6103 (
            .O(N__28138),
            .I(\tok.C_stk.tail_38 ));
    InMux I__6102 (
            .O(N__28135),
            .I(N__28131));
    InMux I__6101 (
            .O(N__28134),
            .I(N__28128));
    LocalMux I__6100 (
            .O(N__28131),
            .I(\tok.tail_46 ));
    LocalMux I__6099 (
            .O(N__28128),
            .I(\tok.tail_46 ));
    InMux I__6098 (
            .O(N__28123),
            .I(N__28119));
    InMux I__6097 (
            .O(N__28122),
            .I(N__28113));
    LocalMux I__6096 (
            .O(N__28119),
            .I(N__28110));
    InMux I__6095 (
            .O(N__28118),
            .I(N__28107));
    InMux I__6094 (
            .O(N__28117),
            .I(N__28104));
    InMux I__6093 (
            .O(N__28116),
            .I(N__28099));
    LocalMux I__6092 (
            .O(N__28113),
            .I(N__28095));
    Span4Mux_s3_v I__6091 (
            .O(N__28110),
            .I(N__28088));
    LocalMux I__6090 (
            .O(N__28107),
            .I(N__28088));
    LocalMux I__6089 (
            .O(N__28104),
            .I(N__28088));
    InMux I__6088 (
            .O(N__28103),
            .I(N__28085));
    InMux I__6087 (
            .O(N__28102),
            .I(N__28082));
    LocalMux I__6086 (
            .O(N__28099),
            .I(N__28079));
    InMux I__6085 (
            .O(N__28098),
            .I(N__28076));
    Span4Mux_s3_v I__6084 (
            .O(N__28095),
            .I(N__28071));
    Span4Mux_h I__6083 (
            .O(N__28088),
            .I(N__28071));
    LocalMux I__6082 (
            .O(N__28085),
            .I(N__28066));
    LocalMux I__6081 (
            .O(N__28082),
            .I(N__28066));
    Span4Mux_s0_v I__6080 (
            .O(N__28079),
            .I(N__28061));
    LocalMux I__6079 (
            .O(N__28076),
            .I(N__28061));
    Odrv4 I__6078 (
            .O(N__28071),
            .I(\tok.C_stk.n449 ));
    Odrv4 I__6077 (
            .O(N__28066),
            .I(\tok.C_stk.n449 ));
    Odrv4 I__6076 (
            .O(N__28061),
            .I(\tok.C_stk.n449 ));
    InMux I__6075 (
            .O(N__28054),
            .I(N__28044));
    InMux I__6074 (
            .O(N__28053),
            .I(N__28041));
    InMux I__6073 (
            .O(N__28052),
            .I(N__28038));
    InMux I__6072 (
            .O(N__28051),
            .I(N__28035));
    InMux I__6071 (
            .O(N__28050),
            .I(N__28032));
    InMux I__6070 (
            .O(N__28049),
            .I(N__28029));
    InMux I__6069 (
            .O(N__28048),
            .I(N__28026));
    InMux I__6068 (
            .O(N__28047),
            .I(N__28023));
    LocalMux I__6067 (
            .O(N__28044),
            .I(N__28020));
    LocalMux I__6066 (
            .O(N__28041),
            .I(N__28015));
    LocalMux I__6065 (
            .O(N__28038),
            .I(N__28015));
    LocalMux I__6064 (
            .O(N__28035),
            .I(N__28010));
    LocalMux I__6063 (
            .O(N__28032),
            .I(N__28010));
    LocalMux I__6062 (
            .O(N__28029),
            .I(N__28005));
    LocalMux I__6061 (
            .O(N__28026),
            .I(N__28005));
    LocalMux I__6060 (
            .O(N__28023),
            .I(N__28001));
    Span4Mux_s3_v I__6059 (
            .O(N__28020),
            .I(N__27996));
    Span4Mux_h I__6058 (
            .O(N__28015),
            .I(N__27996));
    Span4Mux_s2_v I__6057 (
            .O(N__28010),
            .I(N__27991));
    Span4Mux_h I__6056 (
            .O(N__28005),
            .I(N__27991));
    InMux I__6055 (
            .O(N__28004),
            .I(N__27988));
    Odrv12 I__6054 (
            .O(N__28001),
            .I(\tok.n273 ));
    Odrv4 I__6053 (
            .O(N__27996),
            .I(\tok.n273 ));
    Odrv4 I__6052 (
            .O(N__27991),
            .I(\tok.n273 ));
    LocalMux I__6051 (
            .O(N__27988),
            .I(\tok.n273 ));
    InMux I__6050 (
            .O(N__27979),
            .I(N__27974));
    InMux I__6049 (
            .O(N__27978),
            .I(N__27971));
    InMux I__6048 (
            .O(N__27977),
            .I(N__27967));
    LocalMux I__6047 (
            .O(N__27974),
            .I(N__27964));
    LocalMux I__6046 (
            .O(N__27971),
            .I(N__27961));
    InMux I__6045 (
            .O(N__27970),
            .I(N__27958));
    LocalMux I__6044 (
            .O(N__27967),
            .I(N__27955));
    Odrv4 I__6043 (
            .O(N__27964),
            .I(tc_7));
    Odrv12 I__6042 (
            .O(N__27961),
            .I(tc_7));
    LocalMux I__6041 (
            .O(N__27958),
            .I(tc_7));
    Odrv4 I__6040 (
            .O(N__27955),
            .I(tc_7));
    CascadeMux I__6039 (
            .O(N__27946),
            .I(\tok.C_stk.n6227_cascade_ ));
    InMux I__6038 (
            .O(N__27943),
            .I(N__27937));
    InMux I__6037 (
            .O(N__27942),
            .I(N__27934));
    InMux I__6036 (
            .O(N__27941),
            .I(N__27930));
    InMux I__6035 (
            .O(N__27940),
            .I(N__27926));
    LocalMux I__6034 (
            .O(N__27937),
            .I(N__27918));
    LocalMux I__6033 (
            .O(N__27934),
            .I(N__27918));
    InMux I__6032 (
            .O(N__27933),
            .I(N__27915));
    LocalMux I__6031 (
            .O(N__27930),
            .I(N__27912));
    InMux I__6030 (
            .O(N__27929),
            .I(N__27909));
    LocalMux I__6029 (
            .O(N__27926),
            .I(N__27906));
    InMux I__6028 (
            .O(N__27925),
            .I(N__27903));
    InMux I__6027 (
            .O(N__27924),
            .I(N__27900));
    InMux I__6026 (
            .O(N__27923),
            .I(N__27897));
    Span4Mux_v I__6025 (
            .O(N__27918),
            .I(N__27894));
    LocalMux I__6024 (
            .O(N__27915),
            .I(N__27891));
    Span4Mux_v I__6023 (
            .O(N__27912),
            .I(N__27888));
    LocalMux I__6022 (
            .O(N__27909),
            .I(N__27885));
    Span4Mux_s1_v I__6021 (
            .O(N__27906),
            .I(N__27880));
    LocalMux I__6020 (
            .O(N__27903),
            .I(N__27880));
    LocalMux I__6019 (
            .O(N__27900),
            .I(N__27877));
    LocalMux I__6018 (
            .O(N__27897),
            .I(N__27874));
    Odrv4 I__6017 (
            .O(N__27894),
            .I(\tok.n15 ));
    Odrv4 I__6016 (
            .O(N__27891),
            .I(\tok.n15 ));
    Odrv4 I__6015 (
            .O(N__27888),
            .I(\tok.n15 ));
    Odrv12 I__6014 (
            .O(N__27885),
            .I(\tok.n15 ));
    Odrv4 I__6013 (
            .O(N__27880),
            .I(\tok.n15 ));
    Odrv4 I__6012 (
            .O(N__27877),
            .I(\tok.n15 ));
    Odrv12 I__6011 (
            .O(N__27874),
            .I(\tok.n15 ));
    CascadeMux I__6010 (
            .O(N__27859),
            .I(N__27855));
    InMux I__6009 (
            .O(N__27858),
            .I(N__27846));
    InMux I__6008 (
            .O(N__27855),
            .I(N__27846));
    InMux I__6007 (
            .O(N__27854),
            .I(N__27846));
    InMux I__6006 (
            .O(N__27853),
            .I(N__27843));
    LocalMux I__6005 (
            .O(N__27846),
            .I(N__27840));
    LocalMux I__6004 (
            .O(N__27843),
            .I(\tok.c_stk_r_7 ));
    Odrv12 I__6003 (
            .O(N__27840),
            .I(\tok.c_stk_r_7 ));
    InMux I__6002 (
            .O(N__27835),
            .I(N__27829));
    InMux I__6001 (
            .O(N__27834),
            .I(N__27829));
    LocalMux I__6000 (
            .O(N__27829),
            .I(\tok.C_stk.tail_7 ));
    InMux I__5999 (
            .O(N__27826),
            .I(N__27820));
    InMux I__5998 (
            .O(N__27825),
            .I(N__27820));
    LocalMux I__5997 (
            .O(N__27820),
            .I(\tok.tail_15 ));
    CascadeMux I__5996 (
            .O(N__27817),
            .I(N__27814));
    InMux I__5995 (
            .O(N__27814),
            .I(N__27808));
    InMux I__5994 (
            .O(N__27813),
            .I(N__27808));
    LocalMux I__5993 (
            .O(N__27808),
            .I(\tok.C_stk.tail_23 ));
    InMux I__5992 (
            .O(N__27805),
            .I(N__27799));
    InMux I__5991 (
            .O(N__27804),
            .I(N__27799));
    LocalMux I__5990 (
            .O(N__27799),
            .I(\tok.tail_31 ));
    InMux I__5989 (
            .O(N__27796),
            .I(N__27790));
    InMux I__5988 (
            .O(N__27795),
            .I(N__27790));
    LocalMux I__5987 (
            .O(N__27790),
            .I(\tok.C_stk.tail_39 ));
    InMux I__5986 (
            .O(N__27787),
            .I(N__27784));
    LocalMux I__5985 (
            .O(N__27784),
            .I(reset_c));
    InMux I__5984 (
            .O(N__27781),
            .I(N__27778));
    LocalMux I__5983 (
            .O(N__27778),
            .I(N__27774));
    CascadeMux I__5982 (
            .O(N__27777),
            .I(N__27771));
    Span4Mux_h I__5981 (
            .O(N__27774),
            .I(N__27768));
    InMux I__5980 (
            .O(N__27771),
            .I(N__27765));
    Odrv4 I__5979 (
            .O(N__27768),
            .I(\tok.tail_50 ));
    LocalMux I__5978 (
            .O(N__27765),
            .I(\tok.tail_50 ));
    InMux I__5977 (
            .O(N__27760),
            .I(N__27756));
    InMux I__5976 (
            .O(N__27759),
            .I(N__27753));
    LocalMux I__5975 (
            .O(N__27756),
            .I(\tok.tail_58 ));
    LocalMux I__5974 (
            .O(N__27753),
            .I(\tok.tail_58 ));
    InMux I__5973 (
            .O(N__27748),
            .I(N__27745));
    LocalMux I__5972 (
            .O(N__27745),
            .I(N__27742));
    Span4Mux_s2_h I__5971 (
            .O(N__27742),
            .I(N__27739));
    Span4Mux_h I__5970 (
            .O(N__27739),
            .I(N__27733));
    InMux I__5969 (
            .O(N__27738),
            .I(N__27730));
    InMux I__5968 (
            .O(N__27737),
            .I(N__27725));
    InMux I__5967 (
            .O(N__27736),
            .I(N__27725));
    Odrv4 I__5966 (
            .O(N__27733),
            .I(\tok.tc_plus_1_6 ));
    LocalMux I__5965 (
            .O(N__27730),
            .I(\tok.tc_plus_1_6 ));
    LocalMux I__5964 (
            .O(N__27725),
            .I(\tok.tc_plus_1_6 ));
    CascadeMux I__5963 (
            .O(N__27718),
            .I(\tok.C_stk.n6233_cascade_ ));
    InMux I__5962 (
            .O(N__27715),
            .I(N__27712));
    LocalMux I__5961 (
            .O(N__27712),
            .I(N__27708));
    CascadeMux I__5960 (
            .O(N__27711),
            .I(N__27703));
    Span4Mux_h I__5959 (
            .O(N__27708),
            .I(N__27700));
    InMux I__5958 (
            .O(N__27707),
            .I(N__27695));
    InMux I__5957 (
            .O(N__27706),
            .I(N__27695));
    InMux I__5956 (
            .O(N__27703),
            .I(N__27692));
    Odrv4 I__5955 (
            .O(N__27700),
            .I(tc_6));
    LocalMux I__5954 (
            .O(N__27695),
            .I(tc_6));
    LocalMux I__5953 (
            .O(N__27692),
            .I(tc_6));
    CascadeMux I__5952 (
            .O(N__27685),
            .I(N__27681));
    InMux I__5951 (
            .O(N__27684),
            .I(N__27673));
    InMux I__5950 (
            .O(N__27681),
            .I(N__27673));
    InMux I__5949 (
            .O(N__27680),
            .I(N__27673));
    LocalMux I__5948 (
            .O(N__27673),
            .I(N__27669));
    InMux I__5947 (
            .O(N__27672),
            .I(N__27666));
    Span4Mux_h I__5946 (
            .O(N__27669),
            .I(N__27663));
    LocalMux I__5945 (
            .O(N__27666),
            .I(\tok.c_stk_r_6 ));
    Odrv4 I__5944 (
            .O(N__27663),
            .I(\tok.c_stk_r_6 ));
    InMux I__5943 (
            .O(N__27658),
            .I(N__27652));
    InMux I__5942 (
            .O(N__27657),
            .I(N__27652));
    LocalMux I__5941 (
            .O(N__27652),
            .I(\tok.C_stk.tail_6 ));
    InMux I__5940 (
            .O(N__27649),
            .I(N__27643));
    InMux I__5939 (
            .O(N__27648),
            .I(N__27643));
    LocalMux I__5938 (
            .O(N__27643),
            .I(\tok.tail_14 ));
    CascadeMux I__5937 (
            .O(N__27640),
            .I(N__27637));
    InMux I__5936 (
            .O(N__27637),
            .I(N__27631));
    InMux I__5935 (
            .O(N__27636),
            .I(N__27631));
    LocalMux I__5934 (
            .O(N__27631),
            .I(\tok.C_stk.tail_22 ));
    InMux I__5933 (
            .O(N__27628),
            .I(N__27622));
    InMux I__5932 (
            .O(N__27627),
            .I(N__27622));
    LocalMux I__5931 (
            .O(N__27622),
            .I(\tok.tail_30 ));
    InMux I__5930 (
            .O(N__27619),
            .I(N__27616));
    LocalMux I__5929 (
            .O(N__27616),
            .I(\tok.n6641 ));
    CascadeMux I__5928 (
            .O(N__27613),
            .I(\tok.n266_cascade_ ));
    InMux I__5927 (
            .O(N__27610),
            .I(N__27604));
    InMux I__5926 (
            .O(N__27609),
            .I(N__27604));
    LocalMux I__5925 (
            .O(N__27604),
            .I(N__27601));
    Span4Mux_v I__5924 (
            .O(N__27601),
            .I(N__27598));
    Sp12to4 I__5923 (
            .O(N__27598),
            .I(N__27595));
    Odrv12 I__5922 (
            .O(N__27595),
            .I(\tok.n5_adj_713 ));
    InMux I__5921 (
            .O(N__27592),
            .I(N__27589));
    LocalMux I__5920 (
            .O(N__27589),
            .I(N__27586));
    Span4Mux_h I__5919 (
            .O(N__27586),
            .I(N__27583));
    Odrv4 I__5918 (
            .O(N__27583),
            .I(\tok.n256 ));
    CascadeMux I__5917 (
            .O(N__27580),
            .I(\tok.n4_adj_718_cascade_ ));
    InMux I__5916 (
            .O(N__27577),
            .I(N__27574));
    LocalMux I__5915 (
            .O(N__27574),
            .I(N__27571));
    Span4Mux_h I__5914 (
            .O(N__27571),
            .I(N__27568));
    Span4Mux_v I__5913 (
            .O(N__27568),
            .I(N__27565));
    Odrv4 I__5912 (
            .O(N__27565),
            .I(\tok.n221 ));
    InMux I__5911 (
            .O(N__27562),
            .I(N__27555));
    CascadeMux I__5910 (
            .O(N__27561),
            .I(N__27548));
    InMux I__5909 (
            .O(N__27560),
            .I(N__27545));
    CascadeMux I__5908 (
            .O(N__27559),
            .I(N__27537));
    CascadeMux I__5907 (
            .O(N__27558),
            .I(N__27533));
    LocalMux I__5906 (
            .O(N__27555),
            .I(N__27530));
    InMux I__5905 (
            .O(N__27554),
            .I(N__27525));
    InMux I__5904 (
            .O(N__27553),
            .I(N__27525));
    InMux I__5903 (
            .O(N__27552),
            .I(N__27520));
    InMux I__5902 (
            .O(N__27551),
            .I(N__27515));
    InMux I__5901 (
            .O(N__27548),
            .I(N__27515));
    LocalMux I__5900 (
            .O(N__27545),
            .I(N__27511));
    InMux I__5899 (
            .O(N__27544),
            .I(N__27506));
    InMux I__5898 (
            .O(N__27543),
            .I(N__27501));
    InMux I__5897 (
            .O(N__27542),
            .I(N__27501));
    InMux I__5896 (
            .O(N__27541),
            .I(N__27498));
    InMux I__5895 (
            .O(N__27540),
            .I(N__27493));
    InMux I__5894 (
            .O(N__27537),
            .I(N__27493));
    InMux I__5893 (
            .O(N__27536),
            .I(N__27490));
    InMux I__5892 (
            .O(N__27533),
            .I(N__27487));
    Span4Mux_s3_v I__5891 (
            .O(N__27530),
            .I(N__27482));
    LocalMux I__5890 (
            .O(N__27525),
            .I(N__27482));
    InMux I__5889 (
            .O(N__27524),
            .I(N__27477));
    InMux I__5888 (
            .O(N__27523),
            .I(N__27477));
    LocalMux I__5887 (
            .O(N__27520),
            .I(N__27472));
    LocalMux I__5886 (
            .O(N__27515),
            .I(N__27472));
    InMux I__5885 (
            .O(N__27514),
            .I(N__27468));
    Sp12to4 I__5884 (
            .O(N__27511),
            .I(N__27465));
    InMux I__5883 (
            .O(N__27510),
            .I(N__27462));
    CascadeMux I__5882 (
            .O(N__27509),
            .I(N__27458));
    LocalMux I__5881 (
            .O(N__27506),
            .I(N__27452));
    LocalMux I__5880 (
            .O(N__27501),
            .I(N__27452));
    LocalMux I__5879 (
            .O(N__27498),
            .I(N__27449));
    LocalMux I__5878 (
            .O(N__27493),
            .I(N__27442));
    LocalMux I__5877 (
            .O(N__27490),
            .I(N__27442));
    LocalMux I__5876 (
            .O(N__27487),
            .I(N__27442));
    Span4Mux_v I__5875 (
            .O(N__27482),
            .I(N__27435));
    LocalMux I__5874 (
            .O(N__27477),
            .I(N__27435));
    Span4Mux_v I__5873 (
            .O(N__27472),
            .I(N__27435));
    InMux I__5872 (
            .O(N__27471),
            .I(N__27432));
    LocalMux I__5871 (
            .O(N__27468),
            .I(N__27425));
    Span12Mux_s6_v I__5870 (
            .O(N__27465),
            .I(N__27425));
    LocalMux I__5869 (
            .O(N__27462),
            .I(N__27425));
    InMux I__5868 (
            .O(N__27461),
            .I(N__27418));
    InMux I__5867 (
            .O(N__27458),
            .I(N__27418));
    InMux I__5866 (
            .O(N__27457),
            .I(N__27418));
    Span4Mux_v I__5865 (
            .O(N__27452),
            .I(N__27409));
    Span4Mux_v I__5864 (
            .O(N__27449),
            .I(N__27409));
    Span4Mux_v I__5863 (
            .O(N__27442),
            .I(N__27409));
    Span4Mux_h I__5862 (
            .O(N__27435),
            .I(N__27409));
    LocalMux I__5861 (
            .O(N__27432),
            .I(\tok.A_low_1 ));
    Odrv12 I__5860 (
            .O(N__27425),
            .I(\tok.A_low_1 ));
    LocalMux I__5859 (
            .O(N__27418),
            .I(\tok.A_low_1 ));
    Odrv4 I__5858 (
            .O(N__27409),
            .I(\tok.A_low_1 ));
    InMux I__5857 (
            .O(N__27400),
            .I(N__27397));
    LocalMux I__5856 (
            .O(N__27397),
            .I(\tok.n2637 ));
    CascadeMux I__5855 (
            .O(N__27394),
            .I(N__27383));
    InMux I__5854 (
            .O(N__27393),
            .I(N__27379));
    CascadeMux I__5853 (
            .O(N__27392),
            .I(N__27375));
    InMux I__5852 (
            .O(N__27391),
            .I(N__27371));
    InMux I__5851 (
            .O(N__27390),
            .I(N__27367));
    InMux I__5850 (
            .O(N__27389),
            .I(N__27364));
    InMux I__5849 (
            .O(N__27388),
            .I(N__27359));
    CascadeMux I__5848 (
            .O(N__27387),
            .I(N__27354));
    InMux I__5847 (
            .O(N__27386),
            .I(N__27350));
    InMux I__5846 (
            .O(N__27383),
            .I(N__27347));
    InMux I__5845 (
            .O(N__27382),
            .I(N__27343));
    LocalMux I__5844 (
            .O(N__27379),
            .I(N__27340));
    InMux I__5843 (
            .O(N__27378),
            .I(N__27337));
    InMux I__5842 (
            .O(N__27375),
            .I(N__27334));
    InMux I__5841 (
            .O(N__27374),
            .I(N__27331));
    LocalMux I__5840 (
            .O(N__27371),
            .I(N__27328));
    InMux I__5839 (
            .O(N__27370),
            .I(N__27325));
    LocalMux I__5838 (
            .O(N__27367),
            .I(N__27320));
    LocalMux I__5837 (
            .O(N__27364),
            .I(N__27320));
    InMux I__5836 (
            .O(N__27363),
            .I(N__27317));
    InMux I__5835 (
            .O(N__27362),
            .I(N__27314));
    LocalMux I__5834 (
            .O(N__27359),
            .I(N__27311));
    InMux I__5833 (
            .O(N__27358),
            .I(N__27308));
    InMux I__5832 (
            .O(N__27357),
            .I(N__27301));
    InMux I__5831 (
            .O(N__27354),
            .I(N__27301));
    InMux I__5830 (
            .O(N__27353),
            .I(N__27301));
    LocalMux I__5829 (
            .O(N__27350),
            .I(N__27298));
    LocalMux I__5828 (
            .O(N__27347),
            .I(N__27295));
    InMux I__5827 (
            .O(N__27346),
            .I(N__27290));
    LocalMux I__5826 (
            .O(N__27343),
            .I(N__27287));
    Span4Mux_h I__5825 (
            .O(N__27340),
            .I(N__27284));
    LocalMux I__5824 (
            .O(N__27337),
            .I(N__27277));
    LocalMux I__5823 (
            .O(N__27334),
            .I(N__27277));
    LocalMux I__5822 (
            .O(N__27331),
            .I(N__27277));
    Span4Mux_v I__5821 (
            .O(N__27328),
            .I(N__27272));
    LocalMux I__5820 (
            .O(N__27325),
            .I(N__27272));
    Span4Mux_h I__5819 (
            .O(N__27320),
            .I(N__27269));
    LocalMux I__5818 (
            .O(N__27317),
            .I(N__27266));
    LocalMux I__5817 (
            .O(N__27314),
            .I(N__27263));
    Span4Mux_h I__5816 (
            .O(N__27311),
            .I(N__27255));
    LocalMux I__5815 (
            .O(N__27308),
            .I(N__27255));
    LocalMux I__5814 (
            .O(N__27301),
            .I(N__27255));
    Span4Mux_v I__5813 (
            .O(N__27298),
            .I(N__27250));
    Span4Mux_h I__5812 (
            .O(N__27295),
            .I(N__27250));
    InMux I__5811 (
            .O(N__27294),
            .I(N__27245));
    InMux I__5810 (
            .O(N__27293),
            .I(N__27245));
    LocalMux I__5809 (
            .O(N__27290),
            .I(N__27242));
    Span4Mux_v I__5808 (
            .O(N__27287),
            .I(N__27233));
    Span4Mux_v I__5807 (
            .O(N__27284),
            .I(N__27233));
    Span4Mux_v I__5806 (
            .O(N__27277),
            .I(N__27233));
    Span4Mux_h I__5805 (
            .O(N__27272),
            .I(N__27233));
    Span4Mux_v I__5804 (
            .O(N__27269),
            .I(N__27226));
    Span4Mux_h I__5803 (
            .O(N__27266),
            .I(N__27226));
    Span4Mux_v I__5802 (
            .O(N__27263),
            .I(N__27226));
    InMux I__5801 (
            .O(N__27262),
            .I(N__27223));
    Span4Mux_h I__5800 (
            .O(N__27255),
            .I(N__27218));
    Span4Mux_h I__5799 (
            .O(N__27250),
            .I(N__27218));
    LocalMux I__5798 (
            .O(N__27245),
            .I(\tok.A_low_4 ));
    Odrv4 I__5797 (
            .O(N__27242),
            .I(\tok.A_low_4 ));
    Odrv4 I__5796 (
            .O(N__27233),
            .I(\tok.A_low_4 ));
    Odrv4 I__5795 (
            .O(N__27226),
            .I(\tok.A_low_4 ));
    LocalMux I__5794 (
            .O(N__27223),
            .I(\tok.A_low_4 ));
    Odrv4 I__5793 (
            .O(N__27218),
            .I(\tok.A_low_4 ));
    InMux I__5792 (
            .O(N__27205),
            .I(N__27202));
    LocalMux I__5791 (
            .O(N__27202),
            .I(N__27199));
    Span4Mux_v I__5790 (
            .O(N__27199),
            .I(N__27196));
    Span4Mux_h I__5789 (
            .O(N__27196),
            .I(N__27193));
    Odrv4 I__5788 (
            .O(N__27193),
            .I(\tok.uart.sender_6 ));
    InMux I__5787 (
            .O(N__27190),
            .I(N__27187));
    LocalMux I__5786 (
            .O(N__27187),
            .I(\tok.uart.sender_7 ));
    InMux I__5785 (
            .O(N__27184),
            .I(N__27181));
    LocalMux I__5784 (
            .O(N__27181),
            .I(\tok.uart.sender_8 ));
    CEMux I__5783 (
            .O(N__27178),
            .I(N__27175));
    LocalMux I__5782 (
            .O(N__27175),
            .I(N__27172));
    Span4Mux_s3_h I__5781 (
            .O(N__27172),
            .I(N__27167));
    CEMux I__5780 (
            .O(N__27171),
            .I(N__27164));
    CEMux I__5779 (
            .O(N__27170),
            .I(N__27160));
    Span4Mux_h I__5778 (
            .O(N__27167),
            .I(N__27155));
    LocalMux I__5777 (
            .O(N__27164),
            .I(N__27155));
    CEMux I__5776 (
            .O(N__27163),
            .I(N__27152));
    LocalMux I__5775 (
            .O(N__27160),
            .I(N__27149));
    Span4Mux_h I__5774 (
            .O(N__27155),
            .I(N__27144));
    LocalMux I__5773 (
            .O(N__27152),
            .I(N__27144));
    Span4Mux_h I__5772 (
            .O(N__27149),
            .I(N__27141));
    Span4Mux_s1_v I__5771 (
            .O(N__27144),
            .I(N__27138));
    Odrv4 I__5770 (
            .O(N__27141),
            .I(\tok.uart.n950 ));
    Odrv4 I__5769 (
            .O(N__27138),
            .I(\tok.uart.n950 ));
    InMux I__5768 (
            .O(N__27133),
            .I(N__27130));
    LocalMux I__5767 (
            .O(N__27130),
            .I(N__27126));
    InMux I__5766 (
            .O(N__27129),
            .I(N__27123));
    Span4Mux_v I__5765 (
            .O(N__27126),
            .I(N__27119));
    LocalMux I__5764 (
            .O(N__27123),
            .I(N__27116));
    InMux I__5763 (
            .O(N__27122),
            .I(N__27113));
    Span4Mux_v I__5762 (
            .O(N__27119),
            .I(N__27110));
    Span4Mux_h I__5761 (
            .O(N__27116),
            .I(N__27107));
    LocalMux I__5760 (
            .O(N__27113),
            .I(N__27104));
    Span4Mux_h I__5759 (
            .O(N__27110),
            .I(N__27099));
    Span4Mux_v I__5758 (
            .O(N__27107),
            .I(N__27099));
    Span4Mux_v I__5757 (
            .O(N__27104),
            .I(N__27096));
    Odrv4 I__5756 (
            .O(N__27099),
            .I(\tok.n274 ));
    Odrv4 I__5755 (
            .O(N__27096),
            .I(\tok.n274 ));
    InMux I__5754 (
            .O(N__27091),
            .I(N__27087));
    InMux I__5753 (
            .O(N__27090),
            .I(N__27084));
    LocalMux I__5752 (
            .O(N__27087),
            .I(N__27080));
    LocalMux I__5751 (
            .O(N__27084),
            .I(N__27077));
    InMux I__5750 (
            .O(N__27083),
            .I(N__27074));
    Span4Mux_s2_h I__5749 (
            .O(N__27080),
            .I(N__27069));
    Span4Mux_h I__5748 (
            .O(N__27077),
            .I(N__27069));
    LocalMux I__5747 (
            .O(N__27074),
            .I(N__27066));
    Span4Mux_v I__5746 (
            .O(N__27069),
            .I(N__27063));
    Odrv4 I__5745 (
            .O(N__27066),
            .I(\tok.n185 ));
    Odrv4 I__5744 (
            .O(N__27063),
            .I(\tok.n185 ));
    InMux I__5743 (
            .O(N__27058),
            .I(N__27055));
    LocalMux I__5742 (
            .O(N__27055),
            .I(N__27052));
    Span4Mux_h I__5741 (
            .O(N__27052),
            .I(N__27049));
    Odrv4 I__5740 (
            .O(N__27049),
            .I(\tok.n7410 ));
    CascadeMux I__5739 (
            .O(N__27046),
            .I(\tok.n2598_cascade_ ));
    InMux I__5738 (
            .O(N__27043),
            .I(N__27040));
    LocalMux I__5737 (
            .O(N__27040),
            .I(N__27033));
    InMux I__5736 (
            .O(N__27039),
            .I(N__27030));
    InMux I__5735 (
            .O(N__27038),
            .I(N__27027));
    InMux I__5734 (
            .O(N__27037),
            .I(N__27024));
    InMux I__5733 (
            .O(N__27036),
            .I(N__27019));
    Span4Mux_v I__5732 (
            .O(N__27033),
            .I(N__27013));
    LocalMux I__5731 (
            .O(N__27030),
            .I(N__27013));
    LocalMux I__5730 (
            .O(N__27027),
            .I(N__27008));
    LocalMux I__5729 (
            .O(N__27024),
            .I(N__27005));
    InMux I__5728 (
            .O(N__27023),
            .I(N__27000));
    InMux I__5727 (
            .O(N__27022),
            .I(N__27000));
    LocalMux I__5726 (
            .O(N__27019),
            .I(N__26997));
    InMux I__5725 (
            .O(N__27018),
            .I(N__26994));
    Span4Mux_s3_h I__5724 (
            .O(N__27013),
            .I(N__26991));
    CascadeMux I__5723 (
            .O(N__27012),
            .I(N__26988));
    InMux I__5722 (
            .O(N__27011),
            .I(N__26984));
    Span12Mux_s8_v I__5721 (
            .O(N__27008),
            .I(N__26981));
    Span4Mux_h I__5720 (
            .O(N__27005),
            .I(N__26976));
    LocalMux I__5719 (
            .O(N__27000),
            .I(N__26976));
    Span4Mux_h I__5718 (
            .O(N__26997),
            .I(N__26973));
    LocalMux I__5717 (
            .O(N__26994),
            .I(N__26970));
    Span4Mux_h I__5716 (
            .O(N__26991),
            .I(N__26967));
    InMux I__5715 (
            .O(N__26988),
            .I(N__26962));
    InMux I__5714 (
            .O(N__26987),
            .I(N__26962));
    LocalMux I__5713 (
            .O(N__26984),
            .I(\tok.n45 ));
    Odrv12 I__5712 (
            .O(N__26981),
            .I(\tok.n45 ));
    Odrv4 I__5711 (
            .O(N__26976),
            .I(\tok.n45 ));
    Odrv4 I__5710 (
            .O(N__26973),
            .I(\tok.n45 ));
    Odrv12 I__5709 (
            .O(N__26970),
            .I(\tok.n45 ));
    Odrv4 I__5708 (
            .O(N__26967),
            .I(\tok.n45 ));
    LocalMux I__5707 (
            .O(N__26962),
            .I(\tok.n45 ));
    InMux I__5706 (
            .O(N__26947),
            .I(N__26944));
    LocalMux I__5705 (
            .O(N__26944),
            .I(N__26941));
    Odrv4 I__5704 (
            .O(N__26941),
            .I(\tok.n6390 ));
    InMux I__5703 (
            .O(N__26938),
            .I(N__26934));
    CascadeMux I__5702 (
            .O(N__26937),
            .I(N__26928));
    LocalMux I__5701 (
            .O(N__26934),
            .I(N__26923));
    InMux I__5700 (
            .O(N__26933),
            .I(N__26920));
    InMux I__5699 (
            .O(N__26932),
            .I(N__26917));
    InMux I__5698 (
            .O(N__26931),
            .I(N__26912));
    InMux I__5697 (
            .O(N__26928),
            .I(N__26912));
    InMux I__5696 (
            .O(N__26927),
            .I(N__26907));
    InMux I__5695 (
            .O(N__26926),
            .I(N__26907));
    Span4Mux_h I__5694 (
            .O(N__26923),
            .I(N__26899));
    LocalMux I__5693 (
            .O(N__26920),
            .I(N__26899));
    LocalMux I__5692 (
            .O(N__26917),
            .I(N__26899));
    LocalMux I__5691 (
            .O(N__26912),
            .I(N__26894));
    LocalMux I__5690 (
            .O(N__26907),
            .I(N__26894));
    InMux I__5689 (
            .O(N__26906),
            .I(N__26891));
    Span4Mux_h I__5688 (
            .O(N__26899),
            .I(N__26888));
    Span4Mux_h I__5687 (
            .O(N__26894),
            .I(N__26883));
    LocalMux I__5686 (
            .O(N__26891),
            .I(N__26883));
    Odrv4 I__5685 (
            .O(N__26888),
            .I(\tok.n821 ));
    Odrv4 I__5684 (
            .O(N__26883),
            .I(\tok.n821 ));
    CascadeMux I__5683 (
            .O(N__26878),
            .I(\tok.n215_cascade_ ));
    InMux I__5682 (
            .O(N__26875),
            .I(N__26872));
    LocalMux I__5681 (
            .O(N__26872),
            .I(N__26869));
    Span4Mux_v I__5680 (
            .O(N__26869),
            .I(N__26866));
    Odrv4 I__5679 (
            .O(N__26866),
            .I(\tok.n6547 ));
    InMux I__5678 (
            .O(N__26863),
            .I(N__26860));
    LocalMux I__5677 (
            .O(N__26860),
            .I(N__26857));
    Span4Mux_s2_h I__5676 (
            .O(N__26857),
            .I(N__26853));
    InMux I__5675 (
            .O(N__26856),
            .I(N__26850));
    Span4Mux_v I__5674 (
            .O(N__26853),
            .I(N__26845));
    LocalMux I__5673 (
            .O(N__26850),
            .I(N__26845));
    Odrv4 I__5672 (
            .O(N__26845),
            .I(\tok.n4_adj_712 ));
    InMux I__5671 (
            .O(N__26842),
            .I(N__26839));
    LocalMux I__5670 (
            .O(N__26839),
            .I(N__26835));
    InMux I__5669 (
            .O(N__26838),
            .I(N__26832));
    Span4Mux_s3_h I__5668 (
            .O(N__26835),
            .I(N__26828));
    LocalMux I__5667 (
            .O(N__26832),
            .I(N__26825));
    InMux I__5666 (
            .O(N__26831),
            .I(N__26822));
    Span4Mux_v I__5665 (
            .O(N__26828),
            .I(N__26815));
    Span4Mux_s3_h I__5664 (
            .O(N__26825),
            .I(N__26815));
    LocalMux I__5663 (
            .O(N__26822),
            .I(N__26815));
    Span4Mux_h I__5662 (
            .O(N__26815),
            .I(N__26812));
    Span4Mux_h I__5661 (
            .O(N__26812),
            .I(N__26809));
    Odrv4 I__5660 (
            .O(N__26809),
            .I(\tok.n238 ));
    CascadeMux I__5659 (
            .O(N__26806),
            .I(\tok.n6650_cascade_ ));
    InMux I__5658 (
            .O(N__26803),
            .I(N__26799));
    CascadeMux I__5657 (
            .O(N__26802),
            .I(N__26794));
    LocalMux I__5656 (
            .O(N__26799),
            .I(N__26789));
    InMux I__5655 (
            .O(N__26798),
            .I(N__26786));
    InMux I__5654 (
            .O(N__26797),
            .I(N__26781));
    InMux I__5653 (
            .O(N__26794),
            .I(N__26781));
    InMux I__5652 (
            .O(N__26793),
            .I(N__26776));
    InMux I__5651 (
            .O(N__26792),
            .I(N__26769));
    Span4Mux_v I__5650 (
            .O(N__26789),
            .I(N__26762));
    LocalMux I__5649 (
            .O(N__26786),
            .I(N__26762));
    LocalMux I__5648 (
            .O(N__26781),
            .I(N__26759));
    InMux I__5647 (
            .O(N__26780),
            .I(N__26755));
    InMux I__5646 (
            .O(N__26779),
            .I(N__26752));
    LocalMux I__5645 (
            .O(N__26776),
            .I(N__26749));
    InMux I__5644 (
            .O(N__26775),
            .I(N__26746));
    InMux I__5643 (
            .O(N__26774),
            .I(N__26739));
    InMux I__5642 (
            .O(N__26773),
            .I(N__26739));
    InMux I__5641 (
            .O(N__26772),
            .I(N__26739));
    LocalMux I__5640 (
            .O(N__26769),
            .I(N__26733));
    InMux I__5639 (
            .O(N__26768),
            .I(N__26728));
    InMux I__5638 (
            .O(N__26767),
            .I(N__26728));
    Span4Mux_h I__5637 (
            .O(N__26762),
            .I(N__26723));
    Span4Mux_h I__5636 (
            .O(N__26759),
            .I(N__26723));
    InMux I__5635 (
            .O(N__26758),
            .I(N__26720));
    LocalMux I__5634 (
            .O(N__26755),
            .I(N__26717));
    LocalMux I__5633 (
            .O(N__26752),
            .I(N__26714));
    Span4Mux_v I__5632 (
            .O(N__26749),
            .I(N__26709));
    LocalMux I__5631 (
            .O(N__26746),
            .I(N__26709));
    LocalMux I__5630 (
            .O(N__26739),
            .I(N__26706));
    InMux I__5629 (
            .O(N__26738),
            .I(N__26703));
    InMux I__5628 (
            .O(N__26737),
            .I(N__26698));
    InMux I__5627 (
            .O(N__26736),
            .I(N__26698));
    Span4Mux_s1_v I__5626 (
            .O(N__26733),
            .I(N__26689));
    LocalMux I__5625 (
            .O(N__26728),
            .I(N__26689));
    Span4Mux_h I__5624 (
            .O(N__26723),
            .I(N__26689));
    LocalMux I__5623 (
            .O(N__26720),
            .I(N__26689));
    Span4Mux_v I__5622 (
            .O(N__26717),
            .I(N__26680));
    Span4Mux_v I__5621 (
            .O(N__26714),
            .I(N__26680));
    Span4Mux_h I__5620 (
            .O(N__26709),
            .I(N__26680));
    Span4Mux_v I__5619 (
            .O(N__26706),
            .I(N__26680));
    LocalMux I__5618 (
            .O(N__26703),
            .I(\tok.n48 ));
    LocalMux I__5617 (
            .O(N__26698),
            .I(\tok.n48 ));
    Odrv4 I__5616 (
            .O(N__26689),
            .I(\tok.n48 ));
    Odrv4 I__5615 (
            .O(N__26680),
            .I(\tok.n48 ));
    CascadeMux I__5614 (
            .O(N__26671),
            .I(\tok.n211_cascade_ ));
    CascadeMux I__5613 (
            .O(N__26668),
            .I(N__26665));
    InMux I__5612 (
            .O(N__26665),
            .I(N__26662));
    LocalMux I__5611 (
            .O(N__26662),
            .I(N__26659));
    Span4Mux_s3_v I__5610 (
            .O(N__26659),
            .I(N__26656));
    Span4Mux_h I__5609 (
            .O(N__26656),
            .I(N__26653));
    Span4Mux_h I__5608 (
            .O(N__26653),
            .I(N__26650));
    Span4Mux_v I__5607 (
            .O(N__26650),
            .I(N__26647));
    Odrv4 I__5606 (
            .O(N__26647),
            .I(\tok.n6644 ));
    CascadeMux I__5605 (
            .O(N__26644),
            .I(\tok.n260_cascade_ ));
    CascadeMux I__5604 (
            .O(N__26641),
            .I(N__26638));
    InMux I__5603 (
            .O(N__26638),
            .I(N__26635));
    LocalMux I__5602 (
            .O(N__26635),
            .I(N__26632));
    Odrv4 I__5601 (
            .O(N__26632),
            .I(\tok.n6501 ));
    CascadeMux I__5600 (
            .O(N__26629),
            .I(\tok.n186_adj_798_cascade_ ));
    InMux I__5599 (
            .O(N__26626),
            .I(N__26623));
    LocalMux I__5598 (
            .O(N__26623),
            .I(N__26620));
    Odrv4 I__5597 (
            .O(N__26620),
            .I(\tok.n6496 ));
    CascadeMux I__5596 (
            .O(N__26617),
            .I(N__26612));
    CascadeMux I__5595 (
            .O(N__26616),
            .I(N__26605));
    CascadeMux I__5594 (
            .O(N__26615),
            .I(N__26602));
    InMux I__5593 (
            .O(N__26612),
            .I(N__26597));
    InMux I__5592 (
            .O(N__26611),
            .I(N__26597));
    InMux I__5591 (
            .O(N__26610),
            .I(N__26594));
    InMux I__5590 (
            .O(N__26609),
            .I(N__26591));
    InMux I__5589 (
            .O(N__26608),
            .I(N__26588));
    InMux I__5588 (
            .O(N__26605),
            .I(N__26578));
    InMux I__5587 (
            .O(N__26602),
            .I(N__26578));
    LocalMux I__5586 (
            .O(N__26597),
            .I(N__26575));
    LocalMux I__5585 (
            .O(N__26594),
            .I(N__26570));
    LocalMux I__5584 (
            .O(N__26591),
            .I(N__26570));
    LocalMux I__5583 (
            .O(N__26588),
            .I(N__26567));
    InMux I__5582 (
            .O(N__26587),
            .I(N__26564));
    InMux I__5581 (
            .O(N__26586),
            .I(N__26561));
    InMux I__5580 (
            .O(N__26585),
            .I(N__26556));
    InMux I__5579 (
            .O(N__26584),
            .I(N__26556));
    InMux I__5578 (
            .O(N__26583),
            .I(N__26553));
    LocalMux I__5577 (
            .O(N__26578),
            .I(N__26548));
    Span4Mux_h I__5576 (
            .O(N__26575),
            .I(N__26548));
    Span4Mux_h I__5575 (
            .O(N__26570),
            .I(N__26543));
    Span4Mux_h I__5574 (
            .O(N__26567),
            .I(N__26543));
    LocalMux I__5573 (
            .O(N__26564),
            .I(\tok.n194 ));
    LocalMux I__5572 (
            .O(N__26561),
            .I(\tok.n194 ));
    LocalMux I__5571 (
            .O(N__26556),
            .I(\tok.n194 ));
    LocalMux I__5570 (
            .O(N__26553),
            .I(\tok.n194 ));
    Odrv4 I__5569 (
            .O(N__26548),
            .I(\tok.n194 ));
    Odrv4 I__5568 (
            .O(N__26543),
            .I(\tok.n194 ));
    CascadeMux I__5567 (
            .O(N__26530),
            .I(\tok.n338_adj_805_cascade_ ));
    InMux I__5566 (
            .O(N__26527),
            .I(N__26524));
    LocalMux I__5565 (
            .O(N__26524),
            .I(N__26521));
    Span4Mux_h I__5564 (
            .O(N__26521),
            .I(N__26518));
    Span4Mux_v I__5563 (
            .O(N__26518),
            .I(N__26515));
    Odrv4 I__5562 (
            .O(N__26515),
            .I(\tok.n6608 ));
    InMux I__5561 (
            .O(N__26512),
            .I(N__26508));
    CascadeMux I__5560 (
            .O(N__26511),
            .I(N__26505));
    LocalMux I__5559 (
            .O(N__26508),
            .I(N__26501));
    InMux I__5558 (
            .O(N__26505),
            .I(N__26497));
    InMux I__5557 (
            .O(N__26504),
            .I(N__26493));
    Span4Mux_h I__5556 (
            .O(N__26501),
            .I(N__26490));
    InMux I__5555 (
            .O(N__26500),
            .I(N__26487));
    LocalMux I__5554 (
            .O(N__26497),
            .I(N__26484));
    InMux I__5553 (
            .O(N__26496),
            .I(N__26480));
    LocalMux I__5552 (
            .O(N__26493),
            .I(N__26477));
    Span4Mux_v I__5551 (
            .O(N__26490),
            .I(N__26474));
    LocalMux I__5550 (
            .O(N__26487),
            .I(N__26469));
    Span4Mux_h I__5549 (
            .O(N__26484),
            .I(N__26469));
    InMux I__5548 (
            .O(N__26483),
            .I(N__26466));
    LocalMux I__5547 (
            .O(N__26480),
            .I(N__26463));
    Span4Mux_h I__5546 (
            .O(N__26477),
            .I(N__26458));
    Span4Mux_h I__5545 (
            .O(N__26474),
            .I(N__26458));
    Span4Mux_v I__5544 (
            .O(N__26469),
            .I(N__26453));
    LocalMux I__5543 (
            .O(N__26466),
            .I(N__26453));
    Odrv4 I__5542 (
            .O(N__26463),
            .I(\tok.n219 ));
    Odrv4 I__5541 (
            .O(N__26458),
            .I(\tok.n219 ));
    Odrv4 I__5540 (
            .O(N__26453),
            .I(\tok.n219 ));
    InMux I__5539 (
            .O(N__26446),
            .I(N__26440));
    InMux I__5538 (
            .O(N__26445),
            .I(N__26440));
    LocalMux I__5537 (
            .O(N__26440),
            .I(N__26437));
    Odrv4 I__5536 (
            .O(N__26437),
            .I(\tok.n190_adj_792 ));
    InMux I__5535 (
            .O(N__26434),
            .I(N__26431));
    LocalMux I__5534 (
            .O(N__26431),
            .I(N__26428));
    Odrv12 I__5533 (
            .O(N__26428),
            .I(\tok.n4_adj_804 ));
    InMux I__5532 (
            .O(N__26425),
            .I(N__26422));
    LocalMux I__5531 (
            .O(N__26422),
            .I(N__26419));
    Odrv4 I__5530 (
            .O(N__26419),
            .I(\tok.n174_adj_803 ));
    InMux I__5529 (
            .O(N__26416),
            .I(N__26413));
    LocalMux I__5528 (
            .O(N__26413),
            .I(\tok.n205_adj_806 ));
    InMux I__5527 (
            .O(N__26410),
            .I(N__26407));
    LocalMux I__5526 (
            .O(N__26407),
            .I(N__26404));
    Span4Mux_v I__5525 (
            .O(N__26404),
            .I(N__26401));
    Span4Mux_h I__5524 (
            .O(N__26401),
            .I(N__26398));
    Odrv4 I__5523 (
            .O(N__26398),
            .I(\tok.n177_adj_813 ));
    CascadeMux I__5522 (
            .O(N__26395),
            .I(\tok.n252_adj_801_cascade_ ));
    CascadeMux I__5521 (
            .O(N__26392),
            .I(N__26388));
    CascadeMux I__5520 (
            .O(N__26391),
            .I(N__26385));
    InMux I__5519 (
            .O(N__26388),
            .I(N__26380));
    InMux I__5518 (
            .O(N__26385),
            .I(N__26377));
    InMux I__5517 (
            .O(N__26384),
            .I(N__26374));
    InMux I__5516 (
            .O(N__26383),
            .I(N__26371));
    LocalMux I__5515 (
            .O(N__26380),
            .I(N__26368));
    LocalMux I__5514 (
            .O(N__26377),
            .I(N__26365));
    LocalMux I__5513 (
            .O(N__26374),
            .I(N__26360));
    LocalMux I__5512 (
            .O(N__26371),
            .I(N__26360));
    Span4Mux_h I__5511 (
            .O(N__26368),
            .I(N__26355));
    Span4Mux_s3_h I__5510 (
            .O(N__26365),
            .I(N__26355));
    Odrv12 I__5509 (
            .O(N__26360),
            .I(\tok.n867 ));
    Odrv4 I__5508 (
            .O(N__26355),
            .I(\tok.n867 ));
    InMux I__5507 (
            .O(N__26350),
            .I(N__26346));
    InMux I__5506 (
            .O(N__26349),
            .I(N__26343));
    LocalMux I__5505 (
            .O(N__26346),
            .I(N__26340));
    LocalMux I__5504 (
            .O(N__26343),
            .I(N__26337));
    Span4Mux_s2_h I__5503 (
            .O(N__26340),
            .I(N__26334));
    Span4Mux_h I__5502 (
            .O(N__26337),
            .I(N__26331));
    Span4Mux_h I__5501 (
            .O(N__26334),
            .I(N__26328));
    Span4Mux_h I__5500 (
            .O(N__26331),
            .I(N__26325));
    Span4Mux_h I__5499 (
            .O(N__26328),
            .I(N__26322));
    Odrv4 I__5498 (
            .O(N__26325),
            .I(\tok.n233 ));
    Odrv4 I__5497 (
            .O(N__26322),
            .I(\tok.n233 ));
    InMux I__5496 (
            .O(N__26317),
            .I(N__26312));
    InMux I__5495 (
            .O(N__26316),
            .I(N__26309));
    InMux I__5494 (
            .O(N__26315),
            .I(N__26306));
    LocalMux I__5493 (
            .O(N__26312),
            .I(N__26302));
    LocalMux I__5492 (
            .O(N__26309),
            .I(N__26299));
    LocalMux I__5491 (
            .O(N__26306),
            .I(N__26296));
    InMux I__5490 (
            .O(N__26305),
            .I(N__26293));
    Span4Mux_v I__5489 (
            .O(N__26302),
            .I(N__26288));
    Span4Mux_v I__5488 (
            .O(N__26299),
            .I(N__26288));
    Span4Mux_v I__5487 (
            .O(N__26296),
            .I(N__26282));
    LocalMux I__5486 (
            .O(N__26293),
            .I(N__26282));
    Span4Mux_h I__5485 (
            .O(N__26288),
            .I(N__26279));
    InMux I__5484 (
            .O(N__26287),
            .I(N__26276));
    Odrv4 I__5483 (
            .O(N__26282),
            .I(\tok.n5_adj_745 ));
    Odrv4 I__5482 (
            .O(N__26279),
            .I(\tok.n5_adj_745 ));
    LocalMux I__5481 (
            .O(N__26276),
            .I(\tok.n5_adj_745 ));
    CascadeMux I__5480 (
            .O(N__26269),
            .I(\tok.n255_adj_793_cascade_ ));
    InMux I__5479 (
            .O(N__26266),
            .I(N__26263));
    LocalMux I__5478 (
            .O(N__26263),
            .I(\tok.n258_adj_800 ));
    InMux I__5477 (
            .O(N__26260),
            .I(N__26256));
    InMux I__5476 (
            .O(N__26259),
            .I(N__26253));
    LocalMux I__5475 (
            .O(N__26256),
            .I(N__26250));
    LocalMux I__5474 (
            .O(N__26253),
            .I(N__26247));
    Sp12to4 I__5473 (
            .O(N__26250),
            .I(N__26244));
    Span12Mux_s11_v I__5472 (
            .O(N__26247),
            .I(N__26241));
    Odrv12 I__5471 (
            .O(N__26244),
            .I(\tok.n6183 ));
    Odrv12 I__5470 (
            .O(N__26241),
            .I(\tok.n6183 ));
    CascadeMux I__5469 (
            .O(N__26236),
            .I(\tok.n6162_cascade_ ));
    CascadeMux I__5468 (
            .O(N__26233),
            .I(\tok.n865_cascade_ ));
    CascadeMux I__5467 (
            .O(N__26230),
            .I(\tok.n222_cascade_ ));
    CascadeMux I__5466 (
            .O(N__26227),
            .I(N__26223));
    CascadeMux I__5465 (
            .O(N__26226),
            .I(N__26218));
    InMux I__5464 (
            .O(N__26223),
            .I(N__26214));
    CascadeMux I__5463 (
            .O(N__26222),
            .I(N__26211));
    CascadeMux I__5462 (
            .O(N__26221),
            .I(N__26208));
    InMux I__5461 (
            .O(N__26218),
            .I(N__26204));
    CascadeMux I__5460 (
            .O(N__26217),
            .I(N__26201));
    LocalMux I__5459 (
            .O(N__26214),
            .I(N__26198));
    InMux I__5458 (
            .O(N__26211),
            .I(N__26195));
    InMux I__5457 (
            .O(N__26208),
            .I(N__26192));
    InMux I__5456 (
            .O(N__26207),
            .I(N__26189));
    LocalMux I__5455 (
            .O(N__26204),
            .I(N__26186));
    InMux I__5454 (
            .O(N__26201),
            .I(N__26183));
    Span4Mux_h I__5453 (
            .O(N__26198),
            .I(N__26176));
    LocalMux I__5452 (
            .O(N__26195),
            .I(N__26176));
    LocalMux I__5451 (
            .O(N__26192),
            .I(N__26173));
    LocalMux I__5450 (
            .O(N__26189),
            .I(N__26166));
    Span4Mux_h I__5449 (
            .O(N__26186),
            .I(N__26166));
    LocalMux I__5448 (
            .O(N__26183),
            .I(N__26166));
    InMux I__5447 (
            .O(N__26182),
            .I(N__26163));
    InMux I__5446 (
            .O(N__26181),
            .I(N__26160));
    Span4Mux_v I__5445 (
            .O(N__26176),
            .I(N__26157));
    Span4Mux_v I__5444 (
            .O(N__26173),
            .I(N__26152));
    Span4Mux_v I__5443 (
            .O(N__26166),
            .I(N__26152));
    LocalMux I__5442 (
            .O(N__26163),
            .I(N__26147));
    LocalMux I__5441 (
            .O(N__26160),
            .I(N__26147));
    Span4Mux_h I__5440 (
            .O(N__26157),
            .I(N__26144));
    Span4Mux_h I__5439 (
            .O(N__26152),
            .I(N__26141));
    Span12Mux_s4_h I__5438 (
            .O(N__26147),
            .I(N__26138));
    Odrv4 I__5437 (
            .O(N__26144),
            .I(\tok.n245 ));
    Odrv4 I__5436 (
            .O(N__26141),
            .I(\tok.n245 ));
    Odrv12 I__5435 (
            .O(N__26138),
            .I(\tok.n245 ));
    CascadeMux I__5434 (
            .O(N__26131),
            .I(N__26126));
    InMux I__5433 (
            .O(N__26130),
            .I(N__26123));
    InMux I__5432 (
            .O(N__26129),
            .I(N__26120));
    InMux I__5431 (
            .O(N__26126),
            .I(N__26117));
    LocalMux I__5430 (
            .O(N__26123),
            .I(N__26114));
    LocalMux I__5429 (
            .O(N__26120),
            .I(N__26111));
    LocalMux I__5428 (
            .O(N__26117),
            .I(N__26106));
    Span4Mux_h I__5427 (
            .O(N__26114),
            .I(N__26106));
    Span4Mux_h I__5426 (
            .O(N__26111),
            .I(N__26103));
    Odrv4 I__5425 (
            .O(N__26106),
            .I(\tok.n4_adj_648 ));
    Odrv4 I__5424 (
            .O(N__26103),
            .I(\tok.n4_adj_648 ));
    InMux I__5423 (
            .O(N__26098),
            .I(N__26095));
    LocalMux I__5422 (
            .O(N__26095),
            .I(N__26092));
    Span4Mux_v I__5421 (
            .O(N__26092),
            .I(N__26089));
    Span4Mux_h I__5420 (
            .O(N__26089),
            .I(N__26086));
    Span4Mux_h I__5419 (
            .O(N__26086),
            .I(N__26083));
    Odrv4 I__5418 (
            .O(N__26083),
            .I(\tok.n2635 ));
    CascadeMux I__5417 (
            .O(N__26080),
            .I(\tok.n6653_cascade_ ));
    CascadeMux I__5416 (
            .O(N__26077),
            .I(\tok.n6646_cascade_ ));
    CascadeMux I__5415 (
            .O(N__26074),
            .I(N__26071));
    InMux I__5414 (
            .O(N__26071),
            .I(N__26068));
    LocalMux I__5413 (
            .O(N__26068),
            .I(\tok.n6167 ));
    InMux I__5412 (
            .O(N__26065),
            .I(N__26062));
    LocalMux I__5411 (
            .O(N__26062),
            .I(N__26059));
    Span4Mux_v I__5410 (
            .O(N__26059),
            .I(N__26056));
    Odrv4 I__5409 (
            .O(N__26056),
            .I(\tok.n6645 ));
    CascadeMux I__5408 (
            .O(N__26053),
            .I(N__26050));
    InMux I__5407 (
            .O(N__26050),
            .I(N__26047));
    LocalMux I__5406 (
            .O(N__26047),
            .I(N__26044));
    Span4Mux_h I__5405 (
            .O(N__26044),
            .I(N__26041));
    Odrv4 I__5404 (
            .O(N__26041),
            .I(\tok.n247 ));
    InMux I__5403 (
            .O(N__26038),
            .I(N__26035));
    LocalMux I__5402 (
            .O(N__26035),
            .I(\tok.n6639 ));
    InMux I__5401 (
            .O(N__26032),
            .I(N__26029));
    LocalMux I__5400 (
            .O(N__26029),
            .I(\tok.n280 ));
    CascadeMux I__5399 (
            .O(N__26026),
            .I(\tok.n6638_cascade_ ));
    InMux I__5398 (
            .O(N__26023),
            .I(N__26020));
    LocalMux I__5397 (
            .O(N__26020),
            .I(N__26017));
    Odrv4 I__5396 (
            .O(N__26017),
            .I(\tok.n6636 ));
    InMux I__5395 (
            .O(N__26014),
            .I(N__26010));
    InMux I__5394 (
            .O(N__26013),
            .I(N__26007));
    LocalMux I__5393 (
            .O(N__26010),
            .I(N__26004));
    LocalMux I__5392 (
            .O(N__26007),
            .I(N__25999));
    Span4Mux_v I__5391 (
            .O(N__26004),
            .I(N__25999));
    Span4Mux_h I__5390 (
            .O(N__25999),
            .I(N__25996));
    Odrv4 I__5389 (
            .O(N__25996),
            .I(\tok.n260_adj_717 ));
    InMux I__5388 (
            .O(N__25993),
            .I(N__25989));
    CascadeMux I__5387 (
            .O(N__25992),
            .I(N__25985));
    LocalMux I__5386 (
            .O(N__25989),
            .I(N__25981));
    CascadeMux I__5385 (
            .O(N__25988),
            .I(N__25978));
    InMux I__5384 (
            .O(N__25985),
            .I(N__25975));
    CascadeMux I__5383 (
            .O(N__25984),
            .I(N__25972));
    Span4Mux_v I__5382 (
            .O(N__25981),
            .I(N__25968));
    InMux I__5381 (
            .O(N__25978),
            .I(N__25965));
    LocalMux I__5380 (
            .O(N__25975),
            .I(N__25961));
    InMux I__5379 (
            .O(N__25972),
            .I(N__25958));
    CascadeMux I__5378 (
            .O(N__25971),
            .I(N__25955));
    Span4Mux_h I__5377 (
            .O(N__25968),
            .I(N__25950));
    LocalMux I__5376 (
            .O(N__25965),
            .I(N__25950));
    InMux I__5375 (
            .O(N__25964),
            .I(N__25947));
    Span4Mux_v I__5374 (
            .O(N__25961),
            .I(N__25944));
    LocalMux I__5373 (
            .O(N__25958),
            .I(N__25941));
    InMux I__5372 (
            .O(N__25955),
            .I(N__25938));
    Span4Mux_v I__5371 (
            .O(N__25950),
            .I(N__25933));
    LocalMux I__5370 (
            .O(N__25947),
            .I(N__25930));
    Span4Mux_h I__5369 (
            .O(N__25944),
            .I(N__25927));
    Span4Mux_v I__5368 (
            .O(N__25941),
            .I(N__25924));
    LocalMux I__5367 (
            .O(N__25938),
            .I(N__25921));
    InMux I__5366 (
            .O(N__25937),
            .I(N__25918));
    InMux I__5365 (
            .O(N__25936),
            .I(N__25915));
    Span4Mux_h I__5364 (
            .O(N__25933),
            .I(N__25912));
    Span4Mux_h I__5363 (
            .O(N__25930),
            .I(N__25903));
    Span4Mux_h I__5362 (
            .O(N__25927),
            .I(N__25903));
    Span4Mux_v I__5361 (
            .O(N__25924),
            .I(N__25903));
    Span4Mux_v I__5360 (
            .O(N__25921),
            .I(N__25903));
    LocalMux I__5359 (
            .O(N__25918),
            .I(\tok.S_6 ));
    LocalMux I__5358 (
            .O(N__25915),
            .I(\tok.S_6 ));
    Odrv4 I__5357 (
            .O(N__25912),
            .I(\tok.S_6 ));
    Odrv4 I__5356 (
            .O(N__25903),
            .I(\tok.S_6 ));
    InMux I__5355 (
            .O(N__25894),
            .I(N__25889));
    InMux I__5354 (
            .O(N__25893),
            .I(N__25886));
    InMux I__5353 (
            .O(N__25892),
            .I(N__25883));
    LocalMux I__5352 (
            .O(N__25889),
            .I(N__25879));
    LocalMux I__5351 (
            .O(N__25886),
            .I(N__25876));
    LocalMux I__5350 (
            .O(N__25883),
            .I(N__25872));
    InMux I__5349 (
            .O(N__25882),
            .I(N__25869));
    Span4Mux_h I__5348 (
            .O(N__25879),
            .I(N__25864));
    Span4Mux_v I__5347 (
            .O(N__25876),
            .I(N__25864));
    InMux I__5346 (
            .O(N__25875),
            .I(N__25861));
    Span4Mux_v I__5345 (
            .O(N__25872),
            .I(N__25858));
    LocalMux I__5344 (
            .O(N__25869),
            .I(N__25855));
    Span4Mux_v I__5343 (
            .O(N__25864),
            .I(N__25852));
    LocalMux I__5342 (
            .O(N__25861),
            .I(N__25845));
    Span4Mux_h I__5341 (
            .O(N__25858),
            .I(N__25845));
    Span4Mux_v I__5340 (
            .O(N__25855),
            .I(N__25845));
    Odrv4 I__5339 (
            .O(N__25852),
            .I(\tok.n815 ));
    Odrv4 I__5338 (
            .O(N__25845),
            .I(\tok.n815 ));
    InMux I__5337 (
            .O(N__25840),
            .I(N__25837));
    LocalMux I__5336 (
            .O(N__25837),
            .I(N__25834));
    Odrv4 I__5335 (
            .O(N__25834),
            .I(\tok.n6510 ));
    CascadeMux I__5334 (
            .O(N__25831),
            .I(\tok.n177_adj_799_cascade_ ));
    InMux I__5333 (
            .O(N__25828),
            .I(N__25825));
    LocalMux I__5332 (
            .O(N__25825),
            .I(N__25822));
    Odrv12 I__5331 (
            .O(N__25822),
            .I(\tok.n127_adj_772 ));
    CascadeMux I__5330 (
            .O(N__25819),
            .I(\tok.n10_adj_773_cascade_ ));
    CascadeMux I__5329 (
            .O(N__25816),
            .I(\tok.n6146_cascade_ ));
    InMux I__5328 (
            .O(N__25813),
            .I(N__25810));
    LocalMux I__5327 (
            .O(N__25810),
            .I(N__25801));
    InMux I__5326 (
            .O(N__25809),
            .I(N__25798));
    InMux I__5325 (
            .O(N__25808),
            .I(N__25794));
    InMux I__5324 (
            .O(N__25807),
            .I(N__25791));
    InMux I__5323 (
            .O(N__25806),
            .I(N__25788));
    InMux I__5322 (
            .O(N__25805),
            .I(N__25785));
    InMux I__5321 (
            .O(N__25804),
            .I(N__25782));
    Span4Mux_h I__5320 (
            .O(N__25801),
            .I(N__25779));
    LocalMux I__5319 (
            .O(N__25798),
            .I(N__25776));
    InMux I__5318 (
            .O(N__25797),
            .I(N__25773));
    LocalMux I__5317 (
            .O(N__25794),
            .I(N__25768));
    LocalMux I__5316 (
            .O(N__25791),
            .I(N__25768));
    LocalMux I__5315 (
            .O(N__25788),
            .I(N__25763));
    LocalMux I__5314 (
            .O(N__25785),
            .I(N__25763));
    LocalMux I__5313 (
            .O(N__25782),
            .I(N__25756));
    Span4Mux_v I__5312 (
            .O(N__25779),
            .I(N__25756));
    Span4Mux_h I__5311 (
            .O(N__25776),
            .I(N__25756));
    LocalMux I__5310 (
            .O(N__25773),
            .I(N__25749));
    Span4Mux_s3_v I__5309 (
            .O(N__25768),
            .I(N__25749));
    Span4Mux_h I__5308 (
            .O(N__25763),
            .I(N__25749));
    Span4Mux_h I__5307 (
            .O(N__25756),
            .I(N__25746));
    Span4Mux_h I__5306 (
            .O(N__25749),
            .I(N__25743));
    Odrv4 I__5305 (
            .O(N__25746),
            .I(\tok.n86 ));
    Odrv4 I__5304 (
            .O(N__25743),
            .I(\tok.n86 ));
    InMux I__5303 (
            .O(N__25738),
            .I(N__25734));
    InMux I__5302 (
            .O(N__25737),
            .I(N__25731));
    LocalMux I__5301 (
            .O(N__25734),
            .I(N__25728));
    LocalMux I__5300 (
            .O(N__25731),
            .I(N__25724));
    Span4Mux_s2_h I__5299 (
            .O(N__25728),
            .I(N__25721));
    InMux I__5298 (
            .O(N__25727),
            .I(N__25718));
    Span4Mux_h I__5297 (
            .O(N__25724),
            .I(N__25715));
    Span4Mux_h I__5296 (
            .O(N__25721),
            .I(N__25712));
    LocalMux I__5295 (
            .O(N__25718),
            .I(\tok.n5_adj_715 ));
    Odrv4 I__5294 (
            .O(N__25715),
            .I(\tok.n5_adj_715 ));
    Odrv4 I__5293 (
            .O(N__25712),
            .I(\tok.n5_adj_715 ));
    CascadeMux I__5292 (
            .O(N__25705),
            .I(\tok.n369_cascade_ ));
    InMux I__5291 (
            .O(N__25702),
            .I(N__25699));
    LocalMux I__5290 (
            .O(N__25699),
            .I(N__25696));
    Span4Mux_v I__5289 (
            .O(N__25696),
            .I(N__25693));
    Odrv4 I__5288 (
            .O(N__25693),
            .I(\tok.n278 ));
    CascadeMux I__5287 (
            .O(N__25690),
            .I(\tok.n233_adj_716_cascade_ ));
    InMux I__5286 (
            .O(N__25687),
            .I(N__25684));
    LocalMux I__5285 (
            .O(N__25684),
            .I(N__25681));
    Span4Mux_s2_h I__5284 (
            .O(N__25681),
            .I(N__25678));
    Span4Mux_v I__5283 (
            .O(N__25678),
            .I(N__25675));
    Odrv4 I__5282 (
            .O(N__25675),
            .I(\tok.n229 ));
    InMux I__5281 (
            .O(N__25672),
            .I(N__25669));
    LocalMux I__5280 (
            .O(N__25669),
            .I(N__25666));
    Span4Mux_h I__5279 (
            .O(N__25666),
            .I(N__25663));
    Odrv4 I__5278 (
            .O(N__25663),
            .I(\tok.n6156 ));
    InMux I__5277 (
            .O(N__25660),
            .I(N__25657));
    LocalMux I__5276 (
            .O(N__25657),
            .I(\tok.n7 ));
    CascadeMux I__5275 (
            .O(N__25654),
            .I(\tok.n53_cascade_ ));
    CEMux I__5274 (
            .O(N__25651),
            .I(N__25646));
    CEMux I__5273 (
            .O(N__25650),
            .I(N__25636));
    CEMux I__5272 (
            .O(N__25649),
            .I(N__25632));
    LocalMux I__5271 (
            .O(N__25646),
            .I(N__25629));
    CEMux I__5270 (
            .O(N__25645),
            .I(N__25626));
    CEMux I__5269 (
            .O(N__25644),
            .I(N__25623));
    CEMux I__5268 (
            .O(N__25643),
            .I(N__25620));
    CEMux I__5267 (
            .O(N__25642),
            .I(N__25617));
    CEMux I__5266 (
            .O(N__25641),
            .I(N__25614));
    CEMux I__5265 (
            .O(N__25640),
            .I(N__25611));
    CEMux I__5264 (
            .O(N__25639),
            .I(N__25608));
    LocalMux I__5263 (
            .O(N__25636),
            .I(N__25604));
    CEMux I__5262 (
            .O(N__25635),
            .I(N__25601));
    LocalMux I__5261 (
            .O(N__25632),
            .I(N__25598));
    Span4Mux_v I__5260 (
            .O(N__25629),
            .I(N__25593));
    LocalMux I__5259 (
            .O(N__25626),
            .I(N__25593));
    LocalMux I__5258 (
            .O(N__25623),
            .I(N__25590));
    LocalMux I__5257 (
            .O(N__25620),
            .I(N__25587));
    LocalMux I__5256 (
            .O(N__25617),
            .I(N__25584));
    LocalMux I__5255 (
            .O(N__25614),
            .I(N__25577));
    LocalMux I__5254 (
            .O(N__25611),
            .I(N__25577));
    LocalMux I__5253 (
            .O(N__25608),
            .I(N__25577));
    CEMux I__5252 (
            .O(N__25607),
            .I(N__25574));
    Span4Mux_v I__5251 (
            .O(N__25604),
            .I(N__25571));
    LocalMux I__5250 (
            .O(N__25601),
            .I(N__25568));
    Span4Mux_h I__5249 (
            .O(N__25598),
            .I(N__25563));
    Span4Mux_h I__5248 (
            .O(N__25593),
            .I(N__25563));
    Span4Mux_v I__5247 (
            .O(N__25590),
            .I(N__25560));
    Span4Mux_h I__5246 (
            .O(N__25587),
            .I(N__25555));
    Span4Mux_h I__5245 (
            .O(N__25584),
            .I(N__25555));
    Span4Mux_v I__5244 (
            .O(N__25577),
            .I(N__25552));
    LocalMux I__5243 (
            .O(N__25574),
            .I(N__25547));
    Span4Mux_h I__5242 (
            .O(N__25571),
            .I(N__25547));
    Span4Mux_h I__5241 (
            .O(N__25568),
            .I(N__25544));
    Span4Mux_s2_h I__5240 (
            .O(N__25563),
            .I(N__25537));
    Span4Mux_h I__5239 (
            .O(N__25560),
            .I(N__25537));
    Span4Mux_h I__5238 (
            .O(N__25555),
            .I(N__25537));
    Span4Mux_h I__5237 (
            .O(N__25552),
            .I(N__25532));
    Span4Mux_v I__5236 (
            .O(N__25547),
            .I(N__25532));
    Sp12to4 I__5235 (
            .O(N__25544),
            .I(N__25527));
    Sp12to4 I__5234 (
            .O(N__25537),
            .I(N__25527));
    Odrv4 I__5233 (
            .O(N__25532),
            .I(\tok.n992 ));
    Odrv12 I__5232 (
            .O(N__25527),
            .I(\tok.n992 ));
    CascadeMux I__5231 (
            .O(N__25522),
            .I(\tok.n2_cascade_ ));
    InMux I__5230 (
            .O(N__25519),
            .I(N__25512));
    InMux I__5229 (
            .O(N__25518),
            .I(N__25507));
    InMux I__5228 (
            .O(N__25517),
            .I(N__25507));
    InMux I__5227 (
            .O(N__25516),
            .I(N__25504));
    InMux I__5226 (
            .O(N__25515),
            .I(N__25501));
    LocalMux I__5225 (
            .O(N__25512),
            .I(N__25494));
    LocalMux I__5224 (
            .O(N__25507),
            .I(N__25494));
    LocalMux I__5223 (
            .O(N__25504),
            .I(N__25489));
    LocalMux I__5222 (
            .O(N__25501),
            .I(N__25489));
    InMux I__5221 (
            .O(N__25500),
            .I(N__25486));
    InMux I__5220 (
            .O(N__25499),
            .I(N__25483));
    Span4Mux_v I__5219 (
            .O(N__25494),
            .I(N__25468));
    Span4Mux_v I__5218 (
            .O(N__25489),
            .I(N__25468));
    LocalMux I__5217 (
            .O(N__25486),
            .I(N__25468));
    LocalMux I__5216 (
            .O(N__25483),
            .I(N__25468));
    InMux I__5215 (
            .O(N__25482),
            .I(N__25463));
    InMux I__5214 (
            .O(N__25481),
            .I(N__25460));
    InMux I__5213 (
            .O(N__25480),
            .I(N__25455));
    InMux I__5212 (
            .O(N__25479),
            .I(N__25455));
    InMux I__5211 (
            .O(N__25478),
            .I(N__25450));
    InMux I__5210 (
            .O(N__25477),
            .I(N__25450));
    Span4Mux_v I__5209 (
            .O(N__25468),
            .I(N__25446));
    InMux I__5208 (
            .O(N__25467),
            .I(N__25441));
    InMux I__5207 (
            .O(N__25466),
            .I(N__25441));
    LocalMux I__5206 (
            .O(N__25463),
            .I(N__25438));
    LocalMux I__5205 (
            .O(N__25460),
            .I(N__25435));
    LocalMux I__5204 (
            .O(N__25455),
            .I(N__25430));
    LocalMux I__5203 (
            .O(N__25450),
            .I(N__25430));
    InMux I__5202 (
            .O(N__25449),
            .I(N__25427));
    Span4Mux_h I__5201 (
            .O(N__25446),
            .I(N__25424));
    LocalMux I__5200 (
            .O(N__25441),
            .I(N__25419));
    Span4Mux_v I__5199 (
            .O(N__25438),
            .I(N__25419));
    Span4Mux_h I__5198 (
            .O(N__25435),
            .I(N__25416));
    Span4Mux_h I__5197 (
            .O(N__25430),
            .I(N__25413));
    LocalMux I__5196 (
            .O(N__25427),
            .I(N__25410));
    Sp12to4 I__5195 (
            .O(N__25424),
            .I(N__25406));
    Span4Mux_h I__5194 (
            .O(N__25419),
            .I(N__25403));
    Span4Mux_s1_h I__5193 (
            .O(N__25416),
            .I(N__25400));
    Span4Mux_v I__5192 (
            .O(N__25413),
            .I(N__25395));
    Span4Mux_h I__5191 (
            .O(N__25410),
            .I(N__25395));
    InMux I__5190 (
            .O(N__25409),
            .I(N__25392));
    Odrv12 I__5189 (
            .O(N__25406),
            .I(\tok.n23 ));
    Odrv4 I__5188 (
            .O(N__25403),
            .I(\tok.n23 ));
    Odrv4 I__5187 (
            .O(N__25400),
            .I(\tok.n23 ));
    Odrv4 I__5186 (
            .O(N__25395),
            .I(\tok.n23 ));
    LocalMux I__5185 (
            .O(N__25392),
            .I(\tok.n23 ));
    CascadeMux I__5184 (
            .O(N__25381),
            .I(\tok.n174_cascade_ ));
    InMux I__5183 (
            .O(N__25378),
            .I(N__25369));
    InMux I__5182 (
            .O(N__25377),
            .I(N__25369));
    InMux I__5181 (
            .O(N__25376),
            .I(N__25364));
    CascadeMux I__5180 (
            .O(N__25375),
            .I(N__25361));
    CascadeMux I__5179 (
            .O(N__25374),
            .I(N__25355));
    LocalMux I__5178 (
            .O(N__25369),
            .I(N__25350));
    InMux I__5177 (
            .O(N__25368),
            .I(N__25347));
    InMux I__5176 (
            .O(N__25367),
            .I(N__25344));
    LocalMux I__5175 (
            .O(N__25364),
            .I(N__25340));
    InMux I__5174 (
            .O(N__25361),
            .I(N__25333));
    InMux I__5173 (
            .O(N__25360),
            .I(N__25333));
    CascadeMux I__5172 (
            .O(N__25359),
            .I(N__25330));
    CascadeMux I__5171 (
            .O(N__25358),
            .I(N__25326));
    InMux I__5170 (
            .O(N__25355),
            .I(N__25320));
    InMux I__5169 (
            .O(N__25354),
            .I(N__25320));
    InMux I__5168 (
            .O(N__25353),
            .I(N__25317));
    Span4Mux_s3_h I__5167 (
            .O(N__25350),
            .I(N__25312));
    LocalMux I__5166 (
            .O(N__25347),
            .I(N__25312));
    LocalMux I__5165 (
            .O(N__25344),
            .I(N__25309));
    InMux I__5164 (
            .O(N__25343),
            .I(N__25306));
    Span4Mux_h I__5163 (
            .O(N__25340),
            .I(N__25303));
    InMux I__5162 (
            .O(N__25339),
            .I(N__25298));
    InMux I__5161 (
            .O(N__25338),
            .I(N__25298));
    LocalMux I__5160 (
            .O(N__25333),
            .I(N__25295));
    InMux I__5159 (
            .O(N__25330),
            .I(N__25290));
    InMux I__5158 (
            .O(N__25329),
            .I(N__25290));
    InMux I__5157 (
            .O(N__25326),
            .I(N__25285));
    InMux I__5156 (
            .O(N__25325),
            .I(N__25285));
    LocalMux I__5155 (
            .O(N__25320),
            .I(N__25282));
    LocalMux I__5154 (
            .O(N__25317),
            .I(N__25275));
    Span4Mux_h I__5153 (
            .O(N__25312),
            .I(N__25275));
    Span4Mux_v I__5152 (
            .O(N__25309),
            .I(N__25275));
    LocalMux I__5151 (
            .O(N__25306),
            .I(N__25270));
    Span4Mux_v I__5150 (
            .O(N__25303),
            .I(N__25270));
    LocalMux I__5149 (
            .O(N__25298),
            .I(\tok.stall ));
    Odrv12 I__5148 (
            .O(N__25295),
            .I(\tok.stall ));
    LocalMux I__5147 (
            .O(N__25290),
            .I(\tok.stall ));
    LocalMux I__5146 (
            .O(N__25285),
            .I(\tok.stall ));
    Odrv4 I__5145 (
            .O(N__25282),
            .I(\tok.stall ));
    Odrv4 I__5144 (
            .O(N__25275),
            .I(\tok.stall ));
    Odrv4 I__5143 (
            .O(N__25270),
            .I(\tok.stall ));
    InMux I__5142 (
            .O(N__25255),
            .I(N__25249));
    InMux I__5141 (
            .O(N__25254),
            .I(N__25249));
    LocalMux I__5140 (
            .O(N__25249),
            .I(N__25244));
    InMux I__5139 (
            .O(N__25248),
            .I(N__25239));
    InMux I__5138 (
            .O(N__25247),
            .I(N__25239));
    Span4Mux_v I__5137 (
            .O(N__25244),
            .I(N__25235));
    LocalMux I__5136 (
            .O(N__25239),
            .I(N__25232));
    InMux I__5135 (
            .O(N__25238),
            .I(N__25229));
    Sp12to4 I__5134 (
            .O(N__25235),
            .I(N__25226));
    Span4Mux_v I__5133 (
            .O(N__25232),
            .I(N__25221));
    LocalMux I__5132 (
            .O(N__25229),
            .I(N__25221));
    Odrv12 I__5131 (
            .O(N__25226),
            .I(\tok.n6189 ));
    Odrv4 I__5130 (
            .O(N__25221),
            .I(\tok.n6189 ));
    InMux I__5129 (
            .O(N__25216),
            .I(N__25213));
    LocalMux I__5128 (
            .O(N__25213),
            .I(\tok.n6_adj_722 ));
    InMux I__5127 (
            .O(N__25210),
            .I(N__25206));
    InMux I__5126 (
            .O(N__25209),
            .I(N__25203));
    LocalMux I__5125 (
            .O(N__25206),
            .I(N__25200));
    LocalMux I__5124 (
            .O(N__25203),
            .I(tail_49_adj_899));
    Odrv12 I__5123 (
            .O(N__25200),
            .I(tail_49_adj_899));
    InMux I__5122 (
            .O(N__25195),
            .I(N__25189));
    InMux I__5121 (
            .O(N__25194),
            .I(N__25189));
    LocalMux I__5120 (
            .O(N__25189),
            .I(\tok.C_stk.tail_33 ));
    InMux I__5119 (
            .O(N__25186),
            .I(N__25182));
    InMux I__5118 (
            .O(N__25185),
            .I(N__25179));
    LocalMux I__5117 (
            .O(N__25182),
            .I(N__25176));
    LocalMux I__5116 (
            .O(N__25179),
            .I(tail_41));
    Odrv4 I__5115 (
            .O(N__25176),
            .I(tail_41));
    InMux I__5114 (
            .O(N__25171),
            .I(N__25168));
    LocalMux I__5113 (
            .O(N__25168),
            .I(\tok.n156 ));
    CascadeMux I__5112 (
            .O(N__25165),
            .I(\tok.n211_adj_741_cascade_ ));
    CascadeMux I__5111 (
            .O(N__25162),
            .I(\tok.n277_cascade_ ));
    InMux I__5110 (
            .O(N__25159),
            .I(N__25156));
    LocalMux I__5109 (
            .O(N__25156),
            .I(\tok.n265 ));
    InMux I__5108 (
            .O(N__25153),
            .I(N__25150));
    LocalMux I__5107 (
            .O(N__25150),
            .I(N__25147));
    Span4Mux_h I__5106 (
            .O(N__25147),
            .I(N__25144));
    Span4Mux_h I__5105 (
            .O(N__25144),
            .I(N__25141));
    Odrv4 I__5104 (
            .O(N__25141),
            .I(\tok.n6_adj_748 ));
    CascadeMux I__5103 (
            .O(N__25138),
            .I(N__25135));
    InMux I__5102 (
            .O(N__25135),
            .I(N__25132));
    LocalMux I__5101 (
            .O(N__25132),
            .I(N__25129));
    Span4Mux_h I__5100 (
            .O(N__25129),
            .I(N__25126));
    Odrv4 I__5099 (
            .O(N__25126),
            .I(\tok.n6331 ));
    CascadeMux I__5098 (
            .O(N__25123),
            .I(\tok.n238_adj_855_cascade_ ));
    InMux I__5097 (
            .O(N__25120),
            .I(N__25117));
    LocalMux I__5096 (
            .O(N__25117),
            .I(N__25114));
    Odrv12 I__5095 (
            .O(N__25114),
            .I(\tok.n4_adj_859 ));
    CascadeMux I__5094 (
            .O(N__25111),
            .I(N__25107));
    CascadeMux I__5093 (
            .O(N__25110),
            .I(N__25103));
    InMux I__5092 (
            .O(N__25107),
            .I(N__25100));
    InMux I__5091 (
            .O(N__25106),
            .I(N__25097));
    InMux I__5090 (
            .O(N__25103),
            .I(N__25094));
    LocalMux I__5089 (
            .O(N__25100),
            .I(N__25091));
    LocalMux I__5088 (
            .O(N__25097),
            .I(N__25088));
    LocalMux I__5087 (
            .O(N__25094),
            .I(N__25083));
    Span4Mux_s3_h I__5086 (
            .O(N__25091),
            .I(N__25083));
    Span4Mux_h I__5085 (
            .O(N__25088),
            .I(N__25080));
    Odrv4 I__5084 (
            .O(N__25083),
            .I(\tok.n6_adj_676 ));
    Odrv4 I__5083 (
            .O(N__25080),
            .I(\tok.n6_adj_676 ));
    InMux I__5082 (
            .O(N__25075),
            .I(N__25072));
    LocalMux I__5081 (
            .O(N__25072),
            .I(\tok.n298_adj_856 ));
    InMux I__5080 (
            .O(N__25069),
            .I(N__25063));
    InMux I__5079 (
            .O(N__25068),
            .I(N__25063));
    LocalMux I__5078 (
            .O(N__25063),
            .I(N__25060));
    Span4Mux_h I__5077 (
            .O(N__25060),
            .I(N__25057));
    Sp12to4 I__5076 (
            .O(N__25057),
            .I(N__25054));
    Odrv12 I__5075 (
            .O(N__25054),
            .I(\tok.n37 ));
    InMux I__5074 (
            .O(N__25051),
            .I(N__25045));
    InMux I__5073 (
            .O(N__25050),
            .I(N__25045));
    LocalMux I__5072 (
            .O(N__25045),
            .I(N__25042));
    Span4Mux_v I__5071 (
            .O(N__25042),
            .I(N__25039));
    Sp12to4 I__5070 (
            .O(N__25039),
            .I(N__25036));
    Odrv12 I__5069 (
            .O(N__25036),
            .I(\tok.n2559 ));
    InMux I__5068 (
            .O(N__25033),
            .I(N__25030));
    LocalMux I__5067 (
            .O(N__25030),
            .I(N__25026));
    InMux I__5066 (
            .O(N__25029),
            .I(N__25023));
    Span4Mux_h I__5065 (
            .O(N__25026),
            .I(N__25018));
    LocalMux I__5064 (
            .O(N__25023),
            .I(N__25018));
    Odrv4 I__5063 (
            .O(N__25018),
            .I(\tok.tail_53 ));
    CascadeMux I__5062 (
            .O(N__25015),
            .I(rd_7__N_373_cascade_));
    InMux I__5061 (
            .O(N__25012),
            .I(N__25008));
    InMux I__5060 (
            .O(N__25011),
            .I(N__25005));
    LocalMux I__5059 (
            .O(N__25008),
            .I(\tok.tail_61 ));
    LocalMux I__5058 (
            .O(N__25005),
            .I(\tok.tail_61 ));
    InMux I__5057 (
            .O(N__25000),
            .I(N__24997));
    LocalMux I__5056 (
            .O(N__24997),
            .I(N__24992));
    InMux I__5055 (
            .O(N__24996),
            .I(N__24987));
    InMux I__5054 (
            .O(N__24995),
            .I(N__24987));
    Span4Mux_s3_h I__5053 (
            .O(N__24992),
            .I(N__24981));
    LocalMux I__5052 (
            .O(N__24987),
            .I(N__24981));
    InMux I__5051 (
            .O(N__24986),
            .I(N__24978));
    Span4Mux_h I__5050 (
            .O(N__24981),
            .I(N__24975));
    LocalMux I__5049 (
            .O(N__24978),
            .I(tc_plus_1_1));
    Odrv4 I__5048 (
            .O(N__24975),
            .I(tc_plus_1_1));
    CascadeMux I__5047 (
            .O(N__24970),
            .I(\tok.C_stk.n6248_cascade_ ));
    InMux I__5046 (
            .O(N__24967),
            .I(N__24964));
    LocalMux I__5045 (
            .O(N__24964),
            .I(N__24960));
    InMux I__5044 (
            .O(N__24963),
            .I(N__24956));
    Span4Mux_v I__5043 (
            .O(N__24960),
            .I(N__24952));
    InMux I__5042 (
            .O(N__24959),
            .I(N__24949));
    LocalMux I__5041 (
            .O(N__24956),
            .I(N__24946));
    InMux I__5040 (
            .O(N__24955),
            .I(N__24943));
    Odrv4 I__5039 (
            .O(N__24952),
            .I(tc_1));
    LocalMux I__5038 (
            .O(N__24949),
            .I(tc_1));
    Odrv12 I__5037 (
            .O(N__24946),
            .I(tc_1));
    LocalMux I__5036 (
            .O(N__24943),
            .I(tc_1));
    CascadeMux I__5035 (
            .O(N__24934),
            .I(N__24930));
    InMux I__5034 (
            .O(N__24933),
            .I(N__24921));
    InMux I__5033 (
            .O(N__24930),
            .I(N__24921));
    InMux I__5032 (
            .O(N__24929),
            .I(N__24921));
    InMux I__5031 (
            .O(N__24928),
            .I(N__24918));
    LocalMux I__5030 (
            .O(N__24921),
            .I(N__24915));
    LocalMux I__5029 (
            .O(N__24918),
            .I(c_stk_r_1));
    Odrv4 I__5028 (
            .O(N__24915),
            .I(c_stk_r_1));
    InMux I__5027 (
            .O(N__24910),
            .I(N__24904));
    InMux I__5026 (
            .O(N__24909),
            .I(N__24904));
    LocalMux I__5025 (
            .O(N__24904),
            .I(\tok.C_stk.tail_1 ));
    InMux I__5024 (
            .O(N__24901),
            .I(N__24895));
    InMux I__5023 (
            .O(N__24900),
            .I(N__24895));
    LocalMux I__5022 (
            .O(N__24895),
            .I(tail_9));
    CascadeMux I__5021 (
            .O(N__24892),
            .I(N__24889));
    InMux I__5020 (
            .O(N__24889),
            .I(N__24883));
    InMux I__5019 (
            .O(N__24888),
            .I(N__24883));
    LocalMux I__5018 (
            .O(N__24883),
            .I(\tok.C_stk.tail_17 ));
    InMux I__5017 (
            .O(N__24880),
            .I(N__24874));
    InMux I__5016 (
            .O(N__24879),
            .I(N__24874));
    LocalMux I__5015 (
            .O(N__24874),
            .I(tail_25));
    InMux I__5014 (
            .O(N__24871),
            .I(N__24867));
    InMux I__5013 (
            .O(N__24870),
            .I(N__24864));
    LocalMux I__5012 (
            .O(N__24867),
            .I(N__24861));
    LocalMux I__5011 (
            .O(N__24864),
            .I(\tok.tail_44 ));
    Odrv12 I__5010 (
            .O(N__24861),
            .I(\tok.tail_44 ));
    InMux I__5009 (
            .O(N__24856),
            .I(N__24852));
    InMux I__5008 (
            .O(N__24855),
            .I(N__24849));
    LocalMux I__5007 (
            .O(N__24852),
            .I(N__24844));
    LocalMux I__5006 (
            .O(N__24849),
            .I(N__24844));
    Odrv4 I__5005 (
            .O(N__24844),
            .I(\tok.tail_42 ));
    CascadeMux I__5004 (
            .O(N__24841),
            .I(N__24837));
    InMux I__5003 (
            .O(N__24840),
            .I(N__24834));
    InMux I__5002 (
            .O(N__24837),
            .I(N__24831));
    LocalMux I__5001 (
            .O(N__24834),
            .I(N__24828));
    LocalMux I__5000 (
            .O(N__24831),
            .I(N__24825));
    Span4Mux_v I__4999 (
            .O(N__24828),
            .I(N__24822));
    Odrv4 I__4998 (
            .O(N__24825),
            .I(tail_51));
    Odrv4 I__4997 (
            .O(N__24822),
            .I(tail_51));
    InMux I__4996 (
            .O(N__24817),
            .I(N__24813));
    InMux I__4995 (
            .O(N__24816),
            .I(N__24810));
    LocalMux I__4994 (
            .O(N__24813),
            .I(tail_59));
    LocalMux I__4993 (
            .O(N__24810),
            .I(tail_59));
    CascadeMux I__4992 (
            .O(N__24805),
            .I(N__24802));
    InMux I__4991 (
            .O(N__24802),
            .I(N__24798));
    InMux I__4990 (
            .O(N__24801),
            .I(N__24795));
    LocalMux I__4989 (
            .O(N__24798),
            .I(N__24792));
    LocalMux I__4988 (
            .O(N__24795),
            .I(N__24789));
    Odrv4 I__4987 (
            .O(N__24792),
            .I(tail_48_adj_900));
    Odrv4 I__4986 (
            .O(N__24789),
            .I(tail_48_adj_900));
    InMux I__4985 (
            .O(N__24784),
            .I(N__24781));
    LocalMux I__4984 (
            .O(N__24781),
            .I(N__24777));
    InMux I__4983 (
            .O(N__24780),
            .I(N__24774));
    Odrv4 I__4982 (
            .O(N__24777),
            .I(tail_56));
    LocalMux I__4981 (
            .O(N__24774),
            .I(tail_56));
    CascadeMux I__4980 (
            .O(N__24769),
            .I(C_stk_delta_1_cascade_));
    InMux I__4979 (
            .O(N__24766),
            .I(N__24763));
    LocalMux I__4978 (
            .O(N__24763),
            .I(N__24759));
    InMux I__4977 (
            .O(N__24762),
            .I(N__24756));
    Odrv12 I__4976 (
            .O(N__24759),
            .I(tail_57));
    LocalMux I__4975 (
            .O(N__24756),
            .I(tail_57));
    InMux I__4974 (
            .O(N__24751),
            .I(N__24747));
    CascadeMux I__4973 (
            .O(N__24750),
            .I(N__24744));
    LocalMux I__4972 (
            .O(N__24747),
            .I(N__24741));
    InMux I__4971 (
            .O(N__24744),
            .I(N__24738));
    Odrv12 I__4970 (
            .O(N__24741),
            .I(\tok.tail_52 ));
    LocalMux I__4969 (
            .O(N__24738),
            .I(\tok.tail_52 ));
    InMux I__4968 (
            .O(N__24733),
            .I(N__24729));
    InMux I__4967 (
            .O(N__24732),
            .I(N__24726));
    LocalMux I__4966 (
            .O(N__24729),
            .I(\tok.tail_60 ));
    LocalMux I__4965 (
            .O(N__24726),
            .I(\tok.tail_60 ));
    InMux I__4964 (
            .O(N__24721),
            .I(N__24718));
    LocalMux I__4963 (
            .O(N__24718),
            .I(N__24714));
    InMux I__4962 (
            .O(N__24717),
            .I(N__24711));
    Odrv12 I__4961 (
            .O(N__24714),
            .I(\tok.tail_62 ));
    LocalMux I__4960 (
            .O(N__24711),
            .I(\tok.tail_62 ));
    InMux I__4959 (
            .O(N__24706),
            .I(N__24700));
    InMux I__4958 (
            .O(N__24705),
            .I(N__24700));
    LocalMux I__4957 (
            .O(N__24700),
            .I(tail_40));
    InMux I__4956 (
            .O(N__24697),
            .I(N__24693));
    InMux I__4955 (
            .O(N__24696),
            .I(N__24690));
    LocalMux I__4954 (
            .O(N__24693),
            .I(N__24687));
    LocalMux I__4953 (
            .O(N__24690),
            .I(tail_8));
    Odrv4 I__4952 (
            .O(N__24687),
            .I(tail_8));
    InMux I__4951 (
            .O(N__24682),
            .I(N__24678));
    InMux I__4950 (
            .O(N__24681),
            .I(N__24675));
    LocalMux I__4949 (
            .O(N__24678),
            .I(\tok.C_stk.tail_32 ));
    LocalMux I__4948 (
            .O(N__24675),
            .I(\tok.C_stk.tail_32 ));
    InMux I__4947 (
            .O(N__24670),
            .I(N__24667));
    LocalMux I__4946 (
            .O(N__24667),
            .I(N__24664));
    Span4Mux_h I__4945 (
            .O(N__24664),
            .I(N__24660));
    InMux I__4944 (
            .O(N__24663),
            .I(N__24657));
    Odrv4 I__4943 (
            .O(N__24660),
            .I(\tok.C_stk.tail_16 ));
    LocalMux I__4942 (
            .O(N__24657),
            .I(\tok.C_stk.tail_16 ));
    InMux I__4941 (
            .O(N__24652),
            .I(N__24648));
    InMux I__4940 (
            .O(N__24651),
            .I(N__24645));
    LocalMux I__4939 (
            .O(N__24648),
            .I(tail_24));
    LocalMux I__4938 (
            .O(N__24645),
            .I(tail_24));
    InMux I__4937 (
            .O(N__24640),
            .I(N__24637));
    LocalMux I__4936 (
            .O(N__24637),
            .I(N__24633));
    InMux I__4935 (
            .O(N__24636),
            .I(N__24630));
    Span4Mux_s3_h I__4934 (
            .O(N__24633),
            .I(N__24627));
    LocalMux I__4933 (
            .O(N__24630),
            .I(\tok.C_stk.tail_43 ));
    Odrv4 I__4932 (
            .O(N__24627),
            .I(\tok.C_stk.tail_43 ));
    InMux I__4931 (
            .O(N__24622),
            .I(N__24619));
    LocalMux I__4930 (
            .O(N__24619),
            .I(N__24615));
    InMux I__4929 (
            .O(N__24618),
            .I(N__24612));
    Span4Mux_s3_h I__4928 (
            .O(N__24615),
            .I(N__24609));
    LocalMux I__4927 (
            .O(N__24612),
            .I(\tok.tail_45 ));
    Odrv4 I__4926 (
            .O(N__24609),
            .I(\tok.tail_45 ));
    InMux I__4925 (
            .O(N__24604),
            .I(N__24601));
    LocalMux I__4924 (
            .O(N__24601),
            .I(\tok.n6442 ));
    CascadeMux I__4923 (
            .O(N__24598),
            .I(\tok.n6433_cascade_ ));
    InMux I__4922 (
            .O(N__24595),
            .I(N__24592));
    LocalMux I__4921 (
            .O(N__24592),
            .I(N__24589));
    Span4Mux_h I__4920 (
            .O(N__24589),
            .I(N__24586));
    Odrv4 I__4919 (
            .O(N__24586),
            .I(\tok.n215_adj_841 ));
    InMux I__4918 (
            .O(N__24583),
            .I(N__24580));
    LocalMux I__4917 (
            .O(N__24580),
            .I(\tok.n179_adj_842 ));
    CascadeMux I__4916 (
            .O(N__24577),
            .I(\tok.n6602_cascade_ ));
    InMux I__4915 (
            .O(N__24574),
            .I(N__24571));
    LocalMux I__4914 (
            .O(N__24571),
            .I(N__24568));
    Odrv4 I__4913 (
            .O(N__24568),
            .I(\tok.n6601 ));
    InMux I__4912 (
            .O(N__24565),
            .I(N__24562));
    LocalMux I__4911 (
            .O(N__24562),
            .I(N__24559));
    Odrv4 I__4910 (
            .O(N__24559),
            .I(\tok.n6375 ));
    InMux I__4909 (
            .O(N__24556),
            .I(N__24548));
    CascadeMux I__4908 (
            .O(N__24555),
            .I(N__24545));
    CascadeMux I__4907 (
            .O(N__24554),
            .I(N__24542));
    CascadeMux I__4906 (
            .O(N__24553),
            .I(N__24537));
    CascadeMux I__4905 (
            .O(N__24552),
            .I(N__24534));
    CascadeMux I__4904 (
            .O(N__24551),
            .I(N__24531));
    LocalMux I__4903 (
            .O(N__24548),
            .I(N__24528));
    InMux I__4902 (
            .O(N__24545),
            .I(N__24525));
    InMux I__4901 (
            .O(N__24542),
            .I(N__24518));
    InMux I__4900 (
            .O(N__24541),
            .I(N__24518));
    InMux I__4899 (
            .O(N__24540),
            .I(N__24518));
    InMux I__4898 (
            .O(N__24537),
            .I(N__24515));
    InMux I__4897 (
            .O(N__24534),
            .I(N__24512));
    InMux I__4896 (
            .O(N__24531),
            .I(N__24509));
    Span4Mux_v I__4895 (
            .O(N__24528),
            .I(N__24502));
    LocalMux I__4894 (
            .O(N__24525),
            .I(N__24502));
    LocalMux I__4893 (
            .O(N__24518),
            .I(N__24502));
    LocalMux I__4892 (
            .O(N__24515),
            .I(\tok.n847 ));
    LocalMux I__4891 (
            .O(N__24512),
            .I(\tok.n847 ));
    LocalMux I__4890 (
            .O(N__24509),
            .I(\tok.n847 ));
    Odrv4 I__4889 (
            .O(N__24502),
            .I(\tok.n847 ));
    InMux I__4888 (
            .O(N__24493),
            .I(N__24490));
    LocalMux I__4887 (
            .O(N__24490),
            .I(\tok.n6544 ));
    CascadeMux I__4886 (
            .O(N__24487),
            .I(\tok.n179_adj_657_cascade_ ));
    InMux I__4885 (
            .O(N__24484),
            .I(N__24481));
    LocalMux I__4884 (
            .O(N__24481),
            .I(N__24478));
    Span4Mux_h I__4883 (
            .O(N__24478),
            .I(N__24475));
    Odrv4 I__4882 (
            .O(N__24475),
            .I(\tok.n6543 ));
    InMux I__4881 (
            .O(N__24472),
            .I(N__24469));
    LocalMux I__4880 (
            .O(N__24469),
            .I(N__24466));
    Odrv12 I__4879 (
            .O(N__24466),
            .I(\tok.n464 ));
    CascadeMux I__4878 (
            .O(N__24463),
            .I(N__24455));
    CascadeMux I__4877 (
            .O(N__24462),
            .I(N__24449));
    CascadeMux I__4876 (
            .O(N__24461),
            .I(N__24445));
    CascadeMux I__4875 (
            .O(N__24460),
            .I(N__24442));
    CascadeMux I__4874 (
            .O(N__24459),
            .I(N__24438));
    CascadeMux I__4873 (
            .O(N__24458),
            .I(N__24434));
    InMux I__4872 (
            .O(N__24455),
            .I(N__24430));
    InMux I__4871 (
            .O(N__24454),
            .I(N__24427));
    CascadeMux I__4870 (
            .O(N__24453),
            .I(N__24422));
    InMux I__4869 (
            .O(N__24452),
            .I(N__24413));
    InMux I__4868 (
            .O(N__24449),
            .I(N__24413));
    InMux I__4867 (
            .O(N__24448),
            .I(N__24413));
    InMux I__4866 (
            .O(N__24445),
            .I(N__24413));
    InMux I__4865 (
            .O(N__24442),
            .I(N__24410));
    InMux I__4864 (
            .O(N__24441),
            .I(N__24405));
    InMux I__4863 (
            .O(N__24438),
            .I(N__24405));
    CascadeMux I__4862 (
            .O(N__24437),
            .I(N__24402));
    InMux I__4861 (
            .O(N__24434),
            .I(N__24399));
    CascadeMux I__4860 (
            .O(N__24433),
            .I(N__24396));
    LocalMux I__4859 (
            .O(N__24430),
            .I(N__24391));
    LocalMux I__4858 (
            .O(N__24427),
            .I(N__24391));
    InMux I__4857 (
            .O(N__24426),
            .I(N__24384));
    InMux I__4856 (
            .O(N__24425),
            .I(N__24384));
    InMux I__4855 (
            .O(N__24422),
            .I(N__24384));
    LocalMux I__4854 (
            .O(N__24413),
            .I(N__24379));
    LocalMux I__4853 (
            .O(N__24410),
            .I(N__24379));
    LocalMux I__4852 (
            .O(N__24405),
            .I(N__24376));
    InMux I__4851 (
            .O(N__24402),
            .I(N__24373));
    LocalMux I__4850 (
            .O(N__24399),
            .I(N__24370));
    InMux I__4849 (
            .O(N__24396),
            .I(N__24367));
    Span4Mux_h I__4848 (
            .O(N__24391),
            .I(N__24362));
    LocalMux I__4847 (
            .O(N__24384),
            .I(N__24362));
    Span4Mux_v I__4846 (
            .O(N__24379),
            .I(N__24359));
    Span4Mux_h I__4845 (
            .O(N__24376),
            .I(N__24356));
    LocalMux I__4844 (
            .O(N__24373),
            .I(\tok.n8 ));
    Odrv4 I__4843 (
            .O(N__24370),
            .I(\tok.n8 ));
    LocalMux I__4842 (
            .O(N__24367),
            .I(\tok.n8 ));
    Odrv4 I__4841 (
            .O(N__24362),
            .I(\tok.n8 ));
    Odrv4 I__4840 (
            .O(N__24359),
            .I(\tok.n8 ));
    Odrv4 I__4839 (
            .O(N__24356),
            .I(\tok.n8 ));
    InMux I__4838 (
            .O(N__24343),
            .I(N__24340));
    LocalMux I__4837 (
            .O(N__24340),
            .I(\tok.n6382 ));
    CascadeMux I__4836 (
            .O(N__24337),
            .I(N__24334));
    InMux I__4835 (
            .O(N__24334),
            .I(N__24330));
    InMux I__4834 (
            .O(N__24333),
            .I(N__24325));
    LocalMux I__4833 (
            .O(N__24330),
            .I(N__24319));
    InMux I__4832 (
            .O(N__24329),
            .I(N__24314));
    InMux I__4831 (
            .O(N__24328),
            .I(N__24311));
    LocalMux I__4830 (
            .O(N__24325),
            .I(N__24308));
    InMux I__4829 (
            .O(N__24324),
            .I(N__24305));
    InMux I__4828 (
            .O(N__24323),
            .I(N__24300));
    InMux I__4827 (
            .O(N__24322),
            .I(N__24300));
    Span4Mux_v I__4826 (
            .O(N__24319),
            .I(N__24297));
    InMux I__4825 (
            .O(N__24318),
            .I(N__24294));
    CascadeMux I__4824 (
            .O(N__24317),
            .I(N__24291));
    LocalMux I__4823 (
            .O(N__24314),
            .I(N__24284));
    LocalMux I__4822 (
            .O(N__24311),
            .I(N__24279));
    Span4Mux_v I__4821 (
            .O(N__24308),
            .I(N__24279));
    LocalMux I__4820 (
            .O(N__24305),
            .I(N__24274));
    LocalMux I__4819 (
            .O(N__24300),
            .I(N__24274));
    Sp12to4 I__4818 (
            .O(N__24297),
            .I(N__24269));
    LocalMux I__4817 (
            .O(N__24294),
            .I(N__24269));
    InMux I__4816 (
            .O(N__24291),
            .I(N__24266));
    InMux I__4815 (
            .O(N__24290),
            .I(N__24259));
    InMux I__4814 (
            .O(N__24289),
            .I(N__24259));
    InMux I__4813 (
            .O(N__24288),
            .I(N__24259));
    InMux I__4812 (
            .O(N__24287),
            .I(N__24256));
    Span4Mux_s2_v I__4811 (
            .O(N__24284),
            .I(N__24249));
    Span4Mux_s2_v I__4810 (
            .O(N__24279),
            .I(N__24249));
    Span4Mux_v I__4809 (
            .O(N__24274),
            .I(N__24249));
    Span12Mux_h I__4808 (
            .O(N__24269),
            .I(N__24246));
    LocalMux I__4807 (
            .O(N__24266),
            .I(N__24237));
    LocalMux I__4806 (
            .O(N__24259),
            .I(N__24237));
    LocalMux I__4805 (
            .O(N__24256),
            .I(N__24237));
    Sp12to4 I__4804 (
            .O(N__24249),
            .I(N__24237));
    Odrv12 I__4803 (
            .O(N__24246),
            .I(\tok.n4_adj_636 ));
    Odrv12 I__4802 (
            .O(N__24237),
            .I(\tok.n4_adj_636 ));
    InMux I__4801 (
            .O(N__24232),
            .I(N__24229));
    LocalMux I__4800 (
            .O(N__24229),
            .I(\tok.n213_adj_795 ));
    CascadeMux I__4799 (
            .O(N__24226),
            .I(\tok.n207_adj_796_cascade_ ));
    InMux I__4798 (
            .O(N__24223),
            .I(N__24220));
    LocalMux I__4797 (
            .O(N__24220),
            .I(N__24215));
    InMux I__4796 (
            .O(N__24219),
            .I(N__24210));
    InMux I__4795 (
            .O(N__24218),
            .I(N__24210));
    Span4Mux_s3_v I__4794 (
            .O(N__24215),
            .I(N__24205));
    LocalMux I__4793 (
            .O(N__24210),
            .I(N__24205));
    Odrv4 I__4792 (
            .O(N__24205),
            .I(\tok.n872 ));
    CascadeMux I__4791 (
            .O(N__24202),
            .I(\tok.n6505_cascade_ ));
    CascadeMux I__4790 (
            .O(N__24199),
            .I(N__24193));
    InMux I__4789 (
            .O(N__24198),
            .I(N__24190));
    CascadeMux I__4788 (
            .O(N__24197),
            .I(N__24187));
    InMux I__4787 (
            .O(N__24196),
            .I(N__24181));
    InMux I__4786 (
            .O(N__24193),
            .I(N__24176));
    LocalMux I__4785 (
            .O(N__24190),
            .I(N__24173));
    InMux I__4784 (
            .O(N__24187),
            .I(N__24170));
    InMux I__4783 (
            .O(N__24186),
            .I(N__24166));
    InMux I__4782 (
            .O(N__24185),
            .I(N__24161));
    InMux I__4781 (
            .O(N__24184),
            .I(N__24161));
    LocalMux I__4780 (
            .O(N__24181),
            .I(N__24158));
    CascadeMux I__4779 (
            .O(N__24180),
            .I(N__24155));
    InMux I__4778 (
            .O(N__24179),
            .I(N__24152));
    LocalMux I__4777 (
            .O(N__24176),
            .I(N__24149));
    Span4Mux_v I__4776 (
            .O(N__24173),
            .I(N__24144));
    LocalMux I__4775 (
            .O(N__24170),
            .I(N__24144));
    InMux I__4774 (
            .O(N__24169),
            .I(N__24140));
    LocalMux I__4773 (
            .O(N__24166),
            .I(N__24137));
    LocalMux I__4772 (
            .O(N__24161),
            .I(N__24134));
    Span4Mux_v I__4771 (
            .O(N__24158),
            .I(N__24130));
    InMux I__4770 (
            .O(N__24155),
            .I(N__24127));
    LocalMux I__4769 (
            .O(N__24152),
            .I(N__24124));
    Span4Mux_v I__4768 (
            .O(N__24149),
            .I(N__24119));
    Span4Mux_s1_h I__4767 (
            .O(N__24144),
            .I(N__24119));
    InMux I__4766 (
            .O(N__24143),
            .I(N__24116));
    LocalMux I__4765 (
            .O(N__24140),
            .I(N__24113));
    Span4Mux_h I__4764 (
            .O(N__24137),
            .I(N__24108));
    Span4Mux_h I__4763 (
            .O(N__24134),
            .I(N__24108));
    InMux I__4762 (
            .O(N__24133),
            .I(N__24105));
    Span4Mux_v I__4761 (
            .O(N__24130),
            .I(N__24102));
    LocalMux I__4760 (
            .O(N__24127),
            .I(N__24099));
    Span4Mux_h I__4759 (
            .O(N__24124),
            .I(N__24094));
    Span4Mux_h I__4758 (
            .O(N__24119),
            .I(N__24094));
    LocalMux I__4757 (
            .O(N__24116),
            .I(N__24091));
    Span4Mux_h I__4756 (
            .O(N__24113),
            .I(N__24086));
    Span4Mux_v I__4755 (
            .O(N__24108),
            .I(N__24086));
    LocalMux I__4754 (
            .O(N__24105),
            .I(\tok.n42 ));
    Odrv4 I__4753 (
            .O(N__24102),
            .I(\tok.n42 ));
    Odrv12 I__4752 (
            .O(N__24099),
            .I(\tok.n42 ));
    Odrv4 I__4751 (
            .O(N__24094),
            .I(\tok.n42 ));
    Odrv12 I__4750 (
            .O(N__24091),
            .I(\tok.n42 ));
    Odrv4 I__4749 (
            .O(N__24086),
            .I(\tok.n42 ));
    InMux I__4748 (
            .O(N__24073),
            .I(N__24070));
    LocalMux I__4747 (
            .O(N__24070),
            .I(N__24067));
    Span4Mux_s2_v I__4746 (
            .O(N__24067),
            .I(N__24064));
    Odrv4 I__4745 (
            .O(N__24064),
            .I(\tok.n6360 ));
    CascadeMux I__4744 (
            .O(N__24061),
            .I(N__24057));
    CascadeMux I__4743 (
            .O(N__24060),
            .I(N__24054));
    InMux I__4742 (
            .O(N__24057),
            .I(N__24051));
    InMux I__4741 (
            .O(N__24054),
            .I(N__24048));
    LocalMux I__4740 (
            .O(N__24051),
            .I(N__24045));
    LocalMux I__4739 (
            .O(N__24048),
            .I(N__24042));
    Span4Mux_v I__4738 (
            .O(N__24045),
            .I(N__24039));
    Span4Mux_v I__4737 (
            .O(N__24042),
            .I(N__24036));
    Span4Mux_h I__4736 (
            .O(N__24039),
            .I(N__24031));
    Span4Mux_v I__4735 (
            .O(N__24036),
            .I(N__24031));
    Odrv4 I__4734 (
            .O(N__24031),
            .I(\tok.table_rd_6 ));
    InMux I__4733 (
            .O(N__24028),
            .I(N__24025));
    LocalMux I__4732 (
            .O(N__24025),
            .I(N__24022));
    Odrv4 I__4731 (
            .O(N__24022),
            .I(\tok.n210_adj_802 ));
    CascadeMux I__4730 (
            .O(N__24019),
            .I(N__24016));
    InMux I__4729 (
            .O(N__24016),
            .I(N__24013));
    LocalMux I__4728 (
            .O(N__24013),
            .I(N__24010));
    Span4Mux_h I__4727 (
            .O(N__24010),
            .I(N__24007));
    Odrv4 I__4726 (
            .O(N__24007),
            .I(\tok.n316 ));
    CascadeMux I__4725 (
            .O(N__24004),
            .I(\tok.n6409_cascade_ ));
    InMux I__4724 (
            .O(N__24001),
            .I(N__23996));
    InMux I__4723 (
            .O(N__24000),
            .I(N__23989));
    InMux I__4722 (
            .O(N__23999),
            .I(N__23984));
    LocalMux I__4721 (
            .O(N__23996),
            .I(N__23981));
    InMux I__4720 (
            .O(N__23995),
            .I(N__23978));
    InMux I__4719 (
            .O(N__23994),
            .I(N__23975));
    InMux I__4718 (
            .O(N__23993),
            .I(N__23972));
    InMux I__4717 (
            .O(N__23992),
            .I(N__23969));
    LocalMux I__4716 (
            .O(N__23989),
            .I(N__23962));
    InMux I__4715 (
            .O(N__23988),
            .I(N__23957));
    InMux I__4714 (
            .O(N__23987),
            .I(N__23957));
    LocalMux I__4713 (
            .O(N__23984),
            .I(N__23954));
    Span4Mux_v I__4712 (
            .O(N__23981),
            .I(N__23945));
    LocalMux I__4711 (
            .O(N__23978),
            .I(N__23945));
    LocalMux I__4710 (
            .O(N__23975),
            .I(N__23945));
    LocalMux I__4709 (
            .O(N__23972),
            .I(N__23942));
    LocalMux I__4708 (
            .O(N__23969),
            .I(N__23939));
    InMux I__4707 (
            .O(N__23968),
            .I(N__23936));
    InMux I__4706 (
            .O(N__23967),
            .I(N__23929));
    InMux I__4705 (
            .O(N__23966),
            .I(N__23929));
    InMux I__4704 (
            .O(N__23965),
            .I(N__23929));
    Span12Mux_v I__4703 (
            .O(N__23962),
            .I(N__23926));
    LocalMux I__4702 (
            .O(N__23957),
            .I(N__23921));
    Span4Mux_v I__4701 (
            .O(N__23954),
            .I(N__23921));
    InMux I__4700 (
            .O(N__23953),
            .I(N__23916));
    InMux I__4699 (
            .O(N__23952),
            .I(N__23916));
    Span4Mux_v I__4698 (
            .O(N__23945),
            .I(N__23913));
    Span4Mux_v I__4697 (
            .O(N__23942),
            .I(N__23906));
    Span4Mux_h I__4696 (
            .O(N__23939),
            .I(N__23906));
    LocalMux I__4695 (
            .O(N__23936),
            .I(N__23906));
    LocalMux I__4694 (
            .O(N__23929),
            .I(N__23903));
    Odrv12 I__4693 (
            .O(N__23926),
            .I(\tok.n46 ));
    Odrv4 I__4692 (
            .O(N__23921),
            .I(\tok.n46 ));
    LocalMux I__4691 (
            .O(N__23916),
            .I(\tok.n46 ));
    Odrv4 I__4690 (
            .O(N__23913),
            .I(\tok.n46 ));
    Odrv4 I__4689 (
            .O(N__23906),
            .I(\tok.n46 ));
    Odrv12 I__4688 (
            .O(N__23903),
            .I(\tok.n46 ));
    InMux I__4687 (
            .O(N__23890),
            .I(N__23887));
    LocalMux I__4686 (
            .O(N__23887),
            .I(N__23884));
    Odrv4 I__4685 (
            .O(N__23884),
            .I(\tok.n215_adj_887 ));
    CascadeMux I__4684 (
            .O(N__23881),
            .I(\tok.n207_adj_811_cascade_ ));
    InMux I__4683 (
            .O(N__23878),
            .I(N__23875));
    LocalMux I__4682 (
            .O(N__23875),
            .I(\tok.n6481 ));
    CascadeMux I__4681 (
            .O(N__23872),
            .I(N__23869));
    InMux I__4680 (
            .O(N__23869),
            .I(N__23866));
    LocalMux I__4679 (
            .O(N__23866),
            .I(\tok.n6484 ));
    InMux I__4678 (
            .O(N__23863),
            .I(N__23860));
    LocalMux I__4677 (
            .O(N__23860),
            .I(\tok.n213_adj_810 ));
    CascadeMux I__4676 (
            .O(N__23857),
            .I(N__23853));
    InMux I__4675 (
            .O(N__23856),
            .I(N__23848));
    InMux I__4674 (
            .O(N__23853),
            .I(N__23845));
    CascadeMux I__4673 (
            .O(N__23852),
            .I(N__23840));
    InMux I__4672 (
            .O(N__23851),
            .I(N__23836));
    LocalMux I__4671 (
            .O(N__23848),
            .I(N__23831));
    LocalMux I__4670 (
            .O(N__23845),
            .I(N__23831));
    CascadeMux I__4669 (
            .O(N__23844),
            .I(N__23828));
    CascadeMux I__4668 (
            .O(N__23843),
            .I(N__23825));
    InMux I__4667 (
            .O(N__23840),
            .I(N__23822));
    CascadeMux I__4666 (
            .O(N__23839),
            .I(N__23819));
    LocalMux I__4665 (
            .O(N__23836),
            .I(N__23816));
    Span4Mux_v I__4664 (
            .O(N__23831),
            .I(N__23813));
    InMux I__4663 (
            .O(N__23828),
            .I(N__23810));
    InMux I__4662 (
            .O(N__23825),
            .I(N__23807));
    LocalMux I__4661 (
            .O(N__23822),
            .I(N__23804));
    InMux I__4660 (
            .O(N__23819),
            .I(N__23801));
    Span4Mux_s3_v I__4659 (
            .O(N__23816),
            .I(N__23797));
    Span4Mux_h I__4658 (
            .O(N__23813),
            .I(N__23790));
    LocalMux I__4657 (
            .O(N__23810),
            .I(N__23790));
    LocalMux I__4656 (
            .O(N__23807),
            .I(N__23790));
    Span4Mux_v I__4655 (
            .O(N__23804),
            .I(N__23785));
    LocalMux I__4654 (
            .O(N__23801),
            .I(N__23785));
    InMux I__4653 (
            .O(N__23800),
            .I(N__23782));
    Span4Mux_h I__4652 (
            .O(N__23797),
            .I(N__23777));
    Span4Mux_h I__4651 (
            .O(N__23790),
            .I(N__23777));
    Span4Mux_h I__4650 (
            .O(N__23785),
            .I(N__23774));
    LocalMux I__4649 (
            .O(N__23782),
            .I(\tok.S_4 ));
    Odrv4 I__4648 (
            .O(N__23777),
            .I(\tok.S_4 ));
    Odrv4 I__4647 (
            .O(N__23774),
            .I(\tok.S_4 ));
    CascadeMux I__4646 (
            .O(N__23767),
            .I(\tok.n207_cascade_ ));
    InMux I__4645 (
            .O(N__23764),
            .I(N__23761));
    LocalMux I__4644 (
            .O(N__23761),
            .I(N__23758));
    Odrv4 I__4643 (
            .O(N__23758),
            .I(\tok.n210 ));
    CascadeMux I__4642 (
            .O(N__23755),
            .I(\tok.n6572_cascade_ ));
    InMux I__4641 (
            .O(N__23752),
            .I(N__23749));
    LocalMux I__4640 (
            .O(N__23749),
            .I(\tok.n174_adj_768 ));
    CascadeMux I__4639 (
            .O(N__23746),
            .I(N__23743));
    InMux I__4638 (
            .O(N__23743),
            .I(N__23738));
    InMux I__4637 (
            .O(N__23742),
            .I(N__23733));
    InMux I__4636 (
            .O(N__23741),
            .I(N__23733));
    LocalMux I__4635 (
            .O(N__23738),
            .I(N__23721));
    LocalMux I__4634 (
            .O(N__23733),
            .I(N__23721));
    InMux I__4633 (
            .O(N__23732),
            .I(N__23716));
    InMux I__4632 (
            .O(N__23731),
            .I(N__23711));
    InMux I__4631 (
            .O(N__23730),
            .I(N__23711));
    InMux I__4630 (
            .O(N__23729),
            .I(N__23706));
    InMux I__4629 (
            .O(N__23728),
            .I(N__23706));
    InMux I__4628 (
            .O(N__23727),
            .I(N__23701));
    InMux I__4627 (
            .O(N__23726),
            .I(N__23701));
    Span4Mux_h I__4626 (
            .O(N__23721),
            .I(N__23698));
    InMux I__4625 (
            .O(N__23720),
            .I(N__23693));
    InMux I__4624 (
            .O(N__23719),
            .I(N__23693));
    LocalMux I__4623 (
            .O(N__23716),
            .I(N__23690));
    LocalMux I__4622 (
            .O(N__23711),
            .I(\tok.n31 ));
    LocalMux I__4621 (
            .O(N__23706),
            .I(\tok.n31 ));
    LocalMux I__4620 (
            .O(N__23701),
            .I(\tok.n31 ));
    Odrv4 I__4619 (
            .O(N__23698),
            .I(\tok.n31 ));
    LocalMux I__4618 (
            .O(N__23693),
            .I(\tok.n31 ));
    Odrv12 I__4617 (
            .O(N__23690),
            .I(\tok.n31 ));
    CascadeMux I__4616 (
            .O(N__23677),
            .I(N__23672));
    InMux I__4615 (
            .O(N__23676),
            .I(N__23669));
    InMux I__4614 (
            .O(N__23675),
            .I(N__23666));
    InMux I__4613 (
            .O(N__23672),
            .I(N__23663));
    LocalMux I__4612 (
            .O(N__23669),
            .I(\tok.n26_adj_763 ));
    LocalMux I__4611 (
            .O(N__23666),
            .I(\tok.n26_adj_763 ));
    LocalMux I__4610 (
            .O(N__23663),
            .I(\tok.n26_adj_763 ));
    CascadeMux I__4609 (
            .O(N__23656),
            .I(\tok.n26_adj_763_cascade_ ));
    InMux I__4608 (
            .O(N__23653),
            .I(N__23650));
    LocalMux I__4607 (
            .O(N__23650),
            .I(N__23647));
    Span4Mux_v I__4606 (
            .O(N__23647),
            .I(N__23644));
    Sp12to4 I__4605 (
            .O(N__23644),
            .I(N__23641));
    Odrv12 I__4604 (
            .O(N__23641),
            .I(\tok.n6466 ));
    InMux I__4603 (
            .O(N__23638),
            .I(N__23635));
    LocalMux I__4602 (
            .O(N__23635),
            .I(N__23632));
    Odrv12 I__4601 (
            .O(N__23632),
            .I(\tok.n6467 ));
    CascadeMux I__4600 (
            .O(N__23629),
            .I(N__23626));
    InMux I__4599 (
            .O(N__23626),
            .I(N__23623));
    LocalMux I__4598 (
            .O(N__23623),
            .I(N__23620));
    Odrv4 I__4597 (
            .O(N__23620),
            .I(\tok.n6486 ));
    CascadeMux I__4596 (
            .O(N__23617),
            .I(N__23613));
    InMux I__4595 (
            .O(N__23616),
            .I(N__23609));
    InMux I__4594 (
            .O(N__23613),
            .I(N__23606));
    InMux I__4593 (
            .O(N__23612),
            .I(N__23603));
    LocalMux I__4592 (
            .O(N__23609),
            .I(N__23600));
    LocalMux I__4591 (
            .O(N__23606),
            .I(N__23597));
    LocalMux I__4590 (
            .O(N__23603),
            .I(N__23594));
    Span4Mux_h I__4589 (
            .O(N__23600),
            .I(N__23591));
    Span4Mux_v I__4588 (
            .O(N__23597),
            .I(N__23586));
    Span4Mux_v I__4587 (
            .O(N__23594),
            .I(N__23586));
    Odrv4 I__4586 (
            .O(N__23591),
            .I(\tok.n833 ));
    Odrv4 I__4585 (
            .O(N__23586),
            .I(\tok.n833 ));
    InMux I__4584 (
            .O(N__23581),
            .I(N__23578));
    LocalMux I__4583 (
            .O(N__23578),
            .I(N__23575));
    Span4Mux_h I__4582 (
            .O(N__23575),
            .I(N__23572));
    Odrv4 I__4581 (
            .O(N__23572),
            .I(\tok.n6490 ));
    CascadeMux I__4580 (
            .O(N__23569),
            .I(N__23566));
    InMux I__4579 (
            .O(N__23566),
            .I(N__23563));
    LocalMux I__4578 (
            .O(N__23563),
            .I(N__23560));
    Span4Mux_h I__4577 (
            .O(N__23560),
            .I(N__23557));
    Odrv4 I__4576 (
            .O(N__23557),
            .I(\tok.n6491 ));
    CascadeMux I__4575 (
            .O(N__23554),
            .I(N__23550));
    InMux I__4574 (
            .O(N__23553),
            .I(N__23543));
    InMux I__4573 (
            .O(N__23550),
            .I(N__23540));
    InMux I__4572 (
            .O(N__23549),
            .I(N__23537));
    InMux I__4571 (
            .O(N__23548),
            .I(N__23534));
    CascadeMux I__4570 (
            .O(N__23547),
            .I(N__23531));
    CascadeMux I__4569 (
            .O(N__23546),
            .I(N__23528));
    LocalMux I__4568 (
            .O(N__23543),
            .I(N__23525));
    LocalMux I__4567 (
            .O(N__23540),
            .I(N__23520));
    LocalMux I__4566 (
            .O(N__23537),
            .I(N__23520));
    LocalMux I__4565 (
            .O(N__23534),
            .I(N__23517));
    InMux I__4564 (
            .O(N__23531),
            .I(N__23514));
    InMux I__4563 (
            .O(N__23528),
            .I(N__23511));
    Span4Mux_v I__4562 (
            .O(N__23525),
            .I(N__23506));
    Span4Mux_v I__4561 (
            .O(N__23520),
            .I(N__23506));
    Span4Mux_v I__4560 (
            .O(N__23517),
            .I(N__23503));
    LocalMux I__4559 (
            .O(N__23514),
            .I(N__23500));
    LocalMux I__4558 (
            .O(N__23511),
            .I(N__23497));
    Span4Mux_h I__4557 (
            .O(N__23506),
            .I(N__23486));
    Span4Mux_h I__4556 (
            .O(N__23503),
            .I(N__23486));
    Span4Mux_v I__4555 (
            .O(N__23500),
            .I(N__23486));
    Span4Mux_v I__4554 (
            .O(N__23497),
            .I(N__23486));
    InMux I__4553 (
            .O(N__23496),
            .I(N__23483));
    InMux I__4552 (
            .O(N__23495),
            .I(N__23480));
    Span4Mux_v I__4551 (
            .O(N__23486),
            .I(N__23477));
    LocalMux I__4550 (
            .O(N__23483),
            .I(S_1));
    LocalMux I__4549 (
            .O(N__23480),
            .I(S_1));
    Odrv4 I__4548 (
            .O(N__23477),
            .I(S_1));
    InMux I__4547 (
            .O(N__23470),
            .I(N__23467));
    LocalMux I__4546 (
            .O(N__23467),
            .I(N__23464));
    Span4Mux_h I__4545 (
            .O(N__23464),
            .I(N__23461));
    Odrv4 I__4544 (
            .O(N__23461),
            .I(\tok.n208 ));
    CascadeMux I__4543 (
            .O(N__23458),
            .I(N__23455));
    InMux I__4542 (
            .O(N__23455),
            .I(N__23452));
    LocalMux I__4541 (
            .O(N__23452),
            .I(N__23449));
    Span4Mux_h I__4540 (
            .O(N__23449),
            .I(N__23446));
    Span4Mux_s3_h I__4539 (
            .O(N__23446),
            .I(N__23443));
    Odrv4 I__4538 (
            .O(N__23443),
            .I(\tok.n6589 ));
    InMux I__4537 (
            .O(N__23440),
            .I(N__23437));
    LocalMux I__4536 (
            .O(N__23437),
            .I(N__23434));
    Span12Mux_s6_h I__4535 (
            .O(N__23434),
            .I(N__23431));
    Odrv12 I__4534 (
            .O(N__23431),
            .I(\tok.n239_adj_727 ));
    CascadeMux I__4533 (
            .O(N__23428),
            .I(\tok.n6_adj_728_cascade_ ));
    CascadeMux I__4532 (
            .O(N__23425),
            .I(\tok.n200_adj_732_cascade_ ));
    InMux I__4531 (
            .O(N__23422),
            .I(N__23419));
    LocalMux I__4530 (
            .O(N__23419),
            .I(N__23416));
    Odrv12 I__4529 (
            .O(N__23416),
            .I(\tok.n203_adj_731 ));
    InMux I__4528 (
            .O(N__23413),
            .I(N__23410));
    LocalMux I__4527 (
            .O(N__23410),
            .I(N__23407));
    Span4Mux_h I__4526 (
            .O(N__23407),
            .I(N__23404));
    Odrv4 I__4525 (
            .O(N__23404),
            .I(\tok.n6_adj_733 ));
    InMux I__4524 (
            .O(N__23401),
            .I(N__23397));
    InMux I__4523 (
            .O(N__23400),
            .I(N__23394));
    LocalMux I__4522 (
            .O(N__23397),
            .I(N__23389));
    LocalMux I__4521 (
            .O(N__23394),
            .I(N__23389));
    Span4Mux_v I__4520 (
            .O(N__23389),
            .I(N__23386));
    Span4Mux_v I__4519 (
            .O(N__23386),
            .I(N__23383));
    Odrv4 I__4518 (
            .O(N__23383),
            .I(\tok.n206_adj_794 ));
    CascadeMux I__4517 (
            .O(N__23380),
            .I(\tok.n244_cascade_ ));
    CascadeMux I__4516 (
            .O(N__23377),
            .I(\tok.n4_adj_720_cascade_ ));
    InMux I__4515 (
            .O(N__23374),
            .I(N__23371));
    LocalMux I__4514 (
            .O(N__23371),
            .I(N__23368));
    Odrv12 I__4513 (
            .O(N__23368),
            .I(\tok.n145 ));
    InMux I__4512 (
            .O(N__23365),
            .I(N__23362));
    LocalMux I__4511 (
            .O(N__23362),
            .I(\tok.n251 ));
    InMux I__4510 (
            .O(N__23359),
            .I(N__23356));
    LocalMux I__4509 (
            .O(N__23356),
            .I(N__23352));
    InMux I__4508 (
            .O(N__23355),
            .I(N__23349));
    Span4Mux_h I__4507 (
            .O(N__23352),
            .I(N__23346));
    LocalMux I__4506 (
            .O(N__23349),
            .I(N__23343));
    Span4Mux_v I__4505 (
            .O(N__23346),
            .I(N__23340));
    Span4Mux_v I__4504 (
            .O(N__23343),
            .I(N__23337));
    Odrv4 I__4503 (
            .O(N__23340),
            .I(\tok.n2557 ));
    Odrv4 I__4502 (
            .O(N__23337),
            .I(\tok.n2557 ));
    CascadeMux I__4501 (
            .O(N__23332),
            .I(\tok.n4_adj_714_cascade_ ));
    InMux I__4500 (
            .O(N__23329),
            .I(N__23326));
    LocalMux I__4499 (
            .O(N__23326),
            .I(\tok.n218 ));
    InMux I__4498 (
            .O(N__23323),
            .I(N__23320));
    LocalMux I__4497 (
            .O(N__23320),
            .I(\tok.n39 ));
    CascadeMux I__4496 (
            .O(N__23317),
            .I(\tok.n6269_cascade_ ));
    CascadeMux I__4495 (
            .O(N__23314),
            .I(\tok.n197_adj_729_cascade_ ));
    InMux I__4494 (
            .O(N__23311),
            .I(N__23308));
    LocalMux I__4493 (
            .O(N__23308),
            .I(N__23305));
    Odrv4 I__4492 (
            .O(N__23305),
            .I(\tok.n7458 ));
    InMux I__4491 (
            .O(N__23302),
            .I(N__23299));
    LocalMux I__4490 (
            .O(N__23299),
            .I(\tok.n2544 ));
    CascadeMux I__4489 (
            .O(N__23296),
            .I(N__23292));
    InMux I__4488 (
            .O(N__23295),
            .I(N__23289));
    InMux I__4487 (
            .O(N__23292),
            .I(N__23286));
    LocalMux I__4486 (
            .O(N__23289),
            .I(N__23283));
    LocalMux I__4485 (
            .O(N__23286),
            .I(N__23280));
    Span4Mux_v I__4484 (
            .O(N__23283),
            .I(N__23277));
    Sp12to4 I__4483 (
            .O(N__23280),
            .I(N__23274));
    Span4Mux_h I__4482 (
            .O(N__23277),
            .I(N__23271));
    Span12Mux_s10_h I__4481 (
            .O(N__23274),
            .I(N__23268));
    Odrv4 I__4480 (
            .O(N__23271),
            .I(\tok.table_rd_1 ));
    Odrv12 I__4479 (
            .O(N__23268),
            .I(\tok.table_rd_1 ));
    CascadeMux I__4478 (
            .O(N__23263),
            .I(\tok.n7475_cascade_ ));
    InMux I__4477 (
            .O(N__23260),
            .I(N__23256));
    InMux I__4476 (
            .O(N__23259),
            .I(N__23253));
    LocalMux I__4475 (
            .O(N__23256),
            .I(N__23248));
    LocalMux I__4474 (
            .O(N__23253),
            .I(N__23248));
    Span4Mux_h I__4473 (
            .O(N__23248),
            .I(N__23245));
    Span4Mux_h I__4472 (
            .O(N__23245),
            .I(N__23242));
    Odrv4 I__4471 (
            .O(N__23242),
            .I(\tok.n237 ));
    CascadeMux I__4470 (
            .O(N__23239),
            .I(N__23236));
    InMux I__4469 (
            .O(N__23236),
            .I(N__23233));
    LocalMux I__4468 (
            .O(N__23233),
            .I(N__23230));
    Odrv4 I__4467 (
            .O(N__23230),
            .I(\tok.n180 ));
    CascadeMux I__4466 (
            .O(N__23227),
            .I(N__23224));
    InMux I__4465 (
            .O(N__23224),
            .I(N__23221));
    LocalMux I__4464 (
            .O(N__23221),
            .I(\tok.n6628 ));
    InMux I__4463 (
            .O(N__23218),
            .I(N__23212));
    InMux I__4462 (
            .O(N__23217),
            .I(N__23206));
    InMux I__4461 (
            .O(N__23216),
            .I(N__23203));
    CascadeMux I__4460 (
            .O(N__23215),
            .I(N__23200));
    LocalMux I__4459 (
            .O(N__23212),
            .I(N__23197));
    InMux I__4458 (
            .O(N__23211),
            .I(N__23194));
    InMux I__4457 (
            .O(N__23210),
            .I(N__23191));
    InMux I__4456 (
            .O(N__23209),
            .I(N__23188));
    LocalMux I__4455 (
            .O(N__23206),
            .I(N__23185));
    LocalMux I__4454 (
            .O(N__23203),
            .I(N__23182));
    InMux I__4453 (
            .O(N__23200),
            .I(N__23179));
    Span4Mux_v I__4452 (
            .O(N__23197),
            .I(N__23173));
    LocalMux I__4451 (
            .O(N__23194),
            .I(N__23173));
    LocalMux I__4450 (
            .O(N__23191),
            .I(N__23170));
    LocalMux I__4449 (
            .O(N__23188),
            .I(N__23161));
    Span4Mux_h I__4448 (
            .O(N__23185),
            .I(N__23161));
    Span4Mux_v I__4447 (
            .O(N__23182),
            .I(N__23161));
    LocalMux I__4446 (
            .O(N__23179),
            .I(N__23161));
    InMux I__4445 (
            .O(N__23178),
            .I(N__23158));
    Span4Mux_v I__4444 (
            .O(N__23173),
            .I(N__23155));
    Span4Mux_v I__4443 (
            .O(N__23170),
            .I(N__23150));
    Span4Mux_h I__4442 (
            .O(N__23161),
            .I(N__23150));
    LocalMux I__4441 (
            .O(N__23158),
            .I(\tok.S_3 ));
    Odrv4 I__4440 (
            .O(N__23155),
            .I(\tok.S_3 ));
    Odrv4 I__4439 (
            .O(N__23150),
            .I(\tok.S_3 ));
    CascadeMux I__4438 (
            .O(N__23143),
            .I(N__23140));
    InMux I__4437 (
            .O(N__23140),
            .I(N__23137));
    LocalMux I__4436 (
            .O(N__23137),
            .I(N__23134));
    Odrv4 I__4435 (
            .O(N__23134),
            .I(\tok.n241 ));
    InMux I__4434 (
            .O(N__23131),
            .I(N__23128));
    LocalMux I__4433 (
            .O(N__23128),
            .I(N__23125));
    Odrv4 I__4432 (
            .O(N__23125),
            .I(\tok.n6637 ));
    CascadeMux I__4431 (
            .O(N__23122),
            .I(\tok.n284_cascade_ ));
    InMux I__4430 (
            .O(N__23119),
            .I(N__23116));
    LocalMux I__4429 (
            .O(N__23116),
            .I(\tok.n17 ));
    CascadeMux I__4428 (
            .O(N__23113),
            .I(N__23110));
    InMux I__4427 (
            .O(N__23110),
            .I(N__23107));
    LocalMux I__4426 (
            .O(N__23107),
            .I(N__23103));
    InMux I__4425 (
            .O(N__23106),
            .I(N__23100));
    Span12Mux_s9_h I__4424 (
            .O(N__23103),
            .I(N__23097));
    LocalMux I__4423 (
            .O(N__23100),
            .I(\tok.n5_adj_821 ));
    Odrv12 I__4422 (
            .O(N__23097),
            .I(\tok.n5_adj_821 ));
    InMux I__4421 (
            .O(N__23092),
            .I(N__23089));
    LocalMux I__4420 (
            .O(N__23089),
            .I(\tok.n2679 ));
    CascadeMux I__4419 (
            .O(N__23086),
            .I(\tok.n17_cascade_ ));
    CascadeMux I__4418 (
            .O(N__23083),
            .I(N__23080));
    InMux I__4417 (
            .O(N__23080),
            .I(N__23077));
    LocalMux I__4416 (
            .O(N__23077),
            .I(\tok.n864 ));
    InMux I__4415 (
            .O(N__23074),
            .I(N__23071));
    LocalMux I__4414 (
            .O(N__23071),
            .I(N__23068));
    Odrv4 I__4413 (
            .O(N__23068),
            .I(\tok.n186 ));
    CascadeMux I__4412 (
            .O(N__23065),
            .I(\tok.n6562_cascade_ ));
    CascadeMux I__4411 (
            .O(N__23062),
            .I(N__23059));
    InMux I__4410 (
            .O(N__23059),
            .I(N__23056));
    LocalMux I__4409 (
            .O(N__23056),
            .I(N__23053));
    Span4Mux_v I__4408 (
            .O(N__23053),
            .I(N__23050));
    Odrv4 I__4407 (
            .O(N__23050),
            .I(\tok.n338 ));
    InMux I__4406 (
            .O(N__23047),
            .I(N__23044));
    LocalMux I__4405 (
            .O(N__23044),
            .I(\tok.n162 ));
    InMux I__4404 (
            .O(N__23041),
            .I(N__23038));
    LocalMux I__4403 (
            .O(N__23038),
            .I(\tok.n179_adj_730 ));
    InMux I__4402 (
            .O(N__23035),
            .I(N__23032));
    LocalMux I__4401 (
            .O(N__23032),
            .I(N__23029));
    Span4Mux_v I__4400 (
            .O(N__23029),
            .I(N__23026));
    Odrv4 I__4399 (
            .O(N__23026),
            .I(\tok.n4926 ));
    CascadeMux I__4398 (
            .O(N__23023),
            .I(\tok.n2692_cascade_ ));
    InMux I__4397 (
            .O(N__23020),
            .I(N__23017));
    LocalMux I__4396 (
            .O(N__23017),
            .I(N__23014));
    Span4Mux_h I__4395 (
            .O(N__23014),
            .I(N__23011));
    Odrv4 I__4394 (
            .O(N__23011),
            .I(\tok.n217 ));
    InMux I__4393 (
            .O(N__23008),
            .I(N__23005));
    LocalMux I__4392 (
            .O(N__23005),
            .I(\tok.n7154 ));
    InMux I__4391 (
            .O(N__23002),
            .I(N__22999));
    LocalMux I__4390 (
            .O(N__22999),
            .I(\tok.n6_adj_701 ));
    InMux I__4389 (
            .O(N__22996),
            .I(N__22993));
    LocalMux I__4388 (
            .O(N__22993),
            .I(\tok.n2700 ));
    InMux I__4387 (
            .O(N__22990),
            .I(N__22987));
    LocalMux I__4386 (
            .O(N__22987),
            .I(\tok.n236_adj_737 ));
    InMux I__4385 (
            .O(N__22984),
            .I(N__22981));
    LocalMux I__4384 (
            .O(N__22981),
            .I(N__22978));
    Span4Mux_h I__4383 (
            .O(N__22978),
            .I(N__22975));
    Odrv4 I__4382 (
            .O(N__22975),
            .I(\tok.n239_adj_738 ));
    InMux I__4381 (
            .O(N__22972),
            .I(N__22966));
    InMux I__4380 (
            .O(N__22971),
            .I(N__22966));
    LocalMux I__4379 (
            .O(N__22966),
            .I(\tok.C_stk.tail_19 ));
    InMux I__4378 (
            .O(N__22963),
            .I(N__22957));
    InMux I__4377 (
            .O(N__22962),
            .I(N__22957));
    LocalMux I__4376 (
            .O(N__22957),
            .I(\tok.C_stk.tail_27 ));
    InMux I__4375 (
            .O(N__22954),
            .I(N__22948));
    InMux I__4374 (
            .O(N__22953),
            .I(N__22948));
    LocalMux I__4373 (
            .O(N__22948),
            .I(\tok.C_stk.tail_35 ));
    InMux I__4372 (
            .O(N__22945),
            .I(N__22940));
    InMux I__4371 (
            .O(N__22944),
            .I(N__22936));
    InMux I__4370 (
            .O(N__22943),
            .I(N__22933));
    LocalMux I__4369 (
            .O(N__22940),
            .I(N__22928));
    InMux I__4368 (
            .O(N__22939),
            .I(N__22925));
    LocalMux I__4367 (
            .O(N__22936),
            .I(N__22922));
    LocalMux I__4366 (
            .O(N__22933),
            .I(N__22919));
    InMux I__4365 (
            .O(N__22932),
            .I(N__22916));
    InMux I__4364 (
            .O(N__22931),
            .I(N__22911));
    Span4Mux_v I__4363 (
            .O(N__22928),
            .I(N__22906));
    LocalMux I__4362 (
            .O(N__22925),
            .I(N__22906));
    Span4Mux_v I__4361 (
            .O(N__22922),
            .I(N__22903));
    Span4Mux_v I__4360 (
            .O(N__22919),
            .I(N__22898));
    LocalMux I__4359 (
            .O(N__22916),
            .I(N__22898));
    InMux I__4358 (
            .O(N__22915),
            .I(N__22895));
    InMux I__4357 (
            .O(N__22914),
            .I(N__22892));
    LocalMux I__4356 (
            .O(N__22911),
            .I(N__22885));
    Span4Mux_h I__4355 (
            .O(N__22906),
            .I(N__22885));
    Span4Mux_s2_v I__4354 (
            .O(N__22903),
            .I(N__22885));
    Odrv4 I__4353 (
            .O(N__22898),
            .I(\tok.n4_adj_726 ));
    LocalMux I__4352 (
            .O(N__22895),
            .I(\tok.n4_adj_726 ));
    LocalMux I__4351 (
            .O(N__22892),
            .I(\tok.n4_adj_726 ));
    Odrv4 I__4350 (
            .O(N__22885),
            .I(\tok.n4_adj_726 ));
    CascadeMux I__4349 (
            .O(N__22876),
            .I(N__22871));
    InMux I__4348 (
            .O(N__22875),
            .I(N__22865));
    InMux I__4347 (
            .O(N__22874),
            .I(N__22860));
    InMux I__4346 (
            .O(N__22871),
            .I(N__22857));
    InMux I__4345 (
            .O(N__22870),
            .I(N__22854));
    InMux I__4344 (
            .O(N__22869),
            .I(N__22851));
    InMux I__4343 (
            .O(N__22868),
            .I(N__22848));
    LocalMux I__4342 (
            .O(N__22865),
            .I(N__22845));
    InMux I__4341 (
            .O(N__22864),
            .I(N__22842));
    InMux I__4340 (
            .O(N__22863),
            .I(N__22839));
    LocalMux I__4339 (
            .O(N__22860),
            .I(N__22832));
    LocalMux I__4338 (
            .O(N__22857),
            .I(N__22832));
    LocalMux I__4337 (
            .O(N__22854),
            .I(N__22832));
    LocalMux I__4336 (
            .O(N__22851),
            .I(N__22827));
    LocalMux I__4335 (
            .O(N__22848),
            .I(N__22827));
    Span4Mux_h I__4334 (
            .O(N__22845),
            .I(N__22818));
    LocalMux I__4333 (
            .O(N__22842),
            .I(N__22818));
    LocalMux I__4332 (
            .O(N__22839),
            .I(N__22818));
    Span4Mux_h I__4331 (
            .O(N__22832),
            .I(N__22818));
    Span4Mux_h I__4330 (
            .O(N__22827),
            .I(N__22815));
    Span4Mux_v I__4329 (
            .O(N__22818),
            .I(N__22812));
    Odrv4 I__4328 (
            .O(N__22815),
            .I(\tok.tc__7__N_133 ));
    Odrv4 I__4327 (
            .O(N__22812),
            .I(\tok.tc__7__N_133 ));
    InMux I__4326 (
            .O(N__22807),
            .I(N__22803));
    InMux I__4325 (
            .O(N__22806),
            .I(N__22798));
    LocalMux I__4324 (
            .O(N__22803),
            .I(N__22795));
    InMux I__4323 (
            .O(N__22802),
            .I(N__22792));
    InMux I__4322 (
            .O(N__22801),
            .I(N__22787));
    LocalMux I__4321 (
            .O(N__22798),
            .I(N__22780));
    Span4Mux_s3_v I__4320 (
            .O(N__22795),
            .I(N__22780));
    LocalMux I__4319 (
            .O(N__22792),
            .I(N__22780));
    InMux I__4318 (
            .O(N__22791),
            .I(N__22776));
    InMux I__4317 (
            .O(N__22790),
            .I(N__22772));
    LocalMux I__4316 (
            .O(N__22787),
            .I(N__22769));
    Span4Mux_h I__4315 (
            .O(N__22780),
            .I(N__22766));
    InMux I__4314 (
            .O(N__22779),
            .I(N__22763));
    LocalMux I__4313 (
            .O(N__22776),
            .I(N__22760));
    InMux I__4312 (
            .O(N__22775),
            .I(N__22757));
    LocalMux I__4311 (
            .O(N__22772),
            .I(\tok.n2573 ));
    Odrv12 I__4310 (
            .O(N__22769),
            .I(\tok.n2573 ));
    Odrv4 I__4309 (
            .O(N__22766),
            .I(\tok.n2573 ));
    LocalMux I__4308 (
            .O(N__22763),
            .I(\tok.n2573 ));
    Odrv4 I__4307 (
            .O(N__22760),
            .I(\tok.n2573 ));
    LocalMux I__4306 (
            .O(N__22757),
            .I(\tok.n2573 ));
    CascadeMux I__4305 (
            .O(N__22744),
            .I(\tok.n6291_cascade_ ));
    CascadeMux I__4304 (
            .O(N__22741),
            .I(\tok.n80_adj_735_cascade_ ));
    CascadeMux I__4303 (
            .O(N__22738),
            .I(\tok.n83_adj_725_cascade_ ));
    InMux I__4302 (
            .O(N__22735),
            .I(N__22732));
    LocalMux I__4301 (
            .O(N__22732),
            .I(\tok.n6287 ));
    InMux I__4300 (
            .O(N__22729),
            .I(N__22726));
    LocalMux I__4299 (
            .O(N__22726),
            .I(\tok.n89_adj_736 ));
    CascadeMux I__4298 (
            .O(N__22723),
            .I(N__22720));
    InMux I__4297 (
            .O(N__22720),
            .I(N__22716));
    InMux I__4296 (
            .O(N__22719),
            .I(N__22713));
    LocalMux I__4295 (
            .O(N__22716),
            .I(N__22710));
    LocalMux I__4294 (
            .O(N__22713),
            .I(N__22707));
    Span4Mux_h I__4293 (
            .O(N__22710),
            .I(N__22702));
    Span4Mux_h I__4292 (
            .O(N__22707),
            .I(N__22702));
    Odrv4 I__4291 (
            .O(N__22702),
            .I(n92));
    InMux I__4290 (
            .O(N__22699),
            .I(N__22693));
    InMux I__4289 (
            .O(N__22698),
            .I(N__22693));
    LocalMux I__4288 (
            .O(N__22693),
            .I(\tok.tail_10 ));
    CascadeMux I__4287 (
            .O(N__22690),
            .I(N__22687));
    InMux I__4286 (
            .O(N__22687),
            .I(N__22681));
    InMux I__4285 (
            .O(N__22686),
            .I(N__22681));
    LocalMux I__4284 (
            .O(N__22681),
            .I(\tok.C_stk.tail_18 ));
    InMux I__4283 (
            .O(N__22678),
            .I(N__22672));
    InMux I__4282 (
            .O(N__22677),
            .I(N__22672));
    LocalMux I__4281 (
            .O(N__22672),
            .I(\tok.tail_26 ));
    InMux I__4280 (
            .O(N__22669),
            .I(N__22663));
    InMux I__4279 (
            .O(N__22668),
            .I(N__22663));
    LocalMux I__4278 (
            .O(N__22663),
            .I(\tok.C_stk.tail_34 ));
    CascadeMux I__4277 (
            .O(N__22660),
            .I(N__22656));
    InMux I__4276 (
            .O(N__22659),
            .I(N__22650));
    InMux I__4275 (
            .O(N__22656),
            .I(N__22650));
    InMux I__4274 (
            .O(N__22655),
            .I(N__22647));
    LocalMux I__4273 (
            .O(N__22650),
            .I(N__22643));
    LocalMux I__4272 (
            .O(N__22647),
            .I(N__22640));
    InMux I__4271 (
            .O(N__22646),
            .I(N__22637));
    Span4Mux_v I__4270 (
            .O(N__22643),
            .I(N__22634));
    Span4Mux_v I__4269 (
            .O(N__22640),
            .I(N__22627));
    LocalMux I__4268 (
            .O(N__22637),
            .I(N__22627));
    Span4Mux_s1_v I__4267 (
            .O(N__22634),
            .I(N__22627));
    Odrv4 I__4266 (
            .O(N__22627),
            .I(\tok.tc_plus_1_3 ));
    CascadeMux I__4265 (
            .O(N__22624),
            .I(\tok.C_stk.n6242_cascade_ ));
    InMux I__4264 (
            .O(N__22621),
            .I(N__22617));
    InMux I__4263 (
            .O(N__22620),
            .I(N__22614));
    LocalMux I__4262 (
            .O(N__22617),
            .I(N__22611));
    LocalMux I__4261 (
            .O(N__22614),
            .I(N__22607));
    Span4Mux_h I__4260 (
            .O(N__22611),
            .I(N__22603));
    InMux I__4259 (
            .O(N__22610),
            .I(N__22600));
    Span4Mux_v I__4258 (
            .O(N__22607),
            .I(N__22597));
    InMux I__4257 (
            .O(N__22606),
            .I(N__22594));
    Odrv4 I__4256 (
            .O(N__22603),
            .I(tc_3));
    LocalMux I__4255 (
            .O(N__22600),
            .I(tc_3));
    Odrv4 I__4254 (
            .O(N__22597),
            .I(tc_3));
    LocalMux I__4253 (
            .O(N__22594),
            .I(tc_3));
    InMux I__4252 (
            .O(N__22585),
            .I(N__22579));
    InMux I__4251 (
            .O(N__22584),
            .I(N__22572));
    InMux I__4250 (
            .O(N__22583),
            .I(N__22572));
    InMux I__4249 (
            .O(N__22582),
            .I(N__22572));
    LocalMux I__4248 (
            .O(N__22579),
            .I(\tok.c_stk_r_3 ));
    LocalMux I__4247 (
            .O(N__22572),
            .I(\tok.c_stk_r_3 ));
    InMux I__4246 (
            .O(N__22567),
            .I(N__22561));
    InMux I__4245 (
            .O(N__22566),
            .I(N__22561));
    LocalMux I__4244 (
            .O(N__22561),
            .I(\tok.C_stk.tail_3 ));
    InMux I__4243 (
            .O(N__22558),
            .I(N__22552));
    InMux I__4242 (
            .O(N__22557),
            .I(N__22552));
    LocalMux I__4241 (
            .O(N__22552),
            .I(\tok.C_stk.tail_11 ));
    InMux I__4240 (
            .O(N__22549),
            .I(N__22543));
    InMux I__4239 (
            .O(N__22548),
            .I(N__22543));
    LocalMux I__4238 (
            .O(N__22543),
            .I(\tok.C_stk.tail_5 ));
    InMux I__4237 (
            .O(N__22540),
            .I(N__22534));
    InMux I__4236 (
            .O(N__22539),
            .I(N__22534));
    LocalMux I__4235 (
            .O(N__22534),
            .I(\tok.tail_13 ));
    CascadeMux I__4234 (
            .O(N__22531),
            .I(N__22528));
    InMux I__4233 (
            .O(N__22528),
            .I(N__22522));
    InMux I__4232 (
            .O(N__22527),
            .I(N__22522));
    LocalMux I__4231 (
            .O(N__22522),
            .I(\tok.C_stk.tail_21 ));
    InMux I__4230 (
            .O(N__22519),
            .I(N__22513));
    InMux I__4229 (
            .O(N__22518),
            .I(N__22513));
    LocalMux I__4228 (
            .O(N__22513),
            .I(\tok.tail_29 ));
    InMux I__4227 (
            .O(N__22510),
            .I(N__22504));
    InMux I__4226 (
            .O(N__22509),
            .I(N__22504));
    LocalMux I__4225 (
            .O(N__22504),
            .I(\tok.C_stk.tail_37 ));
    CascadeMux I__4224 (
            .O(N__22501),
            .I(N__22498));
    InMux I__4223 (
            .O(N__22498),
            .I(N__22491));
    InMux I__4222 (
            .O(N__22497),
            .I(N__22491));
    InMux I__4221 (
            .O(N__22496),
            .I(N__22488));
    LocalMux I__4220 (
            .O(N__22491),
            .I(N__22484));
    LocalMux I__4219 (
            .O(N__22488),
            .I(N__22481));
    InMux I__4218 (
            .O(N__22487),
            .I(N__22478));
    Span4Mux_h I__4217 (
            .O(N__22484),
            .I(N__22475));
    Odrv4 I__4216 (
            .O(N__22481),
            .I(\tok.tc_plus_1_2 ));
    LocalMux I__4215 (
            .O(N__22478),
            .I(\tok.tc_plus_1_2 ));
    Odrv4 I__4214 (
            .O(N__22475),
            .I(\tok.tc_plus_1_2 ));
    CascadeMux I__4213 (
            .O(N__22468),
            .I(\tok.C_stk.n6245_cascade_ ));
    InMux I__4212 (
            .O(N__22465),
            .I(N__22461));
    InMux I__4211 (
            .O(N__22464),
            .I(N__22457));
    LocalMux I__4210 (
            .O(N__22461),
            .I(N__22453));
    InMux I__4209 (
            .O(N__22460),
            .I(N__22450));
    LocalMux I__4208 (
            .O(N__22457),
            .I(N__22447));
    InMux I__4207 (
            .O(N__22456),
            .I(N__22444));
    Odrv4 I__4206 (
            .O(N__22453),
            .I(tc_2));
    LocalMux I__4205 (
            .O(N__22450),
            .I(tc_2));
    Odrv12 I__4204 (
            .O(N__22447),
            .I(tc_2));
    LocalMux I__4203 (
            .O(N__22444),
            .I(tc_2));
    CascadeMux I__4202 (
            .O(N__22435),
            .I(N__22429));
    InMux I__4201 (
            .O(N__22434),
            .I(N__22426));
    InMux I__4200 (
            .O(N__22433),
            .I(N__22421));
    InMux I__4199 (
            .O(N__22432),
            .I(N__22421));
    InMux I__4198 (
            .O(N__22429),
            .I(N__22418));
    LocalMux I__4197 (
            .O(N__22426),
            .I(\tok.c_stk_r_2 ));
    LocalMux I__4196 (
            .O(N__22421),
            .I(\tok.c_stk_r_2 ));
    LocalMux I__4195 (
            .O(N__22418),
            .I(\tok.c_stk_r_2 ));
    InMux I__4194 (
            .O(N__22411),
            .I(N__22405));
    InMux I__4193 (
            .O(N__22410),
            .I(N__22405));
    LocalMux I__4192 (
            .O(N__22405),
            .I(\tok.C_stk.tail_2 ));
    CascadeMux I__4191 (
            .O(N__22402),
            .I(\tok.n6404_cascade_ ));
    InMux I__4190 (
            .O(N__22399),
            .I(N__22396));
    LocalMux I__4189 (
            .O(N__22396),
            .I(\tok.n179_adj_888 ));
    CascadeMux I__4188 (
            .O(N__22393),
            .I(\tok.n6550_cascade_ ));
    InMux I__4187 (
            .O(N__22390),
            .I(N__22387));
    LocalMux I__4186 (
            .O(N__22387),
            .I(N__22384));
    Odrv4 I__4185 (
            .O(N__22384),
            .I(\tok.n6549 ));
    CascadeMux I__4184 (
            .O(N__22381),
            .I(N__22378));
    InMux I__4183 (
            .O(N__22378),
            .I(N__22375));
    LocalMux I__4182 (
            .O(N__22375),
            .I(\tok.n6419 ));
    InMux I__4181 (
            .O(N__22372),
            .I(N__22369));
    LocalMux I__4180 (
            .O(N__22369),
            .I(N__22366));
    Span4Mux_s1_v I__4179 (
            .O(N__22366),
            .I(N__22363));
    Odrv4 I__4178 (
            .O(N__22363),
            .I(\tok.n215_adj_697 ));
    CascadeMux I__4177 (
            .O(N__22360),
            .I(\tok.n6337_cascade_ ));
    CascadeMux I__4176 (
            .O(N__22357),
            .I(N__22354));
    InMux I__4175 (
            .O(N__22354),
            .I(N__22351));
    LocalMux I__4174 (
            .O(N__22351),
            .I(\tok.n6538 ));
    InMux I__4173 (
            .O(N__22348),
            .I(N__22344));
    InMux I__4172 (
            .O(N__22347),
            .I(N__22341));
    LocalMux I__4171 (
            .O(N__22344),
            .I(N__22338));
    LocalMux I__4170 (
            .O(N__22341),
            .I(N__22335));
    Span4Mux_h I__4169 (
            .O(N__22338),
            .I(N__22328));
    Span4Mux_v I__4168 (
            .O(N__22335),
            .I(N__22328));
    InMux I__4167 (
            .O(N__22334),
            .I(N__22323));
    InMux I__4166 (
            .O(N__22333),
            .I(N__22323));
    Odrv4 I__4165 (
            .O(N__22328),
            .I(\tok.tc_plus_1_5 ));
    LocalMux I__4164 (
            .O(N__22323),
            .I(\tok.tc_plus_1_5 ));
    CascadeMux I__4163 (
            .O(N__22318),
            .I(\tok.C_stk.n6236_cascade_ ));
    InMux I__4162 (
            .O(N__22315),
            .I(N__22312));
    LocalMux I__4161 (
            .O(N__22312),
            .I(N__22309));
    Span4Mux_s2_v I__4160 (
            .O(N__22309),
            .I(N__22303));
    InMux I__4159 (
            .O(N__22308),
            .I(N__22298));
    InMux I__4158 (
            .O(N__22307),
            .I(N__22298));
    InMux I__4157 (
            .O(N__22306),
            .I(N__22295));
    Odrv4 I__4156 (
            .O(N__22303),
            .I(tc_5));
    LocalMux I__4155 (
            .O(N__22298),
            .I(tc_5));
    LocalMux I__4154 (
            .O(N__22295),
            .I(tc_5));
    InMux I__4153 (
            .O(N__22288),
            .I(N__22279));
    InMux I__4152 (
            .O(N__22287),
            .I(N__22279));
    InMux I__4151 (
            .O(N__22286),
            .I(N__22279));
    LocalMux I__4150 (
            .O(N__22279),
            .I(N__22275));
    InMux I__4149 (
            .O(N__22278),
            .I(N__22272));
    Span4Mux_v I__4148 (
            .O(N__22275),
            .I(N__22269));
    LocalMux I__4147 (
            .O(N__22272),
            .I(\tok.c_stk_r_5 ));
    Odrv4 I__4146 (
            .O(N__22269),
            .I(\tok.c_stk_r_5 ));
    CascadeMux I__4145 (
            .O(N__22264),
            .I(N__22261));
    InMux I__4144 (
            .O(N__22261),
            .I(N__22258));
    LocalMux I__4143 (
            .O(N__22258),
            .I(\tok.n6320 ));
    InMux I__4142 (
            .O(N__22255),
            .I(N__22252));
    LocalMux I__4141 (
            .O(N__22252),
            .I(N__22246));
    InMux I__4140 (
            .O(N__22251),
            .I(N__22237));
    CascadeMux I__4139 (
            .O(N__22250),
            .I(N__22234));
    CascadeMux I__4138 (
            .O(N__22249),
            .I(N__22229));
    Span4Mux_v I__4137 (
            .O(N__22246),
            .I(N__22225));
    InMux I__4136 (
            .O(N__22245),
            .I(N__22218));
    InMux I__4135 (
            .O(N__22244),
            .I(N__22218));
    InMux I__4134 (
            .O(N__22243),
            .I(N__22218));
    InMux I__4133 (
            .O(N__22242),
            .I(N__22215));
    InMux I__4132 (
            .O(N__22241),
            .I(N__22212));
    InMux I__4131 (
            .O(N__22240),
            .I(N__22209));
    LocalMux I__4130 (
            .O(N__22237),
            .I(N__22206));
    InMux I__4129 (
            .O(N__22234),
            .I(N__22203));
    InMux I__4128 (
            .O(N__22233),
            .I(N__22200));
    InMux I__4127 (
            .O(N__22232),
            .I(N__22195));
    InMux I__4126 (
            .O(N__22229),
            .I(N__22195));
    InMux I__4125 (
            .O(N__22228),
            .I(N__22192));
    Span4Mux_v I__4124 (
            .O(N__22225),
            .I(N__22185));
    LocalMux I__4123 (
            .O(N__22218),
            .I(N__22182));
    LocalMux I__4122 (
            .O(N__22215),
            .I(N__22179));
    LocalMux I__4121 (
            .O(N__22212),
            .I(N__22176));
    LocalMux I__4120 (
            .O(N__22209),
            .I(N__22173));
    Span4Mux_v I__4119 (
            .O(N__22206),
            .I(N__22168));
    LocalMux I__4118 (
            .O(N__22203),
            .I(N__22168));
    LocalMux I__4117 (
            .O(N__22200),
            .I(N__22162));
    LocalMux I__4116 (
            .O(N__22195),
            .I(N__22162));
    LocalMux I__4115 (
            .O(N__22192),
            .I(N__22159));
    InMux I__4114 (
            .O(N__22191),
            .I(N__22154));
    InMux I__4113 (
            .O(N__22190),
            .I(N__22154));
    InMux I__4112 (
            .O(N__22189),
            .I(N__22149));
    InMux I__4111 (
            .O(N__22188),
            .I(N__22149));
    Span4Mux_s3_h I__4110 (
            .O(N__22185),
            .I(N__22144));
    Span4Mux_s2_v I__4109 (
            .O(N__22182),
            .I(N__22144));
    Span4Mux_h I__4108 (
            .O(N__22179),
            .I(N__22139));
    Span4Mux_h I__4107 (
            .O(N__22176),
            .I(N__22139));
    Span4Mux_h I__4106 (
            .O(N__22173),
            .I(N__22134));
    Span4Mux_h I__4105 (
            .O(N__22168),
            .I(N__22134));
    InMux I__4104 (
            .O(N__22167),
            .I(N__22131));
    Span4Mux_v I__4103 (
            .O(N__22162),
            .I(N__22128));
    Span4Mux_s2_v I__4102 (
            .O(N__22159),
            .I(N__22123));
    LocalMux I__4101 (
            .O(N__22154),
            .I(N__22123));
    LocalMux I__4100 (
            .O(N__22149),
            .I(\tok.n49 ));
    Odrv4 I__4099 (
            .O(N__22144),
            .I(\tok.n49 ));
    Odrv4 I__4098 (
            .O(N__22139),
            .I(\tok.n49 ));
    Odrv4 I__4097 (
            .O(N__22134),
            .I(\tok.n49 ));
    LocalMux I__4096 (
            .O(N__22131),
            .I(\tok.n49 ));
    Odrv4 I__4095 (
            .O(N__22128),
            .I(\tok.n49 ));
    Odrv4 I__4094 (
            .O(N__22123),
            .I(\tok.n49 ));
    CascadeMux I__4093 (
            .O(N__22108),
            .I(\tok.n6380_cascade_ ));
    CascadeMux I__4092 (
            .O(N__22105),
            .I(\tok.n215_adj_656_cascade_ ));
    InMux I__4091 (
            .O(N__22102),
            .I(N__22099));
    LocalMux I__4090 (
            .O(N__22099),
            .I(N__22096));
    Odrv4 I__4089 (
            .O(N__22096),
            .I(\tok.n2665 ));
    CascadeMux I__4088 (
            .O(N__22093),
            .I(N__22090));
    InMux I__4087 (
            .O(N__22090),
            .I(N__22087));
    LocalMux I__4086 (
            .O(N__22087),
            .I(\tok.n4_adj_719 ));
    CascadeMux I__4085 (
            .O(N__22084),
            .I(\tok.n4_adj_719_cascade_ ));
    CascadeMux I__4084 (
            .O(N__22081),
            .I(N__22078));
    InMux I__4083 (
            .O(N__22078),
            .I(N__22075));
    LocalMux I__4082 (
            .O(N__22075),
            .I(N__22072));
    Span12Mux_s7_v I__4081 (
            .O(N__22072),
            .I(N__22069));
    Odrv12 I__4080 (
            .O(N__22069),
            .I(\tok.n10_adj_809 ));
    InMux I__4079 (
            .O(N__22066),
            .I(N__22063));
    LocalMux I__4078 (
            .O(N__22063),
            .I(N__22060));
    Odrv12 I__4077 (
            .O(N__22060),
            .I(\tok.n6411 ));
    InMux I__4076 (
            .O(N__22057),
            .I(N__22054));
    LocalMux I__4075 (
            .O(N__22054),
            .I(N__22051));
    Span4Mux_h I__4074 (
            .O(N__22051),
            .I(N__22048));
    Span4Mux_v I__4073 (
            .O(N__22048),
            .I(N__22045));
    Odrv4 I__4072 (
            .O(N__22045),
            .I(\tok.n6532 ));
    CascadeMux I__4071 (
            .O(N__22042),
            .I(\tok.n207_adj_771_cascade_ ));
    InMux I__4070 (
            .O(N__22039),
            .I(N__22036));
    LocalMux I__4069 (
            .O(N__22036),
            .I(N__22033));
    Odrv12 I__4068 (
            .O(N__22033),
            .I(\tok.n6583 ));
    CascadeMux I__4067 (
            .O(N__22030),
            .I(N__22024));
    InMux I__4066 (
            .O(N__22029),
            .I(N__22021));
    InMux I__4065 (
            .O(N__22028),
            .I(N__22018));
    CascadeMux I__4064 (
            .O(N__22027),
            .I(N__22015));
    InMux I__4063 (
            .O(N__22024),
            .I(N__22011));
    LocalMux I__4062 (
            .O(N__22021),
            .I(N__22006));
    LocalMux I__4061 (
            .O(N__22018),
            .I(N__22006));
    InMux I__4060 (
            .O(N__22015),
            .I(N__22003));
    InMux I__4059 (
            .O(N__22014),
            .I(N__22000));
    LocalMux I__4058 (
            .O(N__22011),
            .I(N__21997));
    Span4Mux_v I__4057 (
            .O(N__22006),
            .I(N__21992));
    LocalMux I__4056 (
            .O(N__22003),
            .I(N__21992));
    LocalMux I__4055 (
            .O(N__22000),
            .I(N__21988));
    Span4Mux_h I__4054 (
            .O(N__21997),
            .I(N__21983));
    Span4Mux_h I__4053 (
            .O(N__21992),
            .I(N__21980));
    InMux I__4052 (
            .O(N__21991),
            .I(N__21977));
    Span4Mux_v I__4051 (
            .O(N__21988),
            .I(N__21974));
    InMux I__4050 (
            .O(N__21987),
            .I(N__21971));
    InMux I__4049 (
            .O(N__21986),
            .I(N__21968));
    Span4Mux_h I__4048 (
            .O(N__21983),
            .I(N__21965));
    Span4Mux_h I__4047 (
            .O(N__21980),
            .I(N__21962));
    LocalMux I__4046 (
            .O(N__21977),
            .I(N__21955));
    Sp12to4 I__4045 (
            .O(N__21974),
            .I(N__21955));
    LocalMux I__4044 (
            .O(N__21971),
            .I(N__21955));
    LocalMux I__4043 (
            .O(N__21968),
            .I(\tok.S_5 ));
    Odrv4 I__4042 (
            .O(N__21965),
            .I(\tok.S_5 ));
    Odrv4 I__4041 (
            .O(N__21962),
            .I(\tok.S_5 ));
    Odrv12 I__4040 (
            .O(N__21955),
            .I(\tok.S_5 ));
    InMux I__4039 (
            .O(N__21946),
            .I(N__21943));
    LocalMux I__4038 (
            .O(N__21943),
            .I(\tok.n213 ));
    CascadeMux I__4037 (
            .O(N__21940),
            .I(\tok.n207_adj_776_cascade_ ));
    CascadeMux I__4036 (
            .O(N__21937),
            .I(\tok.n6529_cascade_ ));
    InMux I__4035 (
            .O(N__21934),
            .I(N__21931));
    LocalMux I__4034 (
            .O(N__21931),
            .I(N__21928));
    Span4Mux_v I__4033 (
            .O(N__21928),
            .I(N__21925));
    Odrv4 I__4032 (
            .O(N__21925),
            .I(\tok.n210_adj_784 ));
    InMux I__4031 (
            .O(N__21922),
            .I(N__21919));
    LocalMux I__4030 (
            .O(N__21919),
            .I(\tok.n174_adj_785 ));
    InMux I__4029 (
            .O(N__21916),
            .I(N__21913));
    LocalMux I__4028 (
            .O(N__21913),
            .I(N__21910));
    Span4Mux_v I__4027 (
            .O(N__21910),
            .I(N__21907));
    Span4Mux_v I__4026 (
            .O(N__21907),
            .I(N__21904));
    Odrv4 I__4025 (
            .O(N__21904),
            .I(\tok.n229_adj_861 ));
    CascadeMux I__4024 (
            .O(N__21901),
            .I(N__21898));
    InMux I__4023 (
            .O(N__21898),
            .I(N__21895));
    LocalMux I__4022 (
            .O(N__21895),
            .I(\tok.n6365 ));
    InMux I__4021 (
            .O(N__21892),
            .I(N__21889));
    LocalMux I__4020 (
            .O(N__21889),
            .I(N__21886));
    Sp12to4 I__4019 (
            .O(N__21886),
            .I(N__21883));
    Odrv12 I__4018 (
            .O(N__21883),
            .I(\tok.n215_adj_672 ));
    InMux I__4017 (
            .O(N__21880),
            .I(N__21877));
    LocalMux I__4016 (
            .O(N__21877),
            .I(N__21874));
    Span4Mux_h I__4015 (
            .O(N__21874),
            .I(N__21871));
    Odrv4 I__4014 (
            .O(N__21871),
            .I(\tok.n252 ));
    CascadeMux I__4013 (
            .O(N__21868),
            .I(\tok.n4_adj_769_cascade_ ));
    InMux I__4012 (
            .O(N__21865),
            .I(N__21862));
    LocalMux I__4011 (
            .O(N__21862),
            .I(\tok.n205_adj_770 ));
    InMux I__4010 (
            .O(N__21859),
            .I(N__21855));
    InMux I__4009 (
            .O(N__21858),
            .I(N__21852));
    LocalMux I__4008 (
            .O(N__21855),
            .I(N__21849));
    LocalMux I__4007 (
            .O(N__21852),
            .I(N__21846));
    Span4Mux_v I__4006 (
            .O(N__21849),
            .I(N__21841));
    Span4Mux_v I__4005 (
            .O(N__21846),
            .I(N__21841));
    Sp12to4 I__4004 (
            .O(N__21841),
            .I(N__21838));
    Odrv12 I__4003 (
            .O(N__21838),
            .I(\tok.n235 ));
    CascadeMux I__4002 (
            .O(N__21835),
            .I(\tok.n190_cascade_ ));
    InMux I__4001 (
            .O(N__21832),
            .I(N__21829));
    LocalMux I__4000 (
            .O(N__21829),
            .I(\tok.n190 ));
    CascadeMux I__3999 (
            .O(N__21826),
            .I(\tok.n255_cascade_ ));
    InMux I__3998 (
            .O(N__21823),
            .I(N__21820));
    LocalMux I__3997 (
            .O(N__21820),
            .I(\tok.n258 ));
    CascadeMux I__3996 (
            .O(N__21817),
            .I(\tok.n6508_cascade_ ));
    InMux I__3995 (
            .O(N__21814),
            .I(N__21811));
    LocalMux I__3994 (
            .O(N__21811),
            .I(\tok.n210_adj_816 ));
    CascadeMux I__3993 (
            .O(N__21808),
            .I(\tok.n872_cascade_ ));
    CascadeMux I__3992 (
            .O(N__21805),
            .I(\tok.n174_adj_817_cascade_ ));
    InMux I__3991 (
            .O(N__21802),
            .I(N__21799));
    LocalMux I__3990 (
            .O(N__21799),
            .I(\tok.n4_adj_818 ));
    InMux I__3989 (
            .O(N__21796),
            .I(N__21793));
    LocalMux I__3988 (
            .O(N__21793),
            .I(\tok.n205_adj_820 ));
    InMux I__3987 (
            .O(N__21790),
            .I(N__21787));
    LocalMux I__3986 (
            .O(N__21787),
            .I(N__21784));
    Odrv12 I__3985 (
            .O(N__21784),
            .I(\tok.n200_adj_840 ));
    CascadeMux I__3984 (
            .O(N__21781),
            .I(\tok.n6_adj_843_cascade_ ));
    InMux I__3983 (
            .O(N__21778),
            .I(N__21774));
    CascadeMux I__3982 (
            .O(N__21777),
            .I(N__21769));
    LocalMux I__3981 (
            .O(N__21774),
            .I(N__21765));
    InMux I__3980 (
            .O(N__21773),
            .I(N__21762));
    CascadeMux I__3979 (
            .O(N__21772),
            .I(N__21758));
    InMux I__3978 (
            .O(N__21769),
            .I(N__21755));
    InMux I__3977 (
            .O(N__21768),
            .I(N__21752));
    Span4Mux_v I__3976 (
            .O(N__21765),
            .I(N__21747));
    LocalMux I__3975 (
            .O(N__21762),
            .I(N__21747));
    InMux I__3974 (
            .O(N__21761),
            .I(N__21744));
    InMux I__3973 (
            .O(N__21758),
            .I(N__21741));
    LocalMux I__3972 (
            .O(N__21755),
            .I(N__21738));
    LocalMux I__3971 (
            .O(N__21752),
            .I(N__21734));
    Span4Mux_h I__3970 (
            .O(N__21747),
            .I(N__21731));
    LocalMux I__3969 (
            .O(N__21744),
            .I(N__21726));
    LocalMux I__3968 (
            .O(N__21741),
            .I(N__21726));
    Span4Mux_v I__3967 (
            .O(N__21738),
            .I(N__21723));
    InMux I__3966 (
            .O(N__21737),
            .I(N__21720));
    Span4Mux_h I__3965 (
            .O(N__21734),
            .I(N__21717));
    Span4Mux_h I__3964 (
            .O(N__21731),
            .I(N__21714));
    Span4Mux_v I__3963 (
            .O(N__21726),
            .I(N__21711));
    Span4Mux_h I__3962 (
            .O(N__21723),
            .I(N__21708));
    LocalMux I__3961 (
            .O(N__21720),
            .I(\tok.S_9 ));
    Odrv4 I__3960 (
            .O(N__21717),
            .I(\tok.S_9 ));
    Odrv4 I__3959 (
            .O(N__21714),
            .I(\tok.S_9 ));
    Odrv4 I__3958 (
            .O(N__21711),
            .I(\tok.S_9 ));
    Odrv4 I__3957 (
            .O(N__21708),
            .I(\tok.S_9 ));
    CascadeMux I__3956 (
            .O(N__21697),
            .I(\tok.n6440_cascade_ ));
    CascadeMux I__3955 (
            .O(N__21694),
            .I(\tok.n6612_cascade_ ));
    CascadeMux I__3954 (
            .O(N__21691),
            .I(\tok.n179_cascade_ ));
    InMux I__3953 (
            .O(N__21688),
            .I(N__21685));
    LocalMux I__3952 (
            .O(N__21685),
            .I(\tok.n6546 ));
    CascadeMux I__3951 (
            .O(N__21682),
            .I(N__21678));
    CascadeMux I__3950 (
            .O(N__21681),
            .I(N__21675));
    InMux I__3949 (
            .O(N__21678),
            .I(N__21672));
    InMux I__3948 (
            .O(N__21675),
            .I(N__21669));
    LocalMux I__3947 (
            .O(N__21672),
            .I(N__21666));
    LocalMux I__3946 (
            .O(N__21669),
            .I(N__21663));
    Span4Mux_v I__3945 (
            .O(N__21666),
            .I(N__21660));
    Span4Mux_v I__3944 (
            .O(N__21663),
            .I(N__21657));
    Span4Mux_h I__3943 (
            .O(N__21660),
            .I(N__21654));
    Span4Mux_v I__3942 (
            .O(N__21657),
            .I(N__21651));
    Odrv4 I__3941 (
            .O(N__21654),
            .I(\tok.table_rd_7 ));
    Odrv4 I__3940 (
            .O(N__21651),
            .I(\tok.table_rd_7 ));
    CascadeMux I__3939 (
            .O(N__21646),
            .I(N__21643));
    InMux I__3938 (
            .O(N__21643),
            .I(N__21639));
    InMux I__3937 (
            .O(N__21642),
            .I(N__21636));
    LocalMux I__3936 (
            .O(N__21639),
            .I(N__21633));
    LocalMux I__3935 (
            .O(N__21636),
            .I(N__21630));
    Span4Mux_v I__3934 (
            .O(N__21633),
            .I(N__21627));
    Span12Mux_s9_v I__3933 (
            .O(N__21630),
            .I(N__21624));
    Span4Mux_h I__3932 (
            .O(N__21627),
            .I(N__21621));
    Odrv12 I__3931 (
            .O(N__21624),
            .I(\tok.table_rd_4 ));
    Odrv4 I__3930 (
            .O(N__21621),
            .I(\tok.table_rd_4 ));
    InMux I__3929 (
            .O(N__21616),
            .I(N__21613));
    LocalMux I__3928 (
            .O(N__21613),
            .I(\tok.n258_adj_814 ));
    CascadeMux I__3927 (
            .O(N__21610),
            .I(\tok.n252_adj_815_cascade_ ));
    InMux I__3926 (
            .O(N__21607),
            .I(N__21603));
    InMux I__3925 (
            .O(N__21606),
            .I(N__21600));
    LocalMux I__3924 (
            .O(N__21603),
            .I(N__21595));
    LocalMux I__3923 (
            .O(N__21600),
            .I(N__21595));
    Span4Mux_v I__3922 (
            .O(N__21595),
            .I(N__21592));
    Span4Mux_h I__3921 (
            .O(N__21592),
            .I(N__21589));
    Odrv4 I__3920 (
            .O(N__21589),
            .I(\tok.n232 ));
    InMux I__3919 (
            .O(N__21586),
            .I(N__21583));
    LocalMux I__3918 (
            .O(N__21583),
            .I(\tok.n255_adj_808 ));
    InMux I__3917 (
            .O(N__21580),
            .I(N__21577));
    LocalMux I__3916 (
            .O(N__21577),
            .I(\tok.n311_adj_721 ));
    CascadeMux I__3915 (
            .O(N__21574),
            .I(\tok.n167_cascade_ ));
    InMux I__3914 (
            .O(N__21571),
            .I(N__21568));
    LocalMux I__3913 (
            .O(N__21568),
            .I(N__21565));
    Odrv4 I__3912 (
            .O(N__21565),
            .I(\tok.n6567 ));
    InMux I__3911 (
            .O(N__21562),
            .I(N__21558));
    CascadeMux I__3910 (
            .O(N__21561),
            .I(N__21555));
    LocalMux I__3909 (
            .O(N__21558),
            .I(N__21552));
    InMux I__3908 (
            .O(N__21555),
            .I(N__21549));
    Span4Mux_v I__3907 (
            .O(N__21552),
            .I(N__21544));
    LocalMux I__3906 (
            .O(N__21549),
            .I(N__21544));
    Span4Mux_v I__3905 (
            .O(N__21544),
            .I(N__21541));
    Span4Mux_h I__3904 (
            .O(N__21541),
            .I(N__21538));
    Odrv4 I__3903 (
            .O(N__21538),
            .I(\tok.table_rd_2 ));
    CascadeMux I__3902 (
            .O(N__21535),
            .I(\tok.n209_cascade_ ));
    CascadeMux I__3901 (
            .O(N__21532),
            .I(\tok.n6625_cascade_ ));
    InMux I__3900 (
            .O(N__21529),
            .I(N__21526));
    LocalMux I__3899 (
            .O(N__21526),
            .I(\tok.n6624 ));
    CascadeMux I__3898 (
            .O(N__21523),
            .I(\tok.n168_adj_700_cascade_ ));
    InMux I__3897 (
            .O(N__21520),
            .I(N__21517));
    LocalMux I__3896 (
            .O(N__21517),
            .I(\tok.n6569 ));
    InMux I__3895 (
            .O(N__21514),
            .I(N__21511));
    LocalMux I__3894 (
            .O(N__21511),
            .I(N__21508));
    Span4Mux_h I__3893 (
            .O(N__21508),
            .I(N__21505));
    Odrv4 I__3892 (
            .O(N__21505),
            .I(\tok.n2548 ));
    CascadeMux I__3891 (
            .O(N__21502),
            .I(N__21499));
    InMux I__3890 (
            .O(N__21499),
            .I(N__21496));
    LocalMux I__3889 (
            .O(N__21496),
            .I(N__21493));
    Span4Mux_v I__3888 (
            .O(N__21493),
            .I(N__21490));
    Odrv4 I__3887 (
            .O(N__21490),
            .I(\tok.n6396 ));
    InMux I__3886 (
            .O(N__21487),
            .I(N__21481));
    InMux I__3885 (
            .O(N__21486),
            .I(N__21481));
    LocalMux I__3884 (
            .O(N__21481),
            .I(N__21477));
    InMux I__3883 (
            .O(N__21480),
            .I(N__21474));
    Span4Mux_v I__3882 (
            .O(N__21477),
            .I(N__21471));
    LocalMux I__3881 (
            .O(N__21474),
            .I(N__21468));
    Span4Mux_v I__3880 (
            .O(N__21471),
            .I(N__21465));
    Span4Mux_h I__3879 (
            .O(N__21468),
            .I(N__21462));
    Span4Mux_h I__3878 (
            .O(N__21465),
            .I(N__21459));
    Span4Mux_h I__3877 (
            .O(N__21462),
            .I(N__21456));
    Odrv4 I__3876 (
            .O(N__21459),
            .I(\tok.n236 ));
    Odrv4 I__3875 (
            .O(N__21456),
            .I(\tok.n236 ));
    InMux I__3874 (
            .O(N__21451),
            .I(N__21448));
    LocalMux I__3873 (
            .O(N__21448),
            .I(\tok.n4925 ));
    InMux I__3872 (
            .O(N__21445),
            .I(N__21442));
    LocalMux I__3871 (
            .O(N__21442),
            .I(N__21439));
    Span4Mux_h I__3870 (
            .O(N__21439),
            .I(N__21436));
    Odrv4 I__3869 (
            .O(N__21436),
            .I(\tok.n288 ));
    InMux I__3868 (
            .O(N__21433),
            .I(N__21430));
    LocalMux I__3867 (
            .O(N__21430),
            .I(N__21427));
    Span4Mux_v I__3866 (
            .O(N__21427),
            .I(N__21424));
    Span4Mux_h I__3865 (
            .O(N__21424),
            .I(N__21421));
    Odrv4 I__3864 (
            .O(N__21421),
            .I(\tok.n2613 ));
    CascadeMux I__3863 (
            .O(N__21418),
            .I(\tok.n6578_cascade_ ));
    InMux I__3862 (
            .O(N__21415),
            .I(N__21412));
    LocalMux I__3861 (
            .O(N__21412),
            .I(N__21409));
    Odrv4 I__3860 (
            .O(N__21409),
            .I(\tok.n6581 ));
    InMux I__3859 (
            .O(N__21406),
            .I(N__21403));
    LocalMux I__3858 (
            .O(N__21403),
            .I(\tok.n4_adj_739 ));
    InMux I__3857 (
            .O(N__21400),
            .I(N__21397));
    LocalMux I__3856 (
            .O(N__21397),
            .I(\tok.n2611 ));
    InMux I__3855 (
            .O(N__21394),
            .I(N__21391));
    LocalMux I__3854 (
            .O(N__21391),
            .I(N__21388));
    Span4Mux_h I__3853 (
            .O(N__21388),
            .I(N__21385));
    Odrv4 I__3852 (
            .O(N__21385),
            .I(\tok.n6580 ));
    InMux I__3851 (
            .O(N__21382),
            .I(N__21376));
    InMux I__3850 (
            .O(N__21381),
            .I(N__21376));
    LocalMux I__3849 (
            .O(N__21376),
            .I(\tok.n4_adj_684 ));
    CascadeMux I__3848 (
            .O(N__21373),
            .I(\tok.n6620_cascade_ ));
    CascadeMux I__3847 (
            .O(N__21370),
            .I(\tok.n14_adj_683_cascade_ ));
    InMux I__3846 (
            .O(N__21367),
            .I(N__21364));
    LocalMux I__3845 (
            .O(N__21364),
            .I(N__21360));
    InMux I__3844 (
            .O(N__21363),
            .I(N__21357));
    Odrv4 I__3843 (
            .O(N__21360),
            .I(\tok.n9_adj_651 ));
    LocalMux I__3842 (
            .O(N__21357),
            .I(\tok.n9_adj_651 ));
    CascadeMux I__3841 (
            .O(N__21352),
            .I(\tok.n15_adj_807_cascade_ ));
    InMux I__3840 (
            .O(N__21349),
            .I(N__21343));
    InMux I__3839 (
            .O(N__21348),
            .I(N__21343));
    LocalMux I__3838 (
            .O(N__21343),
            .I(N__21340));
    Odrv12 I__3837 (
            .O(N__21340),
            .I(\tok.n903 ));
    CascadeMux I__3836 (
            .O(N__21337),
            .I(N__21334));
    InMux I__3835 (
            .O(N__21334),
            .I(N__21331));
    LocalMux I__3834 (
            .O(N__21331),
            .I(N__21328));
    Odrv4 I__3833 (
            .O(N__21328),
            .I(\tok.n14_adj_683 ));
    CascadeMux I__3832 (
            .O(N__21325),
            .I(N__21322));
    InMux I__3831 (
            .O(N__21322),
            .I(N__21319));
    LocalMux I__3830 (
            .O(N__21319),
            .I(\tok.n6621 ));
    InMux I__3829 (
            .O(N__21316),
            .I(N__21313));
    LocalMux I__3828 (
            .O(N__21313),
            .I(\tok.n241_adj_747 ));
    InMux I__3827 (
            .O(N__21310),
            .I(N__21307));
    LocalMux I__3826 (
            .O(N__21307),
            .I(N__21304));
    Odrv4 I__3825 (
            .O(N__21304),
            .I(\tok.n6593 ));
    InMux I__3824 (
            .O(N__21301),
            .I(N__21298));
    LocalMux I__3823 (
            .O(N__21298),
            .I(\tok.n6664 ));
    CascadeMux I__3822 (
            .O(N__21295),
            .I(\tok.n1600_cascade_ ));
    InMux I__3821 (
            .O(N__21292),
            .I(N__21289));
    LocalMux I__3820 (
            .O(N__21289),
            .I(\tok.n13_adj_742 ));
    CascadeMux I__3819 (
            .O(N__21286),
            .I(\tok.n6301_cascade_ ));
    CascadeMux I__3818 (
            .O(N__21283),
            .I(\tok.n80_adj_751_cascade_ ));
    CascadeMux I__3817 (
            .O(N__21280),
            .I(\tok.n83_adj_746_cascade_ ));
    InMux I__3816 (
            .O(N__21277),
            .I(N__21274));
    LocalMux I__3815 (
            .O(N__21274),
            .I(\tok.n6297 ));
    InMux I__3814 (
            .O(N__21271),
            .I(N__21268));
    LocalMux I__3813 (
            .O(N__21268),
            .I(\tok.n89_adj_754 ));
    InMux I__3812 (
            .O(N__21265),
            .I(N__21261));
    InMux I__3811 (
            .O(N__21264),
            .I(N__21258));
    LocalMux I__3810 (
            .O(N__21261),
            .I(N__21255));
    LocalMux I__3809 (
            .O(N__21258),
            .I(N__21252));
    Span4Mux_h I__3808 (
            .O(N__21255),
            .I(N__21249));
    Odrv4 I__3807 (
            .O(N__21252),
            .I(n92_adj_898));
    Odrv4 I__3806 (
            .O(N__21249),
            .I(n92_adj_898));
    CascadeMux I__3805 (
            .O(N__21244),
            .I(N__21240));
    InMux I__3804 (
            .O(N__21243),
            .I(N__21235));
    InMux I__3803 (
            .O(N__21240),
            .I(N__21235));
    LocalMux I__3802 (
            .O(N__21235),
            .I(N__21232));
    Span4Mux_h I__3801 (
            .O(N__21232),
            .I(N__21229));
    Span4Mux_h I__3800 (
            .O(N__21229),
            .I(N__21226));
    Span4Mux_v I__3799 (
            .O(N__21226),
            .I(N__21223));
    Odrv4 I__3798 (
            .O(N__21223),
            .I(\tok.table_rd_3 ));
    InMux I__3797 (
            .O(N__21220),
            .I(N__21214));
    InMux I__3796 (
            .O(N__21219),
            .I(N__21214));
    LocalMux I__3795 (
            .O(N__21214),
            .I(\tok.tail_28 ));
    InMux I__3794 (
            .O(N__21211),
            .I(N__21205));
    InMux I__3793 (
            .O(N__21210),
            .I(N__21205));
    LocalMux I__3792 (
            .O(N__21205),
            .I(\tok.C_stk.tail_36 ));
    CascadeMux I__3791 (
            .O(N__21202),
            .I(\tok.n83_adj_723_cascade_ ));
    InMux I__3790 (
            .O(N__21199),
            .I(N__21195));
    CascadeMux I__3789 (
            .O(N__21198),
            .I(N__21192));
    LocalMux I__3788 (
            .O(N__21195),
            .I(N__21189));
    InMux I__3787 (
            .O(N__21192),
            .I(N__21186));
    Span4Mux_s1_v I__3786 (
            .O(N__21189),
            .I(N__21181));
    LocalMux I__3785 (
            .O(N__21186),
            .I(N__21181));
    Odrv4 I__3784 (
            .O(N__21181),
            .I(n10_adj_908));
    CascadeMux I__3783 (
            .O(N__21178),
            .I(\tok.n4_adj_726_cascade_ ));
    CascadeMux I__3782 (
            .O(N__21175),
            .I(\tok.ram.n6257_cascade_ ));
    InMux I__3781 (
            .O(N__21172),
            .I(N__21168));
    InMux I__3780 (
            .O(N__21171),
            .I(N__21164));
    LocalMux I__3779 (
            .O(N__21168),
            .I(N__21161));
    CascadeMux I__3778 (
            .O(N__21167),
            .I(N__21157));
    LocalMux I__3777 (
            .O(N__21164),
            .I(N__21154));
    Span4Mux_v I__3776 (
            .O(N__21161),
            .I(N__21151));
    InMux I__3775 (
            .O(N__21160),
            .I(N__21146));
    InMux I__3774 (
            .O(N__21157),
            .I(N__21146));
    Span4Mux_s1_v I__3773 (
            .O(N__21154),
            .I(N__21143));
    Span4Mux_h I__3772 (
            .O(N__21151),
            .I(N__21138));
    LocalMux I__3771 (
            .O(N__21146),
            .I(N__21138));
    Odrv4 I__3770 (
            .O(N__21143),
            .I(tc_plus_1_0));
    Odrv4 I__3769 (
            .O(N__21138),
            .I(tc_plus_1_0));
    CascadeMux I__3768 (
            .O(N__21133),
            .I(\tok.C_stk.n6230_cascade_ ));
    InMux I__3767 (
            .O(N__21130),
            .I(N__21125));
    InMux I__3766 (
            .O(N__21129),
            .I(N__21121));
    InMux I__3765 (
            .O(N__21128),
            .I(N__21118));
    LocalMux I__3764 (
            .O(N__21125),
            .I(N__21115));
    InMux I__3763 (
            .O(N__21124),
            .I(N__21112));
    LocalMux I__3762 (
            .O(N__21121),
            .I(tc_0));
    LocalMux I__3761 (
            .O(N__21118),
            .I(tc_0));
    Odrv12 I__3760 (
            .O(N__21115),
            .I(tc_0));
    LocalMux I__3759 (
            .O(N__21112),
            .I(tc_0));
    CascadeMux I__3758 (
            .O(N__21103),
            .I(N__21098));
    InMux I__3757 (
            .O(N__21102),
            .I(N__21095));
    InMux I__3756 (
            .O(N__21101),
            .I(N__21090));
    InMux I__3755 (
            .O(N__21098),
            .I(N__21090));
    LocalMux I__3754 (
            .O(N__21095),
            .I(N__21084));
    LocalMux I__3753 (
            .O(N__21090),
            .I(N__21084));
    InMux I__3752 (
            .O(N__21089),
            .I(N__21081));
    Span4Mux_h I__3751 (
            .O(N__21084),
            .I(N__21078));
    LocalMux I__3750 (
            .O(N__21081),
            .I(c_stk_r_0));
    Odrv4 I__3749 (
            .O(N__21078),
            .I(c_stk_r_0));
    CascadeMux I__3748 (
            .O(N__21073),
            .I(N__21070));
    InMux I__3747 (
            .O(N__21070),
            .I(N__21064));
    InMux I__3746 (
            .O(N__21069),
            .I(N__21064));
    LocalMux I__3745 (
            .O(N__21064),
            .I(\tok.C_stk.tail_0 ));
    InMux I__3744 (
            .O(N__21061),
            .I(N__21058));
    LocalMux I__3743 (
            .O(N__21058),
            .I(N__21052));
    InMux I__3742 (
            .O(N__21057),
            .I(N__21049));
    InMux I__3741 (
            .O(N__21056),
            .I(N__21044));
    InMux I__3740 (
            .O(N__21055),
            .I(N__21044));
    Odrv4 I__3739 (
            .O(N__21052),
            .I(\tok.tc_plus_1_4 ));
    LocalMux I__3738 (
            .O(N__21049),
            .I(\tok.tc_plus_1_4 ));
    LocalMux I__3737 (
            .O(N__21044),
            .I(\tok.tc_plus_1_4 ));
    CascadeMux I__3736 (
            .O(N__21037),
            .I(\tok.C_stk.n6239_cascade_ ));
    CascadeMux I__3735 (
            .O(N__21034),
            .I(N__21030));
    InMux I__3734 (
            .O(N__21033),
            .I(N__21025));
    InMux I__3733 (
            .O(N__21030),
            .I(N__21020));
    InMux I__3732 (
            .O(N__21029),
            .I(N__21020));
    InMux I__3731 (
            .O(N__21028),
            .I(N__21017));
    LocalMux I__3730 (
            .O(N__21025),
            .I(tc_4));
    LocalMux I__3729 (
            .O(N__21020),
            .I(tc_4));
    LocalMux I__3728 (
            .O(N__21017),
            .I(tc_4));
    CascadeMux I__3727 (
            .O(N__21010),
            .I(N__21005));
    InMux I__3726 (
            .O(N__21009),
            .I(N__21001));
    InMux I__3725 (
            .O(N__21008),
            .I(N__20998));
    InMux I__3724 (
            .O(N__21005),
            .I(N__20993));
    InMux I__3723 (
            .O(N__21004),
            .I(N__20993));
    LocalMux I__3722 (
            .O(N__21001),
            .I(\tok.c_stk_r_4 ));
    LocalMux I__3721 (
            .O(N__20998),
            .I(\tok.c_stk_r_4 ));
    LocalMux I__3720 (
            .O(N__20993),
            .I(\tok.c_stk_r_4 ));
    InMux I__3719 (
            .O(N__20986),
            .I(N__20980));
    InMux I__3718 (
            .O(N__20985),
            .I(N__20980));
    LocalMux I__3717 (
            .O(N__20980),
            .I(\tok.C_stk.tail_4 ));
    InMux I__3716 (
            .O(N__20977),
            .I(N__20971));
    InMux I__3715 (
            .O(N__20976),
            .I(N__20971));
    LocalMux I__3714 (
            .O(N__20971),
            .I(\tok.tail_12 ));
    CascadeMux I__3713 (
            .O(N__20968),
            .I(N__20965));
    InMux I__3712 (
            .O(N__20965),
            .I(N__20959));
    InMux I__3711 (
            .O(N__20964),
            .I(N__20959));
    LocalMux I__3710 (
            .O(N__20959),
            .I(\tok.C_stk.tail_20 ));
    InMux I__3709 (
            .O(N__20956),
            .I(N__20953));
    LocalMux I__3708 (
            .O(N__20953),
            .I(\tok.n6425 ));
    InMux I__3707 (
            .O(N__20950),
            .I(N__20947));
    LocalMux I__3706 (
            .O(N__20947),
            .I(\tok.n6346 ));
    InMux I__3705 (
            .O(N__20944),
            .I(N__20941));
    LocalMux I__3704 (
            .O(N__20941),
            .I(N__20938));
    Odrv12 I__3703 (
            .O(N__20938),
            .I(\tok.n215_adj_876 ));
    InMux I__3702 (
            .O(N__20935),
            .I(N__20932));
    LocalMux I__3701 (
            .O(N__20932),
            .I(\tok.n179_adj_877 ));
    CascadeMux I__3700 (
            .O(N__20929),
            .I(\tok.n6553_cascade_ ));
    InMux I__3699 (
            .O(N__20926),
            .I(N__20923));
    LocalMux I__3698 (
            .O(N__20923),
            .I(N__20920));
    Span4Mux_v I__3697 (
            .O(N__20920),
            .I(N__20917));
    Odrv4 I__3696 (
            .O(N__20917),
            .I(\tok.n6552 ));
    InMux I__3695 (
            .O(N__20914),
            .I(N__20911));
    LocalMux I__3694 (
            .O(N__20911),
            .I(\tok.n179_adj_698 ));
    InMux I__3693 (
            .O(N__20908),
            .I(N__20905));
    LocalMux I__3692 (
            .O(N__20905),
            .I(N__20902));
    Odrv12 I__3691 (
            .O(N__20902),
            .I(\tok.n6537 ));
    CascadeMux I__3690 (
            .O(N__20899),
            .I(\tok.n6541_cascade_ ));
    InMux I__3689 (
            .O(N__20896),
            .I(N__20893));
    LocalMux I__3688 (
            .O(N__20893),
            .I(N__20890));
    Span4Mux_h I__3687 (
            .O(N__20890),
            .I(N__20887));
    Odrv4 I__3686 (
            .O(N__20887),
            .I(\tok.n6540 ));
    InMux I__3685 (
            .O(N__20884),
            .I(N__20881));
    LocalMux I__3684 (
            .O(N__20881),
            .I(N__20878));
    Odrv4 I__3683 (
            .O(N__20878),
            .I(\tok.n6367 ));
    InMux I__3682 (
            .O(N__20875),
            .I(N__20872));
    LocalMux I__3681 (
            .O(N__20872),
            .I(\tok.n179_adj_673 ));
    InMux I__3680 (
            .O(N__20869),
            .I(N__20866));
    LocalMux I__3679 (
            .O(N__20866),
            .I(\tok.uart.sender_4 ));
    InMux I__3678 (
            .O(N__20863),
            .I(N__20860));
    LocalMux I__3677 (
            .O(N__20860),
            .I(N__20857));
    Span4Mux_s2_v I__3676 (
            .O(N__20857),
            .I(N__20854));
    Odrv4 I__3675 (
            .O(N__20854),
            .I(\tok.uart.sender_3 ));
    CascadeMux I__3674 (
            .O(N__20851),
            .I(N__20848));
    InMux I__3673 (
            .O(N__20848),
            .I(N__20845));
    LocalMux I__3672 (
            .O(N__20845),
            .I(N__20842));
    Span4Mux_h I__3671 (
            .O(N__20842),
            .I(N__20839));
    Odrv4 I__3670 (
            .O(N__20839),
            .I(\tok.n2602 ));
    InMux I__3669 (
            .O(N__20836),
            .I(N__20833));
    LocalMux I__3668 (
            .O(N__20833),
            .I(\tok.n6450 ));
    CascadeMux I__3667 (
            .O(N__20830),
            .I(\tok.n215_adj_830_cascade_ ));
    CascadeMux I__3666 (
            .O(N__20827),
            .I(\tok.n6605_cascade_ ));
    InMux I__3665 (
            .O(N__20824),
            .I(N__20821));
    LocalMux I__3664 (
            .O(N__20821),
            .I(N__20818));
    Span4Mux_h I__3663 (
            .O(N__20818),
            .I(N__20815));
    Odrv4 I__3662 (
            .O(N__20815),
            .I(\tok.n6604 ));
    InMux I__3661 (
            .O(N__20812),
            .I(N__20809));
    LocalMux I__3660 (
            .O(N__20809),
            .I(N__20806));
    Span4Mux_h I__3659 (
            .O(N__20806),
            .I(N__20803));
    Odrv4 I__3658 (
            .O(N__20803),
            .I(\tok.n6456 ));
    InMux I__3657 (
            .O(N__20800),
            .I(N__20797));
    LocalMux I__3656 (
            .O(N__20797),
            .I(\tok.n179_adj_831 ));
    InMux I__3655 (
            .O(N__20794),
            .I(N__20789));
    InMux I__3654 (
            .O(N__20793),
            .I(N__20786));
    CascadeMux I__3653 (
            .O(N__20792),
            .I(N__20782));
    LocalMux I__3652 (
            .O(N__20789),
            .I(N__20778));
    LocalMux I__3651 (
            .O(N__20786),
            .I(N__20775));
    InMux I__3650 (
            .O(N__20785),
            .I(N__20770));
    InMux I__3649 (
            .O(N__20782),
            .I(N__20770));
    CascadeMux I__3648 (
            .O(N__20781),
            .I(N__20762));
    Span4Mux_h I__3647 (
            .O(N__20778),
            .I(N__20751));
    Span4Mux_h I__3646 (
            .O(N__20775),
            .I(N__20751));
    LocalMux I__3645 (
            .O(N__20770),
            .I(N__20751));
    InMux I__3644 (
            .O(N__20769),
            .I(N__20748));
    InMux I__3643 (
            .O(N__20768),
            .I(N__20741));
    InMux I__3642 (
            .O(N__20767),
            .I(N__20741));
    InMux I__3641 (
            .O(N__20766),
            .I(N__20741));
    InMux I__3640 (
            .O(N__20765),
            .I(N__20737));
    InMux I__3639 (
            .O(N__20762),
            .I(N__20734));
    InMux I__3638 (
            .O(N__20761),
            .I(N__20731));
    InMux I__3637 (
            .O(N__20760),
            .I(N__20724));
    InMux I__3636 (
            .O(N__20759),
            .I(N__20724));
    InMux I__3635 (
            .O(N__20758),
            .I(N__20724));
    Span4Mux_h I__3634 (
            .O(N__20751),
            .I(N__20721));
    LocalMux I__3633 (
            .O(N__20748),
            .I(N__20716));
    LocalMux I__3632 (
            .O(N__20741),
            .I(N__20716));
    InMux I__3631 (
            .O(N__20740),
            .I(N__20713));
    LocalMux I__3630 (
            .O(N__20737),
            .I(\tok.n214 ));
    LocalMux I__3629 (
            .O(N__20734),
            .I(\tok.n214 ));
    LocalMux I__3628 (
            .O(N__20731),
            .I(\tok.n214 ));
    LocalMux I__3627 (
            .O(N__20724),
            .I(\tok.n214 ));
    Odrv4 I__3626 (
            .O(N__20721),
            .I(\tok.n214 ));
    Odrv4 I__3625 (
            .O(N__20716),
            .I(\tok.n214 ));
    LocalMux I__3624 (
            .O(N__20713),
            .I(\tok.n214 ));
    CascadeMux I__3623 (
            .O(N__20698),
            .I(\tok.n6462_cascade_ ));
    InMux I__3622 (
            .O(N__20695),
            .I(N__20692));
    LocalMux I__3621 (
            .O(N__20692),
            .I(N__20686));
    InMux I__3620 (
            .O(N__20691),
            .I(N__20683));
    InMux I__3619 (
            .O(N__20690),
            .I(N__20680));
    InMux I__3618 (
            .O(N__20689),
            .I(N__20674));
    Span4Mux_v I__3617 (
            .O(N__20686),
            .I(N__20671));
    LocalMux I__3616 (
            .O(N__20683),
            .I(N__20665));
    LocalMux I__3615 (
            .O(N__20680),
            .I(N__20665));
    InMux I__3614 (
            .O(N__20679),
            .I(N__20660));
    InMux I__3613 (
            .O(N__20678),
            .I(N__20660));
    InMux I__3612 (
            .O(N__20677),
            .I(N__20657));
    LocalMux I__3611 (
            .O(N__20674),
            .I(N__20653));
    Span4Mux_v I__3610 (
            .O(N__20671),
            .I(N__20650));
    InMux I__3609 (
            .O(N__20670),
            .I(N__20647));
    Span12Mux_s11_h I__3608 (
            .O(N__20665),
            .I(N__20644));
    LocalMux I__3607 (
            .O(N__20660),
            .I(N__20639));
    LocalMux I__3606 (
            .O(N__20657),
            .I(N__20639));
    InMux I__3605 (
            .O(N__20656),
            .I(N__20636));
    Span4Mux_s2_h I__3604 (
            .O(N__20653),
            .I(N__20633));
    Odrv4 I__3603 (
            .O(N__20650),
            .I(\tok.n786 ));
    LocalMux I__3602 (
            .O(N__20647),
            .I(\tok.n786 ));
    Odrv12 I__3601 (
            .O(N__20644),
            .I(\tok.n786 ));
    Odrv4 I__3600 (
            .O(N__20639),
            .I(\tok.n786 ));
    LocalMux I__3599 (
            .O(N__20636),
            .I(\tok.n786 ));
    Odrv4 I__3598 (
            .O(N__20633),
            .I(\tok.n786 ));
    InMux I__3597 (
            .O(N__20620),
            .I(N__20617));
    LocalMux I__3596 (
            .O(N__20617),
            .I(\tok.n206_adj_823 ));
    CascadeMux I__3595 (
            .O(N__20614),
            .I(N__20611));
    InMux I__3594 (
            .O(N__20611),
            .I(N__20607));
    InMux I__3593 (
            .O(N__20610),
            .I(N__20604));
    LocalMux I__3592 (
            .O(N__20607),
            .I(N__20601));
    LocalMux I__3591 (
            .O(N__20604),
            .I(N__20598));
    Span4Mux_h I__3590 (
            .O(N__20601),
            .I(N__20595));
    Span4Mux_h I__3589 (
            .O(N__20598),
            .I(N__20590));
    Span4Mux_v I__3588 (
            .O(N__20595),
            .I(N__20590));
    Odrv4 I__3587 (
            .O(N__20590),
            .I(\tok.n314 ));
    InMux I__3586 (
            .O(N__20587),
            .I(N__20584));
    LocalMux I__3585 (
            .O(N__20584),
            .I(N__20581));
    Span4Mux_v I__3584 (
            .O(N__20581),
            .I(N__20578));
    Odrv4 I__3583 (
            .O(N__20578),
            .I(\tok.n321 ));
    InMux I__3582 (
            .O(N__20575),
            .I(N__20566));
    InMux I__3581 (
            .O(N__20574),
            .I(N__20566));
    InMux I__3580 (
            .O(N__20573),
            .I(N__20566));
    LocalMux I__3579 (
            .O(N__20566),
            .I(N__20563));
    Odrv4 I__3578 (
            .O(N__20563),
            .I(\tok.n4_adj_640 ));
    InMux I__3577 (
            .O(N__20560),
            .I(N__20553));
    InMux I__3576 (
            .O(N__20559),
            .I(N__20553));
    CascadeMux I__3575 (
            .O(N__20558),
            .I(N__20550));
    LocalMux I__3574 (
            .O(N__20553),
            .I(N__20547));
    InMux I__3573 (
            .O(N__20550),
            .I(N__20544));
    Span4Mux_h I__3572 (
            .O(N__20547),
            .I(N__20541));
    LocalMux I__3571 (
            .O(N__20544),
            .I(N__20538));
    Span4Mux_v I__3570 (
            .O(N__20541),
            .I(N__20535));
    Odrv4 I__3569 (
            .O(N__20538),
            .I(\tok.n4_adj_680 ));
    Odrv4 I__3568 (
            .O(N__20535),
            .I(\tok.n4_adj_680 ));
    InMux I__3567 (
            .O(N__20530),
            .I(N__20527));
    LocalMux I__3566 (
            .O(N__20527),
            .I(N__20524));
    Span4Mux_v I__3565 (
            .O(N__20524),
            .I(N__20521));
    Odrv4 I__3564 (
            .O(N__20521),
            .I(\tok.n239_adj_679 ));
    CascadeMux I__3563 (
            .O(N__20518),
            .I(\tok.n238_adj_681_cascade_ ));
    InMux I__3562 (
            .O(N__20515),
            .I(N__20511));
    InMux I__3561 (
            .O(N__20514),
            .I(N__20508));
    LocalMux I__3560 (
            .O(N__20511),
            .I(N__20505));
    LocalMux I__3559 (
            .O(N__20508),
            .I(\tok.n900 ));
    Odrv12 I__3558 (
            .O(N__20505),
            .I(\tok.n900 ));
    InMux I__3557 (
            .O(N__20500),
            .I(N__20497));
    LocalMux I__3556 (
            .O(N__20497),
            .I(N__20494));
    Span4Mux_v I__3555 (
            .O(N__20494),
            .I(N__20491));
    Odrv4 I__3554 (
            .O(N__20491),
            .I(\tok.n317_adj_659 ));
    InMux I__3553 (
            .O(N__20488),
            .I(N__20485));
    LocalMux I__3552 (
            .O(N__20485),
            .I(N__20482));
    Odrv12 I__3551 (
            .O(N__20482),
            .I(\tok.n2663 ));
    InMux I__3550 (
            .O(N__20479),
            .I(N__20476));
    LocalMux I__3549 (
            .O(N__20476),
            .I(\tok.uart.sender_5 ));
    CascadeMux I__3548 (
            .O(N__20473),
            .I(\tok.n2600_cascade_ ));
    CascadeMux I__3547 (
            .O(N__20470),
            .I(\tok.n6610_cascade_ ));
    CascadeMux I__3546 (
            .O(N__20467),
            .I(N__20464));
    InMux I__3545 (
            .O(N__20464),
            .I(N__20461));
    LocalMux I__3544 (
            .O(N__20461),
            .I(\tok.n6344 ));
    CascadeMux I__3543 (
            .O(N__20458),
            .I(\tok.n269_cascade_ ));
    CascadeMux I__3542 (
            .O(N__20455),
            .I(N__20452));
    InMux I__3541 (
            .O(N__20452),
            .I(N__20449));
    LocalMux I__3540 (
            .O(N__20449),
            .I(\tok.n4_adj_786 ));
    InMux I__3539 (
            .O(N__20446),
            .I(N__20443));
    LocalMux I__3538 (
            .O(N__20443),
            .I(N__20440));
    Odrv4 I__3537 (
            .O(N__20440),
            .I(\tok.n205_adj_789 ));
    InMux I__3536 (
            .O(N__20437),
            .I(N__20434));
    LocalMux I__3535 (
            .O(N__20434),
            .I(N__20430));
    CascadeMux I__3534 (
            .O(N__20433),
            .I(N__20427));
    Span4Mux_v I__3533 (
            .O(N__20430),
            .I(N__20422));
    InMux I__3532 (
            .O(N__20427),
            .I(N__20417));
    InMux I__3531 (
            .O(N__20426),
            .I(N__20417));
    CascadeMux I__3530 (
            .O(N__20425),
            .I(N__20413));
    Span4Mux_h I__3529 (
            .O(N__20422),
            .I(N__20407));
    LocalMux I__3528 (
            .O(N__20417),
            .I(N__20407));
    CascadeMux I__3527 (
            .O(N__20416),
            .I(N__20401));
    InMux I__3526 (
            .O(N__20413),
            .I(N__20397));
    CascadeMux I__3525 (
            .O(N__20412),
            .I(N__20393));
    Span4Mux_h I__3524 (
            .O(N__20407),
            .I(N__20390));
    CascadeMux I__3523 (
            .O(N__20406),
            .I(N__20387));
    CascadeMux I__3522 (
            .O(N__20405),
            .I(N__20384));
    InMux I__3521 (
            .O(N__20404),
            .I(N__20377));
    InMux I__3520 (
            .O(N__20401),
            .I(N__20377));
    InMux I__3519 (
            .O(N__20400),
            .I(N__20377));
    LocalMux I__3518 (
            .O(N__20397),
            .I(N__20374));
    InMux I__3517 (
            .O(N__20396),
            .I(N__20369));
    InMux I__3516 (
            .O(N__20393),
            .I(N__20369));
    Span4Mux_h I__3515 (
            .O(N__20390),
            .I(N__20366));
    InMux I__3514 (
            .O(N__20387),
            .I(N__20361));
    InMux I__3513 (
            .O(N__20384),
            .I(N__20361));
    LocalMux I__3512 (
            .O(N__20377),
            .I(N__20356));
    Span4Mux_h I__3511 (
            .O(N__20374),
            .I(N__20356));
    LocalMux I__3510 (
            .O(N__20369),
            .I(\tok.n4_adj_635 ));
    Odrv4 I__3509 (
            .O(N__20366),
            .I(\tok.n4_adj_635 ));
    LocalMux I__3508 (
            .O(N__20361),
            .I(\tok.n4_adj_635 ));
    Odrv4 I__3507 (
            .O(N__20356),
            .I(\tok.n4_adj_635 ));
    CascadeMux I__3506 (
            .O(N__20347),
            .I(\tok.n6341_cascade_ ));
    InMux I__3505 (
            .O(N__20344),
            .I(N__20336));
    InMux I__3504 (
            .O(N__20343),
            .I(N__20329));
    InMux I__3503 (
            .O(N__20342),
            .I(N__20329));
    InMux I__3502 (
            .O(N__20341),
            .I(N__20329));
    InMux I__3501 (
            .O(N__20340),
            .I(N__20326));
    InMux I__3500 (
            .O(N__20339),
            .I(N__20323));
    LocalMux I__3499 (
            .O(N__20336),
            .I(N__20318));
    LocalMux I__3498 (
            .O(N__20329),
            .I(N__20315));
    LocalMux I__3497 (
            .O(N__20326),
            .I(N__20310));
    LocalMux I__3496 (
            .O(N__20323),
            .I(N__20310));
    InMux I__3495 (
            .O(N__20322),
            .I(N__20307));
    InMux I__3494 (
            .O(N__20321),
            .I(N__20304));
    Span4Mux_s3_v I__3493 (
            .O(N__20318),
            .I(N__20301));
    Span4Mux_s3_v I__3492 (
            .O(N__20315),
            .I(N__20298));
    Span4Mux_s3_v I__3491 (
            .O(N__20310),
            .I(N__20291));
    LocalMux I__3490 (
            .O(N__20307),
            .I(N__20291));
    LocalMux I__3489 (
            .O(N__20304),
            .I(N__20291));
    Odrv4 I__3488 (
            .O(N__20301),
            .I(\tok.n170 ));
    Odrv4 I__3487 (
            .O(N__20298),
            .I(\tok.n170 ));
    Odrv4 I__3486 (
            .O(N__20291),
            .I(\tok.n170 ));
    InMux I__3485 (
            .O(N__20284),
            .I(N__20281));
    LocalMux I__3484 (
            .O(N__20281),
            .I(\tok.n197 ));
    InMux I__3483 (
            .O(N__20278),
            .I(N__20275));
    LocalMux I__3482 (
            .O(N__20275),
            .I(\tok.n248 ));
    CascadeMux I__3481 (
            .O(N__20272),
            .I(\tok.n6606_cascade_ ));
    InMux I__3480 (
            .O(N__20269),
            .I(N__20266));
    LocalMux I__3479 (
            .O(N__20266),
            .I(\tok.n200 ));
    CascadeMux I__3478 (
            .O(N__20263),
            .I(\tok.n6_cascade_ ));
    InMux I__3477 (
            .O(N__20260),
            .I(N__20253));
    InMux I__3476 (
            .O(N__20259),
            .I(N__20253));
    CascadeMux I__3475 (
            .O(N__20258),
            .I(N__20250));
    LocalMux I__3474 (
            .O(N__20253),
            .I(N__20245));
    InMux I__3473 (
            .O(N__20250),
            .I(N__20242));
    InMux I__3472 (
            .O(N__20249),
            .I(N__20239));
    InMux I__3471 (
            .O(N__20248),
            .I(N__20235));
    Span4Mux_h I__3470 (
            .O(N__20245),
            .I(N__20230));
    LocalMux I__3469 (
            .O(N__20242),
            .I(N__20230));
    LocalMux I__3468 (
            .O(N__20239),
            .I(N__20227));
    InMux I__3467 (
            .O(N__20238),
            .I(N__20223));
    LocalMux I__3466 (
            .O(N__20235),
            .I(N__20216));
    Span4Mux_v I__3465 (
            .O(N__20230),
            .I(N__20216));
    Span4Mux_h I__3464 (
            .O(N__20227),
            .I(N__20216));
    InMux I__3463 (
            .O(N__20226),
            .I(N__20213));
    LocalMux I__3462 (
            .O(N__20223),
            .I(N__20208));
    Span4Mux_v I__3461 (
            .O(N__20216),
            .I(N__20208));
    LocalMux I__3460 (
            .O(N__20213),
            .I(\tok.S_12 ));
    Odrv4 I__3459 (
            .O(N__20208),
            .I(\tok.S_12 ));
    InMux I__3458 (
            .O(N__20203),
            .I(N__20200));
    LocalMux I__3457 (
            .O(N__20200),
            .I(N__20197));
    Odrv12 I__3456 (
            .O(N__20197),
            .I(\tok.n200_adj_875 ));
    CascadeMux I__3455 (
            .O(N__20194),
            .I(\tok.n6_adj_878_cascade_ ));
    InMux I__3454 (
            .O(N__20191),
            .I(N__20187));
    InMux I__3453 (
            .O(N__20190),
            .I(N__20184));
    LocalMux I__3452 (
            .O(N__20187),
            .I(N__20181));
    LocalMux I__3451 (
            .O(N__20184),
            .I(N__20174));
    Span4Mux_v I__3450 (
            .O(N__20181),
            .I(N__20170));
    InMux I__3449 (
            .O(N__20180),
            .I(N__20167));
    InMux I__3448 (
            .O(N__20179),
            .I(N__20164));
    InMux I__3447 (
            .O(N__20178),
            .I(N__20161));
    InMux I__3446 (
            .O(N__20177),
            .I(N__20158));
    Span4Mux_v I__3445 (
            .O(N__20174),
            .I(N__20155));
    CascadeMux I__3444 (
            .O(N__20173),
            .I(N__20152));
    Span4Mux_h I__3443 (
            .O(N__20170),
            .I(N__20145));
    LocalMux I__3442 (
            .O(N__20167),
            .I(N__20145));
    LocalMux I__3441 (
            .O(N__20164),
            .I(N__20145));
    LocalMux I__3440 (
            .O(N__20161),
            .I(N__20142));
    LocalMux I__3439 (
            .O(N__20158),
            .I(N__20139));
    Span4Mux_h I__3438 (
            .O(N__20155),
            .I(N__20136));
    InMux I__3437 (
            .O(N__20152),
            .I(N__20133));
    Span4Mux_h I__3436 (
            .O(N__20145),
            .I(N__20130));
    Span4Mux_s2_v I__3435 (
            .O(N__20142),
            .I(N__20123));
    Span4Mux_v I__3434 (
            .O(N__20139),
            .I(N__20123));
    Span4Mux_v I__3433 (
            .O(N__20136),
            .I(N__20123));
    LocalMux I__3432 (
            .O(N__20133),
            .I(N__20120));
    Span4Mux_v I__3431 (
            .O(N__20130),
            .I(N__20117));
    Odrv4 I__3430 (
            .O(N__20123),
            .I(\tok.S_10 ));
    Odrv12 I__3429 (
            .O(N__20120),
            .I(\tok.S_10 ));
    Odrv4 I__3428 (
            .O(N__20117),
            .I(\tok.S_10 ));
    CascadeMux I__3427 (
            .O(N__20110),
            .I(\tok.n4842_cascade_ ));
    CascadeMux I__3426 (
            .O(N__20107),
            .I(\tok.n7451_cascade_ ));
    InMux I__3425 (
            .O(N__20104),
            .I(N__20101));
    LocalMux I__3424 (
            .O(N__20101),
            .I(N__20098));
    Odrv4 I__3423 (
            .O(N__20098),
            .I(\tok.n6616 ));
    CascadeMux I__3422 (
            .O(N__20095),
            .I(N__20091));
    InMux I__3421 (
            .O(N__20094),
            .I(N__20084));
    InMux I__3420 (
            .O(N__20091),
            .I(N__20081));
    CascadeMux I__3419 (
            .O(N__20090),
            .I(N__20078));
    InMux I__3418 (
            .O(N__20089),
            .I(N__20071));
    InMux I__3417 (
            .O(N__20088),
            .I(N__20071));
    InMux I__3416 (
            .O(N__20087),
            .I(N__20068));
    LocalMux I__3415 (
            .O(N__20084),
            .I(N__20065));
    LocalMux I__3414 (
            .O(N__20081),
            .I(N__20062));
    InMux I__3413 (
            .O(N__20078),
            .I(N__20059));
    InMux I__3412 (
            .O(N__20077),
            .I(N__20056));
    InMux I__3411 (
            .O(N__20076),
            .I(N__20053));
    LocalMux I__3410 (
            .O(N__20071),
            .I(N__20050));
    LocalMux I__3409 (
            .O(N__20068),
            .I(N__20047));
    Span4Mux_v I__3408 (
            .O(N__20065),
            .I(N__20042));
    Span4Mux_v I__3407 (
            .O(N__20062),
            .I(N__20042));
    LocalMux I__3406 (
            .O(N__20059),
            .I(N__20037));
    LocalMux I__3405 (
            .O(N__20056),
            .I(N__20037));
    LocalMux I__3404 (
            .O(N__20053),
            .I(\tok.S_2 ));
    Odrv4 I__3403 (
            .O(N__20050),
            .I(\tok.S_2 ));
    Odrv4 I__3402 (
            .O(N__20047),
            .I(\tok.S_2 ));
    Odrv4 I__3401 (
            .O(N__20042),
            .I(\tok.S_2 ));
    Odrv12 I__3400 (
            .O(N__20037),
            .I(\tok.S_2 ));
    InMux I__3399 (
            .O(N__20026),
            .I(N__20023));
    LocalMux I__3398 (
            .O(N__20023),
            .I(N__20020));
    Odrv4 I__3397 (
            .O(N__20020),
            .I(\tok.n164 ));
    InMux I__3396 (
            .O(N__20017),
            .I(N__20014));
    LocalMux I__3395 (
            .O(N__20014),
            .I(\tok.n6597 ));
    InMux I__3394 (
            .O(N__20011),
            .I(N__20008));
    LocalMux I__3393 (
            .O(N__20008),
            .I(N__20005));
    Span4Mux_v I__3392 (
            .O(N__20005),
            .I(N__20002));
    Odrv4 I__3391 (
            .O(N__20002),
            .I(\tok.n4_adj_711 ));
    CascadeMux I__3390 (
            .O(N__19999),
            .I(N__19996));
    InMux I__3389 (
            .O(N__19996),
            .I(N__19993));
    LocalMux I__3388 (
            .O(N__19993),
            .I(N__19990));
    Odrv12 I__3387 (
            .O(N__19990),
            .I(\tok.n307 ));
    InMux I__3386 (
            .O(N__19987),
            .I(N__19984));
    LocalMux I__3385 (
            .O(N__19984),
            .I(N__19981));
    Odrv12 I__3384 (
            .O(N__19981),
            .I(\tok.n6397 ));
    CascadeMux I__3383 (
            .O(N__19978),
            .I(\tok.n242_cascade_ ));
    CascadeMux I__3382 (
            .O(N__19975),
            .I(N__19972));
    InMux I__3381 (
            .O(N__19972),
            .I(N__19969));
    LocalMux I__3380 (
            .O(N__19969),
            .I(\tok.n6582 ));
    InMux I__3379 (
            .O(N__19966),
            .I(N__19963));
    LocalMux I__3378 (
            .O(N__19963),
            .I(N__19960));
    Span12Mux_s7_v I__3377 (
            .O(N__19960),
            .I(N__19957));
    Odrv12 I__3376 (
            .O(N__19957),
            .I(\tok.table_wr_data_5 ));
    CascadeMux I__3375 (
            .O(N__19954),
            .I(\tok.n199_cascade_ ));
    InMux I__3374 (
            .O(N__19951),
            .I(N__19948));
    LocalMux I__3373 (
            .O(N__19948),
            .I(\tok.n262 ));
    CascadeMux I__3372 (
            .O(N__19945),
            .I(\tok.n4_adj_648_cascade_ ));
    InMux I__3371 (
            .O(N__19942),
            .I(N__19939));
    LocalMux I__3370 (
            .O(N__19939),
            .I(\tok.n326 ));
    InMux I__3369 (
            .O(N__19936),
            .I(N__19932));
    InMux I__3368 (
            .O(N__19935),
            .I(N__19929));
    LocalMux I__3367 (
            .O(N__19932),
            .I(N__19926));
    LocalMux I__3366 (
            .O(N__19929),
            .I(N__19923));
    Span4Mux_v I__3365 (
            .O(N__19926),
            .I(N__19920));
    Span4Mux_v I__3364 (
            .O(N__19923),
            .I(N__19917));
    Span4Mux_h I__3363 (
            .O(N__19920),
            .I(N__19914));
    Span4Mux_h I__3362 (
            .O(N__19917),
            .I(N__19911));
    Odrv4 I__3361 (
            .O(N__19914),
            .I(\tok.n234 ));
    Odrv4 I__3360 (
            .O(N__19911),
            .I(\tok.n234 ));
    CascadeMux I__3359 (
            .O(N__19906),
            .I(N__19902));
    CascadeMux I__3358 (
            .O(N__19905),
            .I(N__19899));
    InMux I__3357 (
            .O(N__19902),
            .I(N__19896));
    InMux I__3356 (
            .O(N__19899),
            .I(N__19893));
    LocalMux I__3355 (
            .O(N__19896),
            .I(N__19890));
    LocalMux I__3354 (
            .O(N__19893),
            .I(N__19887));
    Span4Mux_h I__3353 (
            .O(N__19890),
            .I(N__19884));
    Span12Mux_s10_h I__3352 (
            .O(N__19887),
            .I(N__19881));
    Span4Mux_v I__3351 (
            .O(N__19884),
            .I(N__19878));
    Odrv12 I__3350 (
            .O(N__19881),
            .I(\tok.table_rd_5 ));
    Odrv4 I__3349 (
            .O(N__19878),
            .I(\tok.table_rd_5 ));
    CascadeMux I__3348 (
            .O(N__19873),
            .I(\tok.n286_cascade_ ));
    CascadeMux I__3347 (
            .O(N__19870),
            .I(N__19867));
    InMux I__3346 (
            .O(N__19867),
            .I(N__19864));
    LocalMux I__3345 (
            .O(N__19864),
            .I(N__19861));
    Span4Mux_h I__3344 (
            .O(N__19861),
            .I(N__19857));
    InMux I__3343 (
            .O(N__19860),
            .I(N__19854));
    Odrv4 I__3342 (
            .O(N__19857),
            .I(\tok.n877 ));
    LocalMux I__3341 (
            .O(N__19854),
            .I(\tok.n877 ));
    CascadeMux I__3340 (
            .O(N__19849),
            .I(\tok.n394_cascade_ ));
    CascadeMux I__3339 (
            .O(N__19846),
            .I(N__19843));
    InMux I__3338 (
            .O(N__19843),
            .I(N__19840));
    LocalMux I__3337 (
            .O(N__19840),
            .I(N__19837));
    Span4Mux_h I__3336 (
            .O(N__19837),
            .I(N__19834));
    Odrv4 I__3335 (
            .O(N__19834),
            .I(\tok.n6143 ));
    CascadeMux I__3334 (
            .O(N__19831),
            .I(N__19828));
    InMux I__3333 (
            .O(N__19828),
            .I(N__19825));
    LocalMux I__3332 (
            .O(N__19825),
            .I(N__19822));
    Span4Mux_h I__3331 (
            .O(N__19822),
            .I(N__19819));
    Span4Mux_v I__3330 (
            .O(N__19819),
            .I(N__19816));
    Odrv4 I__3329 (
            .O(N__19816),
            .I(\tok.tc_3 ));
    CascadeMux I__3328 (
            .O(N__19813),
            .I(N__19810));
    InMux I__3327 (
            .O(N__19810),
            .I(N__19807));
    LocalMux I__3326 (
            .O(N__19807),
            .I(N__19804));
    Span4Mux_v I__3325 (
            .O(N__19804),
            .I(N__19801));
    Span4Mux_h I__3324 (
            .O(N__19801),
            .I(N__19798));
    Odrv4 I__3323 (
            .O(N__19798),
            .I(\tok.tc_1 ));
    CascadeMux I__3322 (
            .O(N__19795),
            .I(N__19791));
    InMux I__3321 (
            .O(N__19794),
            .I(N__19788));
    InMux I__3320 (
            .O(N__19791),
            .I(N__19785));
    LocalMux I__3319 (
            .O(N__19788),
            .I(N__19782));
    LocalMux I__3318 (
            .O(N__19785),
            .I(N__19779));
    Span4Mux_s3_v I__3317 (
            .O(N__19782),
            .I(N__19774));
    Span4Mux_v I__3316 (
            .O(N__19779),
            .I(N__19774));
    Odrv4 I__3315 (
            .O(N__19774),
            .I(n92_adj_897));
    CascadeMux I__3314 (
            .O(N__19771),
            .I(N__19768));
    InMux I__3313 (
            .O(N__19768),
            .I(N__19765));
    LocalMux I__3312 (
            .O(N__19765),
            .I(N__19762));
    Span4Mux_v I__3311 (
            .O(N__19762),
            .I(N__19759));
    Span4Mux_h I__3310 (
            .O(N__19759),
            .I(N__19756));
    Odrv4 I__3309 (
            .O(N__19756),
            .I(\tok.tc_0 ));
    InMux I__3308 (
            .O(N__19753),
            .I(N__19739));
    InMux I__3307 (
            .O(N__19752),
            .I(N__19739));
    InMux I__3306 (
            .O(N__19751),
            .I(N__19739));
    InMux I__3305 (
            .O(N__19750),
            .I(N__19739));
    InMux I__3304 (
            .O(N__19749),
            .I(N__19732));
    InMux I__3303 (
            .O(N__19748),
            .I(N__19732));
    LocalMux I__3302 (
            .O(N__19739),
            .I(N__19725));
    InMux I__3301 (
            .O(N__19738),
            .I(N__19720));
    InMux I__3300 (
            .O(N__19737),
            .I(N__19720));
    LocalMux I__3299 (
            .O(N__19732),
            .I(N__19713));
    InMux I__3298 (
            .O(N__19731),
            .I(N__19708));
    InMux I__3297 (
            .O(N__19730),
            .I(N__19708));
    InMux I__3296 (
            .O(N__19729),
            .I(N__19703));
    InMux I__3295 (
            .O(N__19728),
            .I(N__19703));
    Span4Mux_h I__3294 (
            .O(N__19725),
            .I(N__19698));
    LocalMux I__3293 (
            .O(N__19720),
            .I(N__19698));
    InMux I__3292 (
            .O(N__19719),
            .I(N__19689));
    InMux I__3291 (
            .O(N__19718),
            .I(N__19689));
    InMux I__3290 (
            .O(N__19717),
            .I(N__19689));
    InMux I__3289 (
            .O(N__19716),
            .I(N__19689));
    Span4Mux_v I__3288 (
            .O(N__19713),
            .I(N__19686));
    LocalMux I__3287 (
            .O(N__19708),
            .I(N__19681));
    LocalMux I__3286 (
            .O(N__19703),
            .I(N__19681));
    Span4Mux_v I__3285 (
            .O(N__19698),
            .I(N__19676));
    LocalMux I__3284 (
            .O(N__19689),
            .I(N__19676));
    Odrv4 I__3283 (
            .O(N__19686),
            .I(stall_));
    Odrv4 I__3282 (
            .O(N__19681),
            .I(stall_));
    Odrv4 I__3281 (
            .O(N__19676),
            .I(stall_));
    CascadeMux I__3280 (
            .O(N__19669),
            .I(N__19666));
    InMux I__3279 (
            .O(N__19666),
            .I(N__19663));
    LocalMux I__3278 (
            .O(N__19663),
            .I(N__19660));
    Span4Mux_v I__3277 (
            .O(N__19660),
            .I(N__19657));
    Span4Mux_v I__3276 (
            .O(N__19657),
            .I(N__19654));
    Odrv4 I__3275 (
            .O(N__19654),
            .I(\tok.tc_2 ));
    InMux I__3274 (
            .O(N__19651),
            .I(N__19648));
    LocalMux I__3273 (
            .O(N__19648),
            .I(\tok.n6140 ));
    CascadeMux I__3272 (
            .O(N__19645),
            .I(\tok.n225_adj_678_cascade_ ));
    InMux I__3271 (
            .O(N__19642),
            .I(N__19639));
    LocalMux I__3270 (
            .O(N__19639),
            .I(\tok.n6351 ));
    InMux I__3269 (
            .O(N__19636),
            .I(N__19633));
    LocalMux I__3268 (
            .O(N__19633),
            .I(\tok.n6632 ));
    CascadeMux I__3267 (
            .O(N__19630),
            .I(\tok.n7456_cascade_ ));
    CascadeMux I__3266 (
            .O(N__19627),
            .I(N__19624));
    InMux I__3265 (
            .O(N__19624),
            .I(N__19621));
    LocalMux I__3264 (
            .O(N__19621),
            .I(N__19618));
    Span4Mux_v I__3263 (
            .O(N__19618),
            .I(N__19615));
    Span4Mux_h I__3262 (
            .O(N__19615),
            .I(N__19612));
    Odrv4 I__3261 (
            .O(N__19612),
            .I(\tok.n176 ));
    InMux I__3260 (
            .O(N__19609),
            .I(N__19606));
    LocalMux I__3259 (
            .O(N__19606),
            .I(N__19603));
    Odrv12 I__3258 (
            .O(N__19603),
            .I(\tok.n8_adj_686 ));
    InMux I__3257 (
            .O(N__19600),
            .I(N__19597));
    LocalMux I__3256 (
            .O(N__19597),
            .I(\tok.n6622 ));
    CascadeMux I__3255 (
            .O(N__19594),
            .I(\tok.n237_adj_724_cascade_ ));
    InMux I__3254 (
            .O(N__19591),
            .I(N__19588));
    LocalMux I__3253 (
            .O(N__19588),
            .I(N__19585));
    Span4Mux_v I__3252 (
            .O(N__19585),
            .I(N__19582));
    Odrv4 I__3251 (
            .O(N__19582),
            .I(\tok.n4893 ));
    InMux I__3250 (
            .O(N__19579),
            .I(N__19576));
    LocalMux I__3249 (
            .O(N__19576),
            .I(\tok.n286 ));
    CascadeMux I__3248 (
            .O(N__19573),
            .I(\tok.ram.n6260_cascade_ ));
    InMux I__3247 (
            .O(N__19570),
            .I(N__19567));
    LocalMux I__3246 (
            .O(N__19567),
            .I(\tok.n6295 ));
    CascadeMux I__3245 (
            .O(N__19564),
            .I(\tok.n1565_cascade_ ));
    CascadeMux I__3244 (
            .O(N__19561),
            .I(\tok.n13_adj_757_cascade_ ));
    CascadeMux I__3243 (
            .O(N__19558),
            .I(n10_adj_906_cascade_));
    CascadeMux I__3242 (
            .O(N__19555),
            .I(N__19552));
    InMux I__3241 (
            .O(N__19552),
            .I(N__19549));
    LocalMux I__3240 (
            .O(N__19549),
            .I(N__19546));
    Span4Mux_v I__3239 (
            .O(N__19546),
            .I(N__19543));
    Span4Mux_v I__3238 (
            .O(N__19543),
            .I(N__19540));
    Odrv4 I__3237 (
            .O(N__19540),
            .I(\tok.tc_4 ));
    InMux I__3236 (
            .O(N__19537),
            .I(N__19534));
    LocalMux I__3235 (
            .O(N__19534),
            .I(n10_adj_906));
    CascadeMux I__3234 (
            .O(N__19531),
            .I(\tok.n324_cascade_ ));
    InMux I__3233 (
            .O(N__19528),
            .I(N__19525));
    LocalMux I__3232 (
            .O(N__19525),
            .I(\tok.n225_adj_678 ));
    InMux I__3231 (
            .O(N__19522),
            .I(N__19518));
    CascadeMux I__3230 (
            .O(N__19521),
            .I(N__19515));
    LocalMux I__3229 (
            .O(N__19518),
            .I(N__19511));
    InMux I__3228 (
            .O(N__19515),
            .I(N__19508));
    InMux I__3227 (
            .O(N__19514),
            .I(N__19505));
    Span4Mux_h I__3226 (
            .O(N__19511),
            .I(N__19500));
    LocalMux I__3225 (
            .O(N__19508),
            .I(N__19497));
    LocalMux I__3224 (
            .O(N__19505),
            .I(N__19494));
    InMux I__3223 (
            .O(N__19504),
            .I(N__19491));
    CascadeMux I__3222 (
            .O(N__19503),
            .I(N__19488));
    Span4Mux_s0_v I__3221 (
            .O(N__19500),
            .I(N__19482));
    Span4Mux_h I__3220 (
            .O(N__19497),
            .I(N__19482));
    Span4Mux_v I__3219 (
            .O(N__19494),
            .I(N__19477));
    LocalMux I__3218 (
            .O(N__19491),
            .I(N__19477));
    InMux I__3217 (
            .O(N__19488),
            .I(N__19474));
    CascadeMux I__3216 (
            .O(N__19487),
            .I(N__19471));
    Span4Mux_v I__3215 (
            .O(N__19482),
            .I(N__19463));
    Span4Mux_v I__3214 (
            .O(N__19477),
            .I(N__19463));
    LocalMux I__3213 (
            .O(N__19474),
            .I(N__19463));
    InMux I__3212 (
            .O(N__19471),
            .I(N__19460));
    InMux I__3211 (
            .O(N__19470),
            .I(N__19457));
    Span4Mux_h I__3210 (
            .O(N__19463),
            .I(N__19454));
    LocalMux I__3209 (
            .O(N__19460),
            .I(N__19451));
    LocalMux I__3208 (
            .O(N__19457),
            .I(N__19448));
    Span4Mux_s1_h I__3207 (
            .O(N__19454),
            .I(N__19445));
    Span4Mux_h I__3206 (
            .O(N__19451),
            .I(N__19442));
    Odrv4 I__3205 (
            .O(N__19448),
            .I(\tok.S_11 ));
    Odrv4 I__3204 (
            .O(N__19445),
            .I(\tok.S_11 ));
    Odrv4 I__3203 (
            .O(N__19442),
            .I(\tok.S_11 ));
    InMux I__3202 (
            .O(N__19435),
            .I(N__19432));
    LocalMux I__3201 (
            .O(N__19432),
            .I(N__19429));
    Span4Mux_s1_v I__3200 (
            .O(N__19429),
            .I(N__19426));
    Odrv4 I__3199 (
            .O(N__19426),
            .I(\tok.n197_adj_883 ));
    CascadeMux I__3198 (
            .O(N__19423),
            .I(N__19420));
    InMux I__3197 (
            .O(N__19420),
            .I(N__19417));
    LocalMux I__3196 (
            .O(N__19417),
            .I(\tok.n248_adj_884 ));
    CascadeMux I__3195 (
            .O(N__19414),
            .I(\tok.n83_adj_756_cascade_ ));
    InMux I__3194 (
            .O(N__19411),
            .I(N__19408));
    LocalMux I__3193 (
            .O(N__19408),
            .I(N__19405));
    Span4Mux_s2_v I__3192 (
            .O(N__19405),
            .I(N__19402));
    Odrv4 I__3191 (
            .O(N__19402),
            .I(\tok.n248_adj_827 ));
    CascadeMux I__3190 (
            .O(N__19399),
            .I(\tok.n242_adj_828_cascade_ ));
    InMux I__3189 (
            .O(N__19396),
            .I(N__19393));
    LocalMux I__3188 (
            .O(N__19393),
            .I(\tok.n200_adj_829 ));
    InMux I__3187 (
            .O(N__19390),
            .I(N__19384));
    InMux I__3186 (
            .O(N__19389),
            .I(N__19384));
    LocalMux I__3185 (
            .O(N__19384),
            .I(\tok.n231 ));
    InMux I__3184 (
            .O(N__19381),
            .I(N__19378));
    LocalMux I__3183 (
            .O(N__19378),
            .I(N__19375));
    Odrv4 I__3182 (
            .O(N__19375),
            .I(\tok.n242_adj_885 ));
    CascadeMux I__3181 (
            .O(N__19372),
            .I(\tok.n200_adj_886_cascade_ ));
    CascadeMux I__3180 (
            .O(N__19369),
            .I(\tok.n6_adj_889_cascade_ ));
    CascadeMux I__3179 (
            .O(N__19366),
            .I(\tok.n8_cascade_ ));
    InMux I__3178 (
            .O(N__19363),
            .I(N__19360));
    LocalMux I__3177 (
            .O(N__19360),
            .I(N__19357));
    Odrv12 I__3176 (
            .O(N__19357),
            .I(\tok.n6368 ));
    InMux I__3175 (
            .O(N__19354),
            .I(N__19351));
    LocalMux I__3174 (
            .O(N__19351),
            .I(\tok.n197_adj_668 ));
    CascadeMux I__3173 (
            .O(N__19348),
            .I(\tok.n248_adj_669_cascade_ ));
    InMux I__3172 (
            .O(N__19345),
            .I(N__19342));
    LocalMux I__3171 (
            .O(N__19342),
            .I(\tok.n242_adj_670 ));
    CascadeMux I__3170 (
            .O(N__19339),
            .I(\tok.n200_adj_671_cascade_ ));
    CascadeMux I__3169 (
            .O(N__19336),
            .I(N__19330));
    InMux I__3168 (
            .O(N__19335),
            .I(N__19325));
    InMux I__3167 (
            .O(N__19334),
            .I(N__19325));
    InMux I__3166 (
            .O(N__19333),
            .I(N__19322));
    InMux I__3165 (
            .O(N__19330),
            .I(N__19317));
    LocalMux I__3164 (
            .O(N__19325),
            .I(N__19314));
    LocalMux I__3163 (
            .O(N__19322),
            .I(N__19311));
    InMux I__3162 (
            .O(N__19321),
            .I(N__19308));
    InMux I__3161 (
            .O(N__19320),
            .I(N__19305));
    LocalMux I__3160 (
            .O(N__19317),
            .I(N__19301));
    Span4Mux_v I__3159 (
            .O(N__19314),
            .I(N__19292));
    Span4Mux_v I__3158 (
            .O(N__19311),
            .I(N__19292));
    LocalMux I__3157 (
            .O(N__19308),
            .I(N__19292));
    LocalMux I__3156 (
            .O(N__19305),
            .I(N__19292));
    InMux I__3155 (
            .O(N__19304),
            .I(N__19289));
    Span4Mux_v I__3154 (
            .O(N__19301),
            .I(N__19286));
    Span4Mux_v I__3153 (
            .O(N__19292),
            .I(N__19283));
    LocalMux I__3152 (
            .O(N__19289),
            .I(N__19278));
    Span4Mux_v I__3151 (
            .O(N__19286),
            .I(N__19278));
    Span4Mux_h I__3150 (
            .O(N__19283),
            .I(N__19275));
    Odrv4 I__3149 (
            .O(N__19278),
            .I(\tok.S_14 ));
    Odrv4 I__3148 (
            .O(N__19275),
            .I(\tok.S_14 ));
    CascadeMux I__3147 (
            .O(N__19270),
            .I(\tok.n6_adj_674_cascade_ ));
    CascadeMux I__3146 (
            .O(N__19267),
            .I(N__19264));
    InMux I__3145 (
            .O(N__19264),
            .I(N__19261));
    LocalMux I__3144 (
            .O(N__19261),
            .I(N__19258));
    Span4Mux_v I__3143 (
            .O(N__19258),
            .I(N__19255));
    Odrv4 I__3142 (
            .O(N__19255),
            .I(\tok.table_rd_8 ));
    CascadeMux I__3141 (
            .O(N__19252),
            .I(N__19248));
    CascadeMux I__3140 (
            .O(N__19251),
            .I(N__19241));
    InMux I__3139 (
            .O(N__19248),
            .I(N__19237));
    InMux I__3138 (
            .O(N__19247),
            .I(N__19234));
    InMux I__3137 (
            .O(N__19246),
            .I(N__19231));
    InMux I__3136 (
            .O(N__19245),
            .I(N__19228));
    InMux I__3135 (
            .O(N__19244),
            .I(N__19225));
    InMux I__3134 (
            .O(N__19241),
            .I(N__19222));
    InMux I__3133 (
            .O(N__19240),
            .I(N__19219));
    LocalMux I__3132 (
            .O(N__19237),
            .I(N__19215));
    LocalMux I__3131 (
            .O(N__19234),
            .I(N__19209));
    LocalMux I__3130 (
            .O(N__19231),
            .I(N__19209));
    LocalMux I__3129 (
            .O(N__19228),
            .I(N__19206));
    LocalMux I__3128 (
            .O(N__19225),
            .I(N__19199));
    LocalMux I__3127 (
            .O(N__19222),
            .I(N__19199));
    LocalMux I__3126 (
            .O(N__19219),
            .I(N__19199));
    InMux I__3125 (
            .O(N__19218),
            .I(N__19196));
    Span4Mux_v I__3124 (
            .O(N__19215),
            .I(N__19193));
    InMux I__3123 (
            .O(N__19214),
            .I(N__19190));
    Span4Mux_v I__3122 (
            .O(N__19209),
            .I(N__19187));
    Span4Mux_s2_v I__3121 (
            .O(N__19206),
            .I(N__19180));
    Span4Mux_v I__3120 (
            .O(N__19199),
            .I(N__19180));
    LocalMux I__3119 (
            .O(N__19196),
            .I(N__19180));
    Span4Mux_v I__3118 (
            .O(N__19193),
            .I(N__19177));
    LocalMux I__3117 (
            .O(N__19190),
            .I(\tok.n7269 ));
    Odrv4 I__3116 (
            .O(N__19187),
            .I(\tok.n7269 ));
    Odrv4 I__3115 (
            .O(N__19180),
            .I(\tok.n7269 ));
    Odrv4 I__3114 (
            .O(N__19177),
            .I(\tok.n7269 ));
    CascadeMux I__3113 (
            .O(N__19168),
            .I(\tok.n203_adj_822_cascade_ ));
    CascadeMux I__3112 (
            .O(N__19165),
            .I(\tok.n212_adj_824_cascade_ ));
    CascadeMux I__3111 (
            .O(N__19162),
            .I(\tok.n6457_cascade_ ));
    InMux I__3110 (
            .O(N__19159),
            .I(N__19156));
    LocalMux I__3109 (
            .O(N__19156),
            .I(N__19153));
    Odrv12 I__3108 (
            .O(N__19153),
            .I(\tok.n208_adj_857 ));
    CascadeMux I__3107 (
            .O(N__19150),
            .I(N__19147));
    InMux I__3106 (
            .O(N__19147),
            .I(N__19144));
    LocalMux I__3105 (
            .O(N__19144),
            .I(\tok.n6328 ));
    CascadeMux I__3104 (
            .O(N__19141),
            .I(N__19138));
    InMux I__3103 (
            .O(N__19138),
            .I(N__19135));
    LocalMux I__3102 (
            .O(N__19135),
            .I(N__19132));
    Odrv12 I__3101 (
            .O(N__19132),
            .I(\tok.n250 ));
    CascadeMux I__3100 (
            .O(N__19129),
            .I(\tok.n190_adj_774_cascade_ ));
    InMux I__3099 (
            .O(N__19126),
            .I(N__19123));
    LocalMux I__3098 (
            .O(N__19123),
            .I(N__19120));
    Span4Mux_h I__3097 (
            .O(N__19120),
            .I(N__19117));
    Odrv4 I__3096 (
            .O(N__19117),
            .I(\tok.n6514 ));
    CascadeMux I__3095 (
            .O(N__19114),
            .I(\tok.n833_cascade_ ));
    InMux I__3094 (
            .O(N__19111),
            .I(N__19108));
    LocalMux I__3093 (
            .O(N__19108),
            .I(N__19105));
    Odrv4 I__3092 (
            .O(N__19105),
            .I(\tok.n6515 ));
    CascadeMux I__3091 (
            .O(N__19102),
            .I(\tok.n6534_cascade_ ));
    CascadeMux I__3090 (
            .O(N__19099),
            .I(\tok.n252_adj_783_cascade_ ));
    InMux I__3089 (
            .O(N__19096),
            .I(N__19093));
    LocalMux I__3088 (
            .O(N__19093),
            .I(\tok.n255_adj_775 ));
    CascadeMux I__3087 (
            .O(N__19090),
            .I(N__19087));
    InMux I__3086 (
            .O(N__19087),
            .I(N__19084));
    LocalMux I__3085 (
            .O(N__19084),
            .I(\tok.n190_adj_774 ));
    InMux I__3084 (
            .O(N__19081),
            .I(N__19078));
    LocalMux I__3083 (
            .O(N__19078),
            .I(\tok.n258_adj_780 ));
    InMux I__3082 (
            .O(N__19075),
            .I(N__19072));
    LocalMux I__3081 (
            .O(N__19072),
            .I(\tok.n177_adj_779 ));
    InMux I__3080 (
            .O(N__19069),
            .I(N__19066));
    LocalMux I__3079 (
            .O(N__19066),
            .I(\tok.n22_adj_847 ));
    InMux I__3078 (
            .O(N__19063),
            .I(N__19060));
    LocalMux I__3077 (
            .O(N__19060),
            .I(\tok.n27_adj_782 ));
    InMux I__3076 (
            .O(N__19057),
            .I(N__19054));
    LocalMux I__3075 (
            .O(N__19054),
            .I(\tok.n298 ));
    InMux I__3074 (
            .O(N__19051),
            .I(N__19048));
    LocalMux I__3073 (
            .O(N__19048),
            .I(\tok.n161_adj_870 ));
    CascadeMux I__3072 (
            .O(N__19045),
            .I(\tok.n6429_cascade_ ));
    CascadeMux I__3071 (
            .O(N__19042),
            .I(\tok.n197_adj_872_cascade_ ));
    CascadeMux I__3070 (
            .O(N__19039),
            .I(N__19036));
    InMux I__3069 (
            .O(N__19036),
            .I(N__19033));
    LocalMux I__3068 (
            .O(N__19033),
            .I(N__19030));
    Span4Mux_s3_h I__3067 (
            .O(N__19030),
            .I(N__19027));
    Odrv4 I__3066 (
            .O(N__19027),
            .I(\tok.n248_adj_873 ));
    InMux I__3065 (
            .O(N__19024),
            .I(N__19021));
    LocalMux I__3064 (
            .O(N__19021),
            .I(\tok.n296 ));
    CascadeMux I__3063 (
            .O(N__19018),
            .I(\tok.n6400_cascade_ ));
    InMux I__3062 (
            .O(N__19015),
            .I(N__19012));
    LocalMux I__3061 (
            .O(N__19012),
            .I(\tok.n161 ));
    CascadeMux I__3060 (
            .O(N__19009),
            .I(N__19006));
    InMux I__3059 (
            .O(N__19006),
            .I(N__19003));
    LocalMux I__3058 (
            .O(N__19003),
            .I(N__19000));
    Odrv4 I__3057 (
            .O(N__19000),
            .I(\tok.n6406 ));
    InMux I__3056 (
            .O(N__18997),
            .I(N__18994));
    LocalMux I__3055 (
            .O(N__18994),
            .I(\tok.n6415 ));
    CascadeMux I__3054 (
            .O(N__18991),
            .I(\tok.n161_adj_882_cascade_ ));
    InMux I__3053 (
            .O(N__18988),
            .I(N__18985));
    LocalMux I__3052 (
            .O(N__18985),
            .I(\tok.n26_adj_781 ));
    CascadeMux I__3051 (
            .O(N__18982),
            .I(\tok.n28_adj_778_cascade_ ));
    InMux I__3050 (
            .O(N__18979),
            .I(N__18976));
    LocalMux I__3049 (
            .O(N__18976),
            .I(\tok.n25_adj_788 ));
    CascadeMux I__3048 (
            .O(N__18973),
            .I(N__18969));
    InMux I__3047 (
            .O(N__18972),
            .I(N__18964));
    InMux I__3046 (
            .O(N__18969),
            .I(N__18964));
    LocalMux I__3045 (
            .O(N__18964),
            .I(N__18959));
    InMux I__3044 (
            .O(N__18963),
            .I(N__18956));
    InMux I__3043 (
            .O(N__18962),
            .I(N__18952));
    Span4Mux_s3_v I__3042 (
            .O(N__18959),
            .I(N__18945));
    LocalMux I__3041 (
            .O(N__18956),
            .I(N__18945));
    InMux I__3040 (
            .O(N__18955),
            .I(N__18942));
    LocalMux I__3039 (
            .O(N__18952),
            .I(N__18939));
    InMux I__3038 (
            .O(N__18951),
            .I(N__18936));
    InMux I__3037 (
            .O(N__18950),
            .I(N__18933));
    Sp12to4 I__3036 (
            .O(N__18945),
            .I(N__18928));
    LocalMux I__3035 (
            .O(N__18942),
            .I(N__18928));
    Span4Mux_s3_v I__3034 (
            .O(N__18939),
            .I(N__18923));
    LocalMux I__3033 (
            .O(N__18936),
            .I(N__18923));
    LocalMux I__3032 (
            .O(N__18933),
            .I(N__18920));
    Span12Mux_s6_v I__3031 (
            .O(N__18928),
            .I(N__18917));
    Span4Mux_v I__3030 (
            .O(N__18923),
            .I(N__18912));
    Span4Mux_h I__3029 (
            .O(N__18920),
            .I(N__18912));
    Odrv12 I__3028 (
            .O(N__18917),
            .I(\tok.S_15 ));
    Odrv4 I__3027 (
            .O(N__18912),
            .I(\tok.S_15 ));
    InMux I__3026 (
            .O(N__18907),
            .I(N__18904));
    LocalMux I__3025 (
            .O(N__18904),
            .I(\tok.n6634 ));
    InMux I__3024 (
            .O(N__18901),
            .I(N__18898));
    LocalMux I__3023 (
            .O(N__18898),
            .I(\tok.n23_adj_848 ));
    CascadeMux I__3022 (
            .O(N__18895),
            .I(\tok.n21_adj_849_cascade_ ));
    InMux I__3021 (
            .O(N__18892),
            .I(N__18889));
    LocalMux I__3020 (
            .O(N__18889),
            .I(\tok.n24_adj_846 ));
    CascadeMux I__3019 (
            .O(N__18886),
            .I(N__18883));
    InMux I__3018 (
            .O(N__18883),
            .I(N__18880));
    LocalMux I__3017 (
            .O(N__18880),
            .I(N__18877));
    Odrv4 I__3016 (
            .O(N__18877),
            .I(\tok.n30_adj_852 ));
    CascadeMux I__3015 (
            .O(N__18874),
            .I(N__18871));
    InMux I__3014 (
            .O(N__18871),
            .I(N__18868));
    LocalMux I__3013 (
            .O(N__18868),
            .I(\tok.n323 ));
    InMux I__3012 (
            .O(N__18865),
            .I(N__18862));
    LocalMux I__3011 (
            .O(N__18862),
            .I(\tok.n163 ));
    InMux I__3010 (
            .O(N__18859),
            .I(N__18856));
    LocalMux I__3009 (
            .O(N__18856),
            .I(\tok.n256_adj_862 ));
    InMux I__3008 (
            .O(N__18853),
            .I(N__18850));
    LocalMux I__3007 (
            .O(N__18850),
            .I(N__18847));
    Span4Mux_v I__3006 (
            .O(N__18847),
            .I(N__18844));
    Span4Mux_h I__3005 (
            .O(N__18844),
            .I(N__18841));
    Odrv4 I__3004 (
            .O(N__18841),
            .I(\tok.n5_adj_871 ));
    CascadeMux I__3003 (
            .O(N__18838),
            .I(\tok.n6_adj_868_cascade_ ));
    InMux I__3002 (
            .O(N__18835),
            .I(N__18829));
    InMux I__3001 (
            .O(N__18834),
            .I(N__18823));
    InMux I__3000 (
            .O(N__18833),
            .I(N__18823));
    CascadeMux I__2999 (
            .O(N__18832),
            .I(N__18820));
    LocalMux I__2998 (
            .O(N__18829),
            .I(N__18817));
    InMux I__2997 (
            .O(N__18828),
            .I(N__18814));
    LocalMux I__2996 (
            .O(N__18823),
            .I(N__18809));
    InMux I__2995 (
            .O(N__18820),
            .I(N__18806));
    Span4Mux_v I__2994 (
            .O(N__18817),
            .I(N__18801));
    LocalMux I__2993 (
            .O(N__18814),
            .I(N__18801));
    InMux I__2992 (
            .O(N__18813),
            .I(N__18798));
    InMux I__2991 (
            .O(N__18812),
            .I(N__18795));
    Span4Mux_v I__2990 (
            .O(N__18809),
            .I(N__18792));
    LocalMux I__2989 (
            .O(N__18806),
            .I(N__18789));
    Span4Mux_v I__2988 (
            .O(N__18801),
            .I(N__18786));
    LocalMux I__2987 (
            .O(N__18798),
            .I(N__18783));
    LocalMux I__2986 (
            .O(N__18795),
            .I(N__18776));
    Span4Mux_h I__2985 (
            .O(N__18792),
            .I(N__18776));
    Span4Mux_h I__2984 (
            .O(N__18789),
            .I(N__18776));
    Span4Mux_h I__2983 (
            .O(N__18786),
            .I(N__18773));
    Odrv12 I__2982 (
            .O(N__18783),
            .I(S_0));
    Odrv4 I__2981 (
            .O(N__18776),
            .I(S_0));
    Odrv4 I__2980 (
            .O(N__18773),
            .I(S_0));
    InMux I__2979 (
            .O(N__18766),
            .I(N__18763));
    LocalMux I__2978 (
            .O(N__18763),
            .I(N__18760));
    Span4Mux_h I__2977 (
            .O(N__18760),
            .I(N__18757));
    Odrv4 I__2976 (
            .O(N__18757),
            .I(\tok.n28 ));
    CascadeMux I__2975 (
            .O(N__18754),
            .I(N__18750));
    InMux I__2974 (
            .O(N__18753),
            .I(N__18745));
    InMux I__2973 (
            .O(N__18750),
            .I(N__18745));
    LocalMux I__2972 (
            .O(N__18745),
            .I(N__18742));
    Span4Mux_v I__2971 (
            .O(N__18742),
            .I(N__18739));
    Span4Mux_h I__2970 (
            .O(N__18739),
            .I(N__18736));
    Odrv4 I__2969 (
            .O(N__18736),
            .I(\tok.key_rd_11 ));
    CascadeMux I__2968 (
            .O(N__18733),
            .I(N__18730));
    InMux I__2967 (
            .O(N__18730),
            .I(N__18724));
    InMux I__2966 (
            .O(N__18729),
            .I(N__18724));
    LocalMux I__2965 (
            .O(N__18724),
            .I(N__18721));
    Span4Mux_h I__2964 (
            .O(N__18721),
            .I(N__18718));
    Odrv4 I__2963 (
            .O(N__18718),
            .I(\tok.key_rd_14 ));
    InMux I__2962 (
            .O(N__18715),
            .I(N__18712));
    LocalMux I__2961 (
            .O(N__18712),
            .I(N__18709));
    Odrv12 I__2960 (
            .O(N__18709),
            .I(\tok.n23_adj_638 ));
    CascadeMux I__2959 (
            .O(N__18706),
            .I(N__18702));
    InMux I__2958 (
            .O(N__18705),
            .I(N__18697));
    InMux I__2957 (
            .O(N__18702),
            .I(N__18697));
    LocalMux I__2956 (
            .O(N__18697),
            .I(N__18694));
    Span4Mux_v I__2955 (
            .O(N__18694),
            .I(N__18691));
    Odrv4 I__2954 (
            .O(N__18691),
            .I(\tok.key_rd_15 ));
    InMux I__2953 (
            .O(N__18688),
            .I(N__18682));
    InMux I__2952 (
            .O(N__18687),
            .I(N__18682));
    LocalMux I__2951 (
            .O(N__18682),
            .I(N__18679));
    Span4Mux_h I__2950 (
            .O(N__18679),
            .I(N__18676));
    Odrv4 I__2949 (
            .O(N__18676),
            .I(\tok.key_rd_9 ));
    InMux I__2948 (
            .O(N__18673),
            .I(N__18670));
    LocalMux I__2947 (
            .O(N__18670),
            .I(N__18667));
    Odrv12 I__2946 (
            .O(N__18667),
            .I(\tok.n24 ));
    CascadeMux I__2945 (
            .O(N__18664),
            .I(\tok.n283_cascade_ ));
    CascadeMux I__2944 (
            .O(N__18661),
            .I(\tok.n223_cascade_ ));
    InMux I__2943 (
            .O(N__18658),
            .I(N__18655));
    LocalMux I__2942 (
            .O(N__18655),
            .I(\tok.n4_adj_752 ));
    CascadeMux I__2941 (
            .O(N__18652),
            .I(\tok.n6586_cascade_ ));
    InMux I__2940 (
            .O(N__18649),
            .I(N__18646));
    LocalMux I__2939 (
            .O(N__18646),
            .I(\tok.n226_adj_744 ));
    InMux I__2938 (
            .O(N__18643),
            .I(N__18640));
    LocalMux I__2937 (
            .O(N__18640),
            .I(\tok.n254 ));
    InMux I__2936 (
            .O(N__18637),
            .I(N__18634));
    LocalMux I__2935 (
            .O(N__18634),
            .I(N__18631));
    Odrv4 I__2934 (
            .O(N__18631),
            .I(\tok.n319 ));
    InMux I__2933 (
            .O(N__18628),
            .I(N__18625));
    LocalMux I__2932 (
            .O(N__18625),
            .I(N__18622));
    Span4Mux_h I__2931 (
            .O(N__18622),
            .I(N__18619));
    Odrv4 I__2930 (
            .O(N__18619),
            .I(\tok.n6326 ));
    CascadeMux I__2929 (
            .O(N__18616),
            .I(\tok.n387_cascade_ ));
    CascadeMux I__2928 (
            .O(N__18613),
            .I(\tok.n254_adj_860_cascade_ ));
    CascadeMux I__2927 (
            .O(N__18610),
            .I(N__18607));
    InMux I__2926 (
            .O(N__18607),
            .I(N__18603));
    InMux I__2925 (
            .O(N__18606),
            .I(N__18600));
    LocalMux I__2924 (
            .O(N__18603),
            .I(N__18597));
    LocalMux I__2923 (
            .O(N__18600),
            .I(\tok.n5_adj_675 ));
    Odrv4 I__2922 (
            .O(N__18597),
            .I(\tok.n5_adj_675 ));
    CascadeMux I__2921 (
            .O(N__18592),
            .I(\tok.n6205_cascade_ ));
    InMux I__2920 (
            .O(N__18589),
            .I(N__18578));
    InMux I__2919 (
            .O(N__18588),
            .I(N__18573));
    InMux I__2918 (
            .O(N__18587),
            .I(N__18573));
    InMux I__2917 (
            .O(N__18586),
            .I(N__18570));
    InMux I__2916 (
            .O(N__18585),
            .I(N__18566));
    InMux I__2915 (
            .O(N__18584),
            .I(N__18559));
    InMux I__2914 (
            .O(N__18583),
            .I(N__18556));
    InMux I__2913 (
            .O(N__18582),
            .I(N__18551));
    InMux I__2912 (
            .O(N__18581),
            .I(N__18551));
    LocalMux I__2911 (
            .O(N__18578),
            .I(N__18543));
    LocalMux I__2910 (
            .O(N__18573),
            .I(N__18543));
    LocalMux I__2909 (
            .O(N__18570),
            .I(N__18543));
    InMux I__2908 (
            .O(N__18569),
            .I(N__18540));
    LocalMux I__2907 (
            .O(N__18566),
            .I(N__18537));
    InMux I__2906 (
            .O(N__18565),
            .I(N__18530));
    InMux I__2905 (
            .O(N__18564),
            .I(N__18530));
    InMux I__2904 (
            .O(N__18563),
            .I(N__18530));
    InMux I__2903 (
            .O(N__18562),
            .I(N__18527));
    LocalMux I__2902 (
            .O(N__18559),
            .I(N__18524));
    LocalMux I__2901 (
            .O(N__18556),
            .I(N__18519));
    LocalMux I__2900 (
            .O(N__18551),
            .I(N__18519));
    InMux I__2899 (
            .O(N__18550),
            .I(N__18516));
    Span4Mux_v I__2898 (
            .O(N__18543),
            .I(N__18511));
    LocalMux I__2897 (
            .O(N__18540),
            .I(N__18511));
    Span4Mux_s0_v I__2896 (
            .O(N__18537),
            .I(N__18506));
    LocalMux I__2895 (
            .O(N__18530),
            .I(N__18506));
    LocalMux I__2894 (
            .O(N__18527),
            .I(N__18503));
    Span4Mux_s3_v I__2893 (
            .O(N__18524),
            .I(N__18496));
    Span4Mux_v I__2892 (
            .O(N__18519),
            .I(N__18496));
    LocalMux I__2891 (
            .O(N__18516),
            .I(N__18496));
    Span4Mux_h I__2890 (
            .O(N__18511),
            .I(N__18491));
    Span4Mux_v I__2889 (
            .O(N__18506),
            .I(N__18491));
    Span4Mux_s3_v I__2888 (
            .O(N__18503),
            .I(N__18486));
    Span4Mux_h I__2887 (
            .O(N__18496),
            .I(N__18486));
    Odrv4 I__2886 (
            .O(N__18491),
            .I(\tok.n270 ));
    Odrv4 I__2885 (
            .O(N__18486),
            .I(\tok.n270 ));
    CascadeMux I__2884 (
            .O(N__18481),
            .I(\tok.n270_cascade_ ));
    InMux I__2883 (
            .O(N__18478),
            .I(N__18475));
    LocalMux I__2882 (
            .O(N__18475),
            .I(N__18472));
    Span4Mux_v I__2881 (
            .O(N__18472),
            .I(N__18469));
    Span4Mux_h I__2880 (
            .O(N__18469),
            .I(N__18465));
    InMux I__2879 (
            .O(N__18468),
            .I(N__18462));
    Odrv4 I__2878 (
            .O(N__18465),
            .I(\tok.A_stk.tail_18 ));
    LocalMux I__2877 (
            .O(N__18462),
            .I(\tok.A_stk.tail_18 ));
    InMux I__2876 (
            .O(N__18457),
            .I(N__18424));
    InMux I__2875 (
            .O(N__18456),
            .I(N__18424));
    InMux I__2874 (
            .O(N__18455),
            .I(N__18424));
    InMux I__2873 (
            .O(N__18454),
            .I(N__18424));
    InMux I__2872 (
            .O(N__18453),
            .I(N__18424));
    InMux I__2871 (
            .O(N__18452),
            .I(N__18424));
    InMux I__2870 (
            .O(N__18451),
            .I(N__18424));
    InMux I__2869 (
            .O(N__18450),
            .I(N__18409));
    InMux I__2868 (
            .O(N__18449),
            .I(N__18409));
    InMux I__2867 (
            .O(N__18448),
            .I(N__18409));
    InMux I__2866 (
            .O(N__18447),
            .I(N__18409));
    InMux I__2865 (
            .O(N__18446),
            .I(N__18409));
    InMux I__2864 (
            .O(N__18445),
            .I(N__18409));
    InMux I__2863 (
            .O(N__18444),
            .I(N__18409));
    InMux I__2862 (
            .O(N__18443),
            .I(N__18398));
    InMux I__2861 (
            .O(N__18442),
            .I(N__18398));
    InMux I__2860 (
            .O(N__18441),
            .I(N__18398));
    InMux I__2859 (
            .O(N__18440),
            .I(N__18398));
    InMux I__2858 (
            .O(N__18439),
            .I(N__18398));
    LocalMux I__2857 (
            .O(N__18424),
            .I(N__18338));
    LocalMux I__2856 (
            .O(N__18409),
            .I(N__18338));
    LocalMux I__2855 (
            .O(N__18398),
            .I(N__18338));
    InMux I__2854 (
            .O(N__18397),
            .I(N__18323));
    InMux I__2853 (
            .O(N__18396),
            .I(N__18323));
    InMux I__2852 (
            .O(N__18395),
            .I(N__18323));
    InMux I__2851 (
            .O(N__18394),
            .I(N__18323));
    InMux I__2850 (
            .O(N__18393),
            .I(N__18323));
    InMux I__2849 (
            .O(N__18392),
            .I(N__18323));
    InMux I__2848 (
            .O(N__18391),
            .I(N__18323));
    InMux I__2847 (
            .O(N__18390),
            .I(N__18299));
    InMux I__2846 (
            .O(N__18389),
            .I(N__18299));
    InMux I__2845 (
            .O(N__18388),
            .I(N__18299));
    InMux I__2844 (
            .O(N__18387),
            .I(N__18299));
    InMux I__2843 (
            .O(N__18386),
            .I(N__18299));
    InMux I__2842 (
            .O(N__18385),
            .I(N__18299));
    InMux I__2841 (
            .O(N__18384),
            .I(N__18299));
    InMux I__2840 (
            .O(N__18383),
            .I(N__18299));
    InMux I__2839 (
            .O(N__18382),
            .I(N__18282));
    InMux I__2838 (
            .O(N__18381),
            .I(N__18282));
    InMux I__2837 (
            .O(N__18380),
            .I(N__18282));
    InMux I__2836 (
            .O(N__18379),
            .I(N__18282));
    InMux I__2835 (
            .O(N__18378),
            .I(N__18282));
    InMux I__2834 (
            .O(N__18377),
            .I(N__18282));
    InMux I__2833 (
            .O(N__18376),
            .I(N__18282));
    InMux I__2832 (
            .O(N__18375),
            .I(N__18282));
    InMux I__2831 (
            .O(N__18374),
            .I(N__18277));
    InMux I__2830 (
            .O(N__18373),
            .I(N__18277));
    InMux I__2829 (
            .O(N__18372),
            .I(N__18260));
    InMux I__2828 (
            .O(N__18371),
            .I(N__18260));
    InMux I__2827 (
            .O(N__18370),
            .I(N__18260));
    InMux I__2826 (
            .O(N__18369),
            .I(N__18260));
    InMux I__2825 (
            .O(N__18368),
            .I(N__18260));
    InMux I__2824 (
            .O(N__18367),
            .I(N__18260));
    InMux I__2823 (
            .O(N__18366),
            .I(N__18260));
    InMux I__2822 (
            .O(N__18365),
            .I(N__18260));
    InMux I__2821 (
            .O(N__18364),
            .I(N__18255));
    InMux I__2820 (
            .O(N__18363),
            .I(N__18255));
    InMux I__2819 (
            .O(N__18362),
            .I(N__18238));
    InMux I__2818 (
            .O(N__18361),
            .I(N__18238));
    InMux I__2817 (
            .O(N__18360),
            .I(N__18238));
    InMux I__2816 (
            .O(N__18359),
            .I(N__18238));
    InMux I__2815 (
            .O(N__18358),
            .I(N__18238));
    InMux I__2814 (
            .O(N__18357),
            .I(N__18238));
    InMux I__2813 (
            .O(N__18356),
            .I(N__18238));
    InMux I__2812 (
            .O(N__18355),
            .I(N__18223));
    InMux I__2811 (
            .O(N__18354),
            .I(N__18223));
    InMux I__2810 (
            .O(N__18353),
            .I(N__18223));
    InMux I__2809 (
            .O(N__18352),
            .I(N__18223));
    InMux I__2808 (
            .O(N__18351),
            .I(N__18223));
    InMux I__2807 (
            .O(N__18350),
            .I(N__18223));
    InMux I__2806 (
            .O(N__18349),
            .I(N__18223));
    InMux I__2805 (
            .O(N__18348),
            .I(N__18220));
    InMux I__2804 (
            .O(N__18347),
            .I(N__18209));
    InMux I__2803 (
            .O(N__18346),
            .I(N__18209));
    InMux I__2802 (
            .O(N__18345),
            .I(N__18209));
    Span4Mux_s3_v I__2801 (
            .O(N__18338),
            .I(N__18204));
    LocalMux I__2800 (
            .O(N__18323),
            .I(N__18204));
    InMux I__2799 (
            .O(N__18322),
            .I(N__18152));
    InMux I__2798 (
            .O(N__18321),
            .I(N__18152));
    InMux I__2797 (
            .O(N__18320),
            .I(N__18152));
    InMux I__2796 (
            .O(N__18319),
            .I(N__18152));
    InMux I__2795 (
            .O(N__18318),
            .I(N__18152));
    InMux I__2794 (
            .O(N__18317),
            .I(N__18152));
    InMux I__2793 (
            .O(N__18316),
            .I(N__18152));
    LocalMux I__2792 (
            .O(N__18299),
            .I(N__18145));
    LocalMux I__2791 (
            .O(N__18282),
            .I(N__18145));
    LocalMux I__2790 (
            .O(N__18277),
            .I(N__18145));
    LocalMux I__2789 (
            .O(N__18260),
            .I(N__18140));
    LocalMux I__2788 (
            .O(N__18255),
            .I(N__18140));
    InMux I__2787 (
            .O(N__18254),
            .I(N__18137));
    InMux I__2786 (
            .O(N__18253),
            .I(N__18134));
    LocalMux I__2785 (
            .O(N__18238),
            .I(N__18127));
    LocalMux I__2784 (
            .O(N__18223),
            .I(N__18127));
    LocalMux I__2783 (
            .O(N__18220),
            .I(N__18127));
    InMux I__2782 (
            .O(N__18219),
            .I(N__18118));
    InMux I__2781 (
            .O(N__18218),
            .I(N__18118));
    InMux I__2780 (
            .O(N__18217),
            .I(N__18118));
    InMux I__2779 (
            .O(N__18216),
            .I(N__18118));
    LocalMux I__2778 (
            .O(N__18209),
            .I(N__18108));
    Span4Mux_h I__2777 (
            .O(N__18204),
            .I(N__18108));
    InMux I__2776 (
            .O(N__18203),
            .I(N__18101));
    InMux I__2775 (
            .O(N__18202),
            .I(N__18101));
    InMux I__2774 (
            .O(N__18201),
            .I(N__18101));
    InMux I__2773 (
            .O(N__18200),
            .I(N__18088));
    InMux I__2772 (
            .O(N__18199),
            .I(N__18088));
    InMux I__2771 (
            .O(N__18198),
            .I(N__18088));
    InMux I__2770 (
            .O(N__18197),
            .I(N__18088));
    InMux I__2769 (
            .O(N__18196),
            .I(N__18088));
    InMux I__2768 (
            .O(N__18195),
            .I(N__18088));
    InMux I__2767 (
            .O(N__18194),
            .I(N__18073));
    InMux I__2766 (
            .O(N__18193),
            .I(N__18073));
    InMux I__2765 (
            .O(N__18192),
            .I(N__18073));
    InMux I__2764 (
            .O(N__18191),
            .I(N__18073));
    InMux I__2763 (
            .O(N__18190),
            .I(N__18073));
    InMux I__2762 (
            .O(N__18189),
            .I(N__18073));
    InMux I__2761 (
            .O(N__18188),
            .I(N__18073));
    InMux I__2760 (
            .O(N__18187),
            .I(N__18058));
    InMux I__2759 (
            .O(N__18186),
            .I(N__18058));
    InMux I__2758 (
            .O(N__18185),
            .I(N__18058));
    InMux I__2757 (
            .O(N__18184),
            .I(N__18058));
    InMux I__2756 (
            .O(N__18183),
            .I(N__18058));
    InMux I__2755 (
            .O(N__18182),
            .I(N__18058));
    InMux I__2754 (
            .O(N__18181),
            .I(N__18058));
    InMux I__2753 (
            .O(N__18180),
            .I(N__18045));
    InMux I__2752 (
            .O(N__18179),
            .I(N__18045));
    InMux I__2751 (
            .O(N__18178),
            .I(N__18045));
    InMux I__2750 (
            .O(N__18177),
            .I(N__18045));
    InMux I__2749 (
            .O(N__18176),
            .I(N__18045));
    InMux I__2748 (
            .O(N__18175),
            .I(N__18045));
    InMux I__2747 (
            .O(N__18174),
            .I(N__18028));
    InMux I__2746 (
            .O(N__18173),
            .I(N__18028));
    InMux I__2745 (
            .O(N__18172),
            .I(N__18028));
    InMux I__2744 (
            .O(N__18171),
            .I(N__18028));
    InMux I__2743 (
            .O(N__18170),
            .I(N__18028));
    InMux I__2742 (
            .O(N__18169),
            .I(N__18028));
    InMux I__2741 (
            .O(N__18168),
            .I(N__18028));
    InMux I__2740 (
            .O(N__18167),
            .I(N__18028));
    LocalMux I__2739 (
            .O(N__18152),
            .I(N__18021));
    Span4Mux_h I__2738 (
            .O(N__18145),
            .I(N__18021));
    Span4Mux_s1_v I__2737 (
            .O(N__18140),
            .I(N__18021));
    LocalMux I__2736 (
            .O(N__18137),
            .I(N__18016));
    LocalMux I__2735 (
            .O(N__18134),
            .I(N__18016));
    Span4Mux_v I__2734 (
            .O(N__18127),
            .I(N__18011));
    LocalMux I__2733 (
            .O(N__18118),
            .I(N__18011));
    InMux I__2732 (
            .O(N__18117),
            .I(N__18008));
    InMux I__2731 (
            .O(N__18116),
            .I(N__17999));
    InMux I__2730 (
            .O(N__18115),
            .I(N__17999));
    InMux I__2729 (
            .O(N__18114),
            .I(N__17999));
    InMux I__2728 (
            .O(N__18113),
            .I(N__17999));
    Odrv4 I__2727 (
            .O(N__18108),
            .I(A_stk_delta_1));
    LocalMux I__2726 (
            .O(N__18101),
            .I(A_stk_delta_1));
    LocalMux I__2725 (
            .O(N__18088),
            .I(A_stk_delta_1));
    LocalMux I__2724 (
            .O(N__18073),
            .I(A_stk_delta_1));
    LocalMux I__2723 (
            .O(N__18058),
            .I(A_stk_delta_1));
    LocalMux I__2722 (
            .O(N__18045),
            .I(A_stk_delta_1));
    LocalMux I__2721 (
            .O(N__18028),
            .I(A_stk_delta_1));
    Odrv4 I__2720 (
            .O(N__18021),
            .I(A_stk_delta_1));
    Odrv12 I__2719 (
            .O(N__18016),
            .I(A_stk_delta_1));
    Odrv4 I__2718 (
            .O(N__18011),
            .I(A_stk_delta_1));
    LocalMux I__2717 (
            .O(N__18008),
            .I(A_stk_delta_1));
    LocalMux I__2716 (
            .O(N__17999),
            .I(A_stk_delta_1));
    InMux I__2715 (
            .O(N__17974),
            .I(N__17971));
    LocalMux I__2714 (
            .O(N__17971),
            .I(N__17968));
    Span4Mux_h I__2713 (
            .O(N__17968),
            .I(N__17964));
    InMux I__2712 (
            .O(N__17967),
            .I(N__17961));
    Odrv4 I__2711 (
            .O(N__17964),
            .I(\tok.A_stk.tail_2 ));
    LocalMux I__2710 (
            .O(N__17961),
            .I(\tok.A_stk.tail_2 ));
    CEMux I__2709 (
            .O(N__17956),
            .I(N__17952));
    CEMux I__2708 (
            .O(N__17955),
            .I(N__17949));
    LocalMux I__2707 (
            .O(N__17952),
            .I(N__17943));
    LocalMux I__2706 (
            .O(N__17949),
            .I(N__17940));
    CEMux I__2705 (
            .O(N__17948),
            .I(N__17937));
    CEMux I__2704 (
            .O(N__17947),
            .I(N__17928));
    CEMux I__2703 (
            .O(N__17946),
            .I(N__17920));
    Span4Mux_h I__2702 (
            .O(N__17943),
            .I(N__17916));
    Span4Mux_h I__2701 (
            .O(N__17940),
            .I(N__17911));
    LocalMux I__2700 (
            .O(N__17937),
            .I(N__17911));
    CEMux I__2699 (
            .O(N__17936),
            .I(N__17908));
    InMux I__2698 (
            .O(N__17935),
            .I(N__17905));
    CEMux I__2697 (
            .O(N__17934),
            .I(N__17897));
    CEMux I__2696 (
            .O(N__17933),
            .I(N__17894));
    CEMux I__2695 (
            .O(N__17932),
            .I(N__17891));
    CascadeMux I__2694 (
            .O(N__17931),
            .I(N__17888));
    LocalMux I__2693 (
            .O(N__17928),
            .I(N__17881));
    CEMux I__2692 (
            .O(N__17927),
            .I(N__17878));
    CEMux I__2691 (
            .O(N__17926),
            .I(N__17875));
    CEMux I__2690 (
            .O(N__17925),
            .I(N__17871));
    CEMux I__2689 (
            .O(N__17924),
            .I(N__17868));
    CEMux I__2688 (
            .O(N__17923),
            .I(N__17865));
    LocalMux I__2687 (
            .O(N__17920),
            .I(N__17862));
    CEMux I__2686 (
            .O(N__17919),
            .I(N__17859));
    Span4Mux_h I__2685 (
            .O(N__17916),
            .I(N__17852));
    Span4Mux_v I__2684 (
            .O(N__17911),
            .I(N__17852));
    LocalMux I__2683 (
            .O(N__17908),
            .I(N__17852));
    LocalMux I__2682 (
            .O(N__17905),
            .I(N__17849));
    InMux I__2681 (
            .O(N__17904),
            .I(N__17846));
    InMux I__2680 (
            .O(N__17903),
            .I(N__17841));
    InMux I__2679 (
            .O(N__17902),
            .I(N__17841));
    CEMux I__2678 (
            .O(N__17901),
            .I(N__17838));
    CEMux I__2677 (
            .O(N__17900),
            .I(N__17835));
    LocalMux I__2676 (
            .O(N__17897),
            .I(N__17828));
    LocalMux I__2675 (
            .O(N__17894),
            .I(N__17828));
    LocalMux I__2674 (
            .O(N__17891),
            .I(N__17828));
    InMux I__2673 (
            .O(N__17888),
            .I(N__17823));
    InMux I__2672 (
            .O(N__17887),
            .I(N__17823));
    CascadeMux I__2671 (
            .O(N__17886),
            .I(N__17820));
    CascadeMux I__2670 (
            .O(N__17885),
            .I(N__17817));
    CascadeMux I__2669 (
            .O(N__17884),
            .I(N__17814));
    Span4Mux_s2_v I__2668 (
            .O(N__17881),
            .I(N__17806));
    LocalMux I__2667 (
            .O(N__17878),
            .I(N__17806));
    LocalMux I__2666 (
            .O(N__17875),
            .I(N__17803));
    CEMux I__2665 (
            .O(N__17874),
            .I(N__17800));
    LocalMux I__2664 (
            .O(N__17871),
            .I(N__17795));
    LocalMux I__2663 (
            .O(N__17868),
            .I(N__17795));
    LocalMux I__2662 (
            .O(N__17865),
            .I(N__17792));
    Span4Mux_v I__2661 (
            .O(N__17862),
            .I(N__17787));
    LocalMux I__2660 (
            .O(N__17859),
            .I(N__17787));
    Span4Mux_s2_h I__2659 (
            .O(N__17852),
            .I(N__17782));
    Span4Mux_s2_h I__2658 (
            .O(N__17849),
            .I(N__17782));
    LocalMux I__2657 (
            .O(N__17846),
            .I(N__17779));
    LocalMux I__2656 (
            .O(N__17841),
            .I(N__17776));
    LocalMux I__2655 (
            .O(N__17838),
            .I(N__17767));
    LocalMux I__2654 (
            .O(N__17835),
            .I(N__17767));
    Span4Mux_v I__2653 (
            .O(N__17828),
            .I(N__17767));
    LocalMux I__2652 (
            .O(N__17823),
            .I(N__17767));
    InMux I__2651 (
            .O(N__17820),
            .I(N__17758));
    InMux I__2650 (
            .O(N__17817),
            .I(N__17758));
    InMux I__2649 (
            .O(N__17814),
            .I(N__17758));
    InMux I__2648 (
            .O(N__17813),
            .I(N__17758));
    CascadeMux I__2647 (
            .O(N__17812),
            .I(N__17754));
    CascadeMux I__2646 (
            .O(N__17811),
            .I(N__17750));
    Span4Mux_h I__2645 (
            .O(N__17806),
            .I(N__17746));
    Span4Mux_h I__2644 (
            .O(N__17803),
            .I(N__17741));
    LocalMux I__2643 (
            .O(N__17800),
            .I(N__17741));
    Span4Mux_v I__2642 (
            .O(N__17795),
            .I(N__17734));
    Span4Mux_v I__2641 (
            .O(N__17792),
            .I(N__17734));
    Span4Mux_v I__2640 (
            .O(N__17787),
            .I(N__17734));
    Span4Mux_v I__2639 (
            .O(N__17782),
            .I(N__17729));
    Span4Mux_h I__2638 (
            .O(N__17779),
            .I(N__17729));
    Span4Mux_h I__2637 (
            .O(N__17776),
            .I(N__17722));
    Span4Mux_s1_v I__2636 (
            .O(N__17767),
            .I(N__17722));
    LocalMux I__2635 (
            .O(N__17758),
            .I(N__17722));
    InMux I__2634 (
            .O(N__17757),
            .I(N__17719));
    InMux I__2633 (
            .O(N__17754),
            .I(N__17710));
    InMux I__2632 (
            .O(N__17753),
            .I(N__17710));
    InMux I__2631 (
            .O(N__17750),
            .I(N__17710));
    InMux I__2630 (
            .O(N__17749),
            .I(N__17710));
    Odrv4 I__2629 (
            .O(N__17746),
            .I(rd_15__N_300));
    Odrv4 I__2628 (
            .O(N__17741),
            .I(rd_15__N_300));
    Odrv4 I__2627 (
            .O(N__17734),
            .I(rd_15__N_300));
    Odrv4 I__2626 (
            .O(N__17729),
            .I(rd_15__N_300));
    Odrv4 I__2625 (
            .O(N__17722),
            .I(rd_15__N_300));
    LocalMux I__2624 (
            .O(N__17719),
            .I(rd_15__N_300));
    LocalMux I__2623 (
            .O(N__17710),
            .I(rd_15__N_300));
    InMux I__2622 (
            .O(N__17695),
            .I(N__17692));
    LocalMux I__2621 (
            .O(N__17692),
            .I(n10_adj_905));
    CascadeMux I__2620 (
            .O(N__17689),
            .I(\tok.n83_adj_764_cascade_ ));
    CascadeMux I__2619 (
            .O(N__17686),
            .I(\tok.ram.n6277_cascade_ ));
    CascadeMux I__2618 (
            .O(N__17683),
            .I(n10_cascade_));
    CascadeMux I__2617 (
            .O(N__17680),
            .I(N__17677));
    InMux I__2616 (
            .O(N__17677),
            .I(N__17674));
    LocalMux I__2615 (
            .O(N__17674),
            .I(N__17671));
    Span4Mux_h I__2614 (
            .O(N__17671),
            .I(N__17668));
    Span4Mux_v I__2613 (
            .O(N__17668),
            .I(N__17665));
    Odrv4 I__2612 (
            .O(N__17665),
            .I(\tok.tc_7 ));
    InMux I__2611 (
            .O(N__17662),
            .I(N__17659));
    LocalMux I__2610 (
            .O(N__17659),
            .I(\tok.n1635 ));
    CascadeMux I__2609 (
            .O(N__17656),
            .I(N__17653));
    InMux I__2608 (
            .O(N__17653),
            .I(N__17650));
    LocalMux I__2607 (
            .O(N__17650),
            .I(\tok.n6662 ));
    InMux I__2606 (
            .O(N__17647),
            .I(N__17644));
    LocalMux I__2605 (
            .O(N__17644),
            .I(\tok.n13_adj_790 ));
    InMux I__2604 (
            .O(N__17641),
            .I(N__17638));
    LocalMux I__2603 (
            .O(N__17638),
            .I(n10));
    InMux I__2602 (
            .O(N__17635),
            .I(\tok.n4817 ));
    InMux I__2601 (
            .O(N__17632),
            .I(\tok.n4818 ));
    CascadeMux I__2600 (
            .O(N__17629),
            .I(\tok.n13_adj_760_cascade_ ));
    CascadeMux I__2599 (
            .O(N__17626),
            .I(n10_adj_905_cascade_));
    CascadeMux I__2598 (
            .O(N__17623),
            .I(N__17620));
    InMux I__2597 (
            .O(N__17620),
            .I(N__17617));
    LocalMux I__2596 (
            .O(N__17617),
            .I(N__17614));
    Span4Mux_v I__2595 (
            .O(N__17614),
            .I(N__17611));
    Span4Mux_v I__2594 (
            .O(N__17611),
            .I(N__17608));
    Odrv4 I__2593 (
            .O(N__17608),
            .I(\tok.tc_5 ));
    CascadeMux I__2592 (
            .O(N__17605),
            .I(\tok.ram.n6263_cascade_ ));
    InMux I__2591 (
            .O(N__17602),
            .I(N__17599));
    LocalMux I__2590 (
            .O(N__17599),
            .I(\tok.n1530 ));
    CascadeMux I__2589 (
            .O(N__17596),
            .I(\tok.n83_adj_759_cascade_ ));
    CascadeMux I__2588 (
            .O(N__17593),
            .I(N__17590));
    InMux I__2587 (
            .O(N__17590),
            .I(N__17587));
    LocalMux I__2586 (
            .O(N__17587),
            .I(\tok.n6660 ));
    CascadeMux I__2585 (
            .O(N__17584),
            .I(\tok.n6_adj_699_cascade_ ));
    InMux I__2584 (
            .O(N__17581),
            .I(bfn_6_2_0_));
    InMux I__2583 (
            .O(N__17578),
            .I(\tok.n4812 ));
    InMux I__2582 (
            .O(N__17575),
            .I(\tok.n4813 ));
    InMux I__2581 (
            .O(N__17572),
            .I(\tok.n4814 ));
    InMux I__2580 (
            .O(N__17569),
            .I(\tok.n4815 ));
    InMux I__2579 (
            .O(N__17566),
            .I(\tok.n4816 ));
    CascadeMux I__2578 (
            .O(N__17563),
            .I(\tok.n262_adj_858_cascade_ ));
    InMux I__2577 (
            .O(N__17560),
            .I(N__17557));
    LocalMux I__2576 (
            .O(N__17557),
            .I(N__17554));
    Span12Mux_s7_v I__2575 (
            .O(N__17554),
            .I(N__17551));
    Odrv12 I__2574 (
            .O(N__17551),
            .I(\tok.n268 ));
    CascadeMux I__2573 (
            .O(N__17548),
            .I(N__17545));
    InMux I__2572 (
            .O(N__17545),
            .I(N__17542));
    LocalMux I__2571 (
            .O(N__17542),
            .I(N__17539));
    Odrv4 I__2570 (
            .O(N__17539),
            .I(\tok.n6315 ));
    DummyBuf I__2569 (
            .O(N__17536),
            .I(N__17532));
    DummyBuf I__2568 (
            .O(N__17535),
            .I(N__17529));
    InMux I__2567 (
            .O(N__17532),
            .I(N__17525));
    InMux I__2566 (
            .O(N__17529),
            .I(N__17522));
    SRMux I__2565 (
            .O(N__17528),
            .I(N__17519));
    LocalMux I__2564 (
            .O(N__17525),
            .I(N__17510));
    LocalMux I__2563 (
            .O(N__17522),
            .I(N__17510));
    LocalMux I__2562 (
            .O(N__17519),
            .I(N__17504));
    SRMux I__2561 (
            .O(N__17518),
            .I(N__17501));
    InMux I__2560 (
            .O(N__17517),
            .I(N__17498));
    InMux I__2559 (
            .O(N__17516),
            .I(N__17492));
    InMux I__2558 (
            .O(N__17515),
            .I(N__17492));
    Span4Mux_s1_h I__2557 (
            .O(N__17510),
            .I(N__17489));
    CascadeMux I__2556 (
            .O(N__17509),
            .I(N__17486));
    InMux I__2555 (
            .O(N__17508),
            .I(N__17482));
    InMux I__2554 (
            .O(N__17507),
            .I(N__17479));
    Span4Mux_v I__2553 (
            .O(N__17504),
            .I(N__17472));
    LocalMux I__2552 (
            .O(N__17501),
            .I(N__17472));
    LocalMux I__2551 (
            .O(N__17498),
            .I(N__17472));
    SRMux I__2550 (
            .O(N__17497),
            .I(N__17469));
    LocalMux I__2549 (
            .O(N__17492),
            .I(N__17466));
    Span4Mux_h I__2548 (
            .O(N__17489),
            .I(N__17463));
    InMux I__2547 (
            .O(N__17486),
            .I(N__17460));
    InMux I__2546 (
            .O(N__17485),
            .I(N__17457));
    LocalMux I__2545 (
            .O(N__17482),
            .I(N__17448));
    LocalMux I__2544 (
            .O(N__17479),
            .I(N__17448));
    Span4Mux_h I__2543 (
            .O(N__17472),
            .I(N__17448));
    LocalMux I__2542 (
            .O(N__17469),
            .I(N__17448));
    Span4Mux_v I__2541 (
            .O(N__17466),
            .I(N__17445));
    Sp12to4 I__2540 (
            .O(N__17463),
            .I(N__17440));
    LocalMux I__2539 (
            .O(N__17460),
            .I(N__17440));
    LocalMux I__2538 (
            .O(N__17457),
            .I(N__17437));
    Span4Mux_v I__2537 (
            .O(N__17448),
            .I(N__17434));
    Odrv4 I__2536 (
            .O(N__17445),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__2535 (
            .O(N__17440),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2534 (
            .O(N__17437),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2533 (
            .O(N__17434),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__2532 (
            .O(N__17425),
            .I(CONSTANT_ONE_NET_cascade_));
    InMux I__2531 (
            .O(N__17422),
            .I(N__17418));
    InMux I__2530 (
            .O(N__17421),
            .I(N__17415));
    LocalMux I__2529 (
            .O(N__17418),
            .I(N__17409));
    LocalMux I__2528 (
            .O(N__17415),
            .I(N__17409));
    InMux I__2527 (
            .O(N__17414),
            .I(N__17406));
    Span12Mux_s5_v I__2526 (
            .O(N__17409),
            .I(N__17403));
    LocalMux I__2525 (
            .O(N__17406),
            .I(\tok.n239 ));
    Odrv12 I__2524 (
            .O(N__17403),
            .I(\tok.n239 ));
    CascadeMux I__2523 (
            .O(N__17398),
            .I(N__17395));
    InMux I__2522 (
            .O(N__17395),
            .I(N__17392));
    LocalMux I__2521 (
            .O(N__17392),
            .I(N__17389));
    Span4Mux_s2_h I__2520 (
            .O(N__17389),
            .I(N__17386));
    Span4Mux_h I__2519 (
            .O(N__17386),
            .I(N__17383));
    Odrv4 I__2518 (
            .O(N__17383),
            .I(sender_2));
    InMux I__2517 (
            .O(N__17380),
            .I(N__17377));
    LocalMux I__2516 (
            .O(N__17377),
            .I(N__17374));
    Span4Mux_h I__2515 (
            .O(N__17374),
            .I(N__17371));
    Odrv4 I__2514 (
            .O(N__17371),
            .I(\tok.n6347 ));
    InMux I__2513 (
            .O(N__17368),
            .I(N__17365));
    LocalMux I__2512 (
            .O(N__17365),
            .I(\tok.n197_adj_693 ));
    CascadeMux I__2511 (
            .O(N__17362),
            .I(\tok.n248_adj_694_cascade_ ));
    InMux I__2510 (
            .O(N__17359),
            .I(N__17356));
    LocalMux I__2509 (
            .O(N__17356),
            .I(\tok.n242_adj_695 ));
    CascadeMux I__2508 (
            .O(N__17353),
            .I(\tok.n200_adj_696_cascade_ ));
    CascadeMux I__2507 (
            .O(N__17350),
            .I(\tok.n200_adj_655_cascade_ ));
    CascadeMux I__2506 (
            .O(N__17347),
            .I(\tok.n6_adj_658_cascade_ ));
    CascadeMux I__2505 (
            .O(N__17344),
            .I(\tok.n6_adj_832_cascade_ ));
    InMux I__2504 (
            .O(N__17341),
            .I(N__17338));
    LocalMux I__2503 (
            .O(N__17338),
            .I(N__17335));
    Span4Mux_h I__2502 (
            .O(N__17335),
            .I(N__17332));
    Span4Mux_s2_h I__2501 (
            .O(N__17332),
            .I(N__17329));
    Odrv4 I__2500 (
            .O(N__17329),
            .I(\tok.n6383 ));
    InMux I__2499 (
            .O(N__17326),
            .I(N__17323));
    LocalMux I__2498 (
            .O(N__17323),
            .I(\tok.n242_adj_654 ));
    CascadeMux I__2497 (
            .O(N__17320),
            .I(N__17315));
    InMux I__2496 (
            .O(N__17319),
            .I(N__17310));
    InMux I__2495 (
            .O(N__17318),
            .I(N__17307));
    InMux I__2494 (
            .O(N__17315),
            .I(N__17304));
    InMux I__2493 (
            .O(N__17314),
            .I(N__17299));
    InMux I__2492 (
            .O(N__17313),
            .I(N__17299));
    LocalMux I__2491 (
            .O(N__17310),
            .I(N__17289));
    LocalMux I__2490 (
            .O(N__17307),
            .I(N__17289));
    LocalMux I__2489 (
            .O(N__17304),
            .I(N__17289));
    LocalMux I__2488 (
            .O(N__17299),
            .I(N__17289));
    InMux I__2487 (
            .O(N__17298),
            .I(N__17285));
    Span4Mux_v I__2486 (
            .O(N__17289),
            .I(N__17282));
    InMux I__2485 (
            .O(N__17288),
            .I(N__17279));
    LocalMux I__2484 (
            .O(N__17285),
            .I(N__17276));
    Span4Mux_h I__2483 (
            .O(N__17282),
            .I(N__17273));
    LocalMux I__2482 (
            .O(N__17279),
            .I(\tok.S_13 ));
    Odrv4 I__2481 (
            .O(N__17276),
            .I(\tok.S_13 ));
    Odrv4 I__2480 (
            .O(N__17273),
            .I(\tok.S_13 ));
    CascadeMux I__2479 (
            .O(N__17266),
            .I(N__17262));
    CascadeMux I__2478 (
            .O(N__17265),
            .I(N__17258));
    InMux I__2477 (
            .O(N__17262),
            .I(N__17255));
    CascadeMux I__2476 (
            .O(N__17261),
            .I(N__17252));
    InMux I__2475 (
            .O(N__17258),
            .I(N__17246));
    LocalMux I__2474 (
            .O(N__17255),
            .I(N__17243));
    InMux I__2473 (
            .O(N__17252),
            .I(N__17240));
    InMux I__2472 (
            .O(N__17251),
            .I(N__17235));
    InMux I__2471 (
            .O(N__17250),
            .I(N__17235));
    InMux I__2470 (
            .O(N__17249),
            .I(N__17232));
    LocalMux I__2469 (
            .O(N__17246),
            .I(N__17229));
    Span4Mux_s3_v I__2468 (
            .O(N__17243),
            .I(N__17224));
    LocalMux I__2467 (
            .O(N__17240),
            .I(N__17224));
    LocalMux I__2466 (
            .O(N__17235),
            .I(N__17221));
    LocalMux I__2465 (
            .O(N__17232),
            .I(N__17217));
    Span4Mux_v I__2464 (
            .O(N__17229),
            .I(N__17214));
    Span4Mux_v I__2463 (
            .O(N__17224),
            .I(N__17209));
    Span4Mux_s3_v I__2462 (
            .O(N__17221),
            .I(N__17209));
    InMux I__2461 (
            .O(N__17220),
            .I(N__17206));
    Span4Mux_v I__2460 (
            .O(N__17217),
            .I(N__17203));
    Span4Mux_h I__2459 (
            .O(N__17214),
            .I(N__17198));
    Span4Mux_h I__2458 (
            .O(N__17209),
            .I(N__17198));
    LocalMux I__2457 (
            .O(N__17206),
            .I(\tok.S_8 ));
    Odrv4 I__2456 (
            .O(N__17203),
            .I(\tok.S_8 ));
    Odrv4 I__2455 (
            .O(N__17198),
            .I(\tok.S_8 ));
    CascadeMux I__2454 (
            .O(N__17191),
            .I(\tok.n14_adj_844_cascade_ ));
    InMux I__2453 (
            .O(N__17188),
            .I(N__17185));
    LocalMux I__2452 (
            .O(N__17185),
            .I(N__17182));
    Odrv12 I__2451 (
            .O(N__17182),
            .I(\tok.n20_adj_845 ));
    InMux I__2450 (
            .O(N__17179),
            .I(N__17176));
    LocalMux I__2449 (
            .O(N__17176),
            .I(\tok.n26_adj_851 ));
    CascadeMux I__2448 (
            .O(N__17173),
            .I(\tok.n6324_cascade_ ));
    InMux I__2447 (
            .O(N__17170),
            .I(N__17167));
    LocalMux I__2446 (
            .O(N__17167),
            .I(\tok.n6460 ));
    CascadeMux I__2445 (
            .O(N__17164),
            .I(N__17161));
    InMux I__2444 (
            .O(N__17161),
            .I(N__17158));
    LocalMux I__2443 (
            .O(N__17158),
            .I(\tok.n161_adj_825 ));
    InMux I__2442 (
            .O(N__17155),
            .I(N__17152));
    LocalMux I__2441 (
            .O(N__17152),
            .I(\tok.n197_adj_826 ));
    InMux I__2440 (
            .O(N__17149),
            .I(N__17146));
    LocalMux I__2439 (
            .O(N__17146),
            .I(N__17143));
    Span4Mux_h I__2438 (
            .O(N__17143),
            .I(N__17140));
    Odrv4 I__2437 (
            .O(N__17140),
            .I(\tok.n18_adj_850 ));
    InMux I__2436 (
            .O(N__17137),
            .I(N__17134));
    LocalMux I__2435 (
            .O(N__17134),
            .I(\tok.n17_adj_853 ));
    CascadeMux I__2434 (
            .O(N__17131),
            .I(\tok.n31_cascade_ ));
    InMux I__2433 (
            .O(N__17128),
            .I(N__17125));
    LocalMux I__2432 (
            .O(N__17125),
            .I(N__17122));
    Odrv4 I__2431 (
            .O(N__17122),
            .I(\tok.n299 ));
    CascadeMux I__2430 (
            .O(N__17119),
            .I(N__17116));
    InMux I__2429 (
            .O(N__17116),
            .I(N__17113));
    LocalMux I__2428 (
            .O(N__17113),
            .I(\tok.n6446 ));
    InMux I__2427 (
            .O(N__17110),
            .I(N__17107));
    LocalMux I__2426 (
            .O(N__17107),
            .I(N__17104));
    Odrv12 I__2425 (
            .O(N__17104),
            .I(\tok.n308 ));
    InMux I__2424 (
            .O(N__17101),
            .I(N__17098));
    LocalMux I__2423 (
            .O(N__17098),
            .I(N__17095));
    Odrv4 I__2422 (
            .O(N__17095),
            .I(\tok.n294 ));
    InMux I__2421 (
            .O(N__17092),
            .I(N__17089));
    LocalMux I__2420 (
            .O(N__17089),
            .I(\tok.n161_adj_667 ));
    CascadeMux I__2419 (
            .O(N__17086),
            .I(\tok.n6371_cascade_ ));
    CascadeMux I__2418 (
            .O(N__17083),
            .I(N__17080));
    InMux I__2417 (
            .O(N__17080),
            .I(N__17077));
    LocalMux I__2416 (
            .O(N__17077),
            .I(\tok.n248_adj_653 ));
    InMux I__2415 (
            .O(N__17074),
            .I(\tok.n4795 ));
    InMux I__2414 (
            .O(N__17071),
            .I(bfn_5_10_0_));
    InMux I__2413 (
            .O(N__17068),
            .I(N__17065));
    LocalMux I__2412 (
            .O(N__17065),
            .I(N__17062));
    Odrv4 I__2411 (
            .O(N__17062),
            .I(\tok.n293 ));
    InMux I__2410 (
            .O(N__17059),
            .I(N__17056));
    LocalMux I__2409 (
            .O(N__17056),
            .I(\tok.n297 ));
    InMux I__2408 (
            .O(N__17053),
            .I(N__17050));
    LocalMux I__2407 (
            .O(N__17050),
            .I(\tok.n310 ));
    InMux I__2406 (
            .O(N__17047),
            .I(N__17044));
    LocalMux I__2405 (
            .O(N__17044),
            .I(\tok.n6452 ));
    InMux I__2404 (
            .O(N__17041),
            .I(N__17038));
    LocalMux I__2403 (
            .O(N__17038),
            .I(\tok.n2579 ));
    InMux I__2402 (
            .O(N__17035),
            .I(N__17032));
    LocalMux I__2401 (
            .O(N__17032),
            .I(\tok.n6392 ));
    InMux I__2400 (
            .O(N__17029),
            .I(N__17026));
    LocalMux I__2399 (
            .O(N__17026),
            .I(\tok.n6421 ));
    InMux I__2398 (
            .O(N__17023),
            .I(N__17020));
    LocalMux I__2397 (
            .O(N__17020),
            .I(\tok.n300 ));
    InMux I__2396 (
            .O(N__17017),
            .I(\tok.n4787 ));
    InMux I__2395 (
            .O(N__17014),
            .I(N__17008));
    InMux I__2394 (
            .O(N__17013),
            .I(N__17005));
    InMux I__2393 (
            .O(N__17012),
            .I(N__17000));
    InMux I__2392 (
            .O(N__17011),
            .I(N__17000));
    LocalMux I__2391 (
            .O(N__17008),
            .I(N__16997));
    LocalMux I__2390 (
            .O(N__17005),
            .I(N__16992));
    LocalMux I__2389 (
            .O(N__17000),
            .I(N__16992));
    Span4Mux_v I__2388 (
            .O(N__16997),
            .I(N__16989));
    Span4Mux_v I__2387 (
            .O(N__16992),
            .I(N__16986));
    Odrv4 I__2386 (
            .O(N__16989),
            .I(\tok.n21_adj_660 ));
    Odrv4 I__2385 (
            .O(N__16986),
            .I(\tok.n21_adj_660 ));
    CascadeMux I__2384 (
            .O(N__16981),
            .I(N__16978));
    InMux I__2383 (
            .O(N__16978),
            .I(N__16975));
    LocalMux I__2382 (
            .O(N__16975),
            .I(N__16972));
    Odrv4 I__2381 (
            .O(N__16972),
            .I(\tok.n318 ));
    InMux I__2380 (
            .O(N__16969),
            .I(bfn_5_9_0_));
    InMux I__2379 (
            .O(N__16966),
            .I(\tok.n4789 ));
    InMux I__2378 (
            .O(N__16963),
            .I(\tok.n4790 ));
    CascadeMux I__2377 (
            .O(N__16960),
            .I(N__16957));
    InMux I__2376 (
            .O(N__16957),
            .I(N__16954));
    LocalMux I__2375 (
            .O(N__16954),
            .I(N__16951));
    Odrv4 I__2374 (
            .O(N__16951),
            .I(\tok.n315 ));
    InMux I__2373 (
            .O(N__16948),
            .I(\tok.n4791 ));
    InMux I__2372 (
            .O(N__16945),
            .I(\tok.n4792 ));
    CascadeMux I__2371 (
            .O(N__16942),
            .I(N__16939));
    InMux I__2370 (
            .O(N__16939),
            .I(N__16936));
    LocalMux I__2369 (
            .O(N__16936),
            .I(N__16933));
    Odrv4 I__2368 (
            .O(N__16933),
            .I(\tok.n313 ));
    InMux I__2367 (
            .O(N__16930),
            .I(\tok.n4793 ));
    InMux I__2366 (
            .O(N__16927),
            .I(N__16923));
    CascadeMux I__2365 (
            .O(N__16926),
            .I(N__16920));
    LocalMux I__2364 (
            .O(N__16923),
            .I(N__16917));
    InMux I__2363 (
            .O(N__16920),
            .I(N__16914));
    Span4Mux_s2_h I__2362 (
            .O(N__16917),
            .I(N__16909));
    LocalMux I__2361 (
            .O(N__16914),
            .I(N__16909));
    Span4Mux_h I__2360 (
            .O(N__16909),
            .I(N__16906));
    Sp12to4 I__2359 (
            .O(N__16906),
            .I(N__16903));
    Odrv12 I__2358 (
            .O(N__16903),
            .I(\tok.n312 ));
    InMux I__2357 (
            .O(N__16900),
            .I(N__16897));
    LocalMux I__2356 (
            .O(N__16897),
            .I(N__16894));
    Span4Mux_h I__2355 (
            .O(N__16894),
            .I(N__16891));
    Odrv4 I__2354 (
            .O(N__16891),
            .I(\tok.n295 ));
    InMux I__2353 (
            .O(N__16888),
            .I(\tok.n4794 ));
    InMux I__2352 (
            .O(N__16885),
            .I(N__16881));
    CascadeMux I__2351 (
            .O(N__16884),
            .I(N__16878));
    LocalMux I__2350 (
            .O(N__16881),
            .I(N__16875));
    InMux I__2349 (
            .O(N__16878),
            .I(N__16872));
    Odrv4 I__2348 (
            .O(N__16875),
            .I(\tok.key_rd_8 ));
    LocalMux I__2347 (
            .O(N__16872),
            .I(\tok.key_rd_8 ));
    CascadeMux I__2346 (
            .O(N__16867),
            .I(\tok.n20_cascade_ ));
    InMux I__2345 (
            .O(N__16864),
            .I(N__16861));
    LocalMux I__2344 (
            .O(N__16861),
            .I(N__16858));
    Odrv4 I__2343 (
            .O(N__16858),
            .I(\tok.n26_adj_645 ));
    InMux I__2342 (
            .O(N__16855),
            .I(N__16851));
    InMux I__2341 (
            .O(N__16854),
            .I(N__16848));
    LocalMux I__2340 (
            .O(N__16851),
            .I(N__16845));
    LocalMux I__2339 (
            .O(N__16848),
            .I(\tok.key_rd_13 ));
    Odrv4 I__2338 (
            .O(N__16845),
            .I(\tok.key_rd_13 ));
    InMux I__2337 (
            .O(N__16840),
            .I(N__16837));
    LocalMux I__2336 (
            .O(N__16837),
            .I(\tok.n14_adj_644 ));
    InMux I__2335 (
            .O(N__16834),
            .I(bfn_5_8_0_));
    InMux I__2334 (
            .O(N__16831),
            .I(\tok.n4782 ));
    InMux I__2333 (
            .O(N__16828),
            .I(\tok.n4783 ));
    CascadeMux I__2332 (
            .O(N__16825),
            .I(N__16822));
    InMux I__2331 (
            .O(N__16822),
            .I(N__16819));
    LocalMux I__2330 (
            .O(N__16819),
            .I(\tok.n127 ));
    InMux I__2329 (
            .O(N__16816),
            .I(\tok.n4784 ));
    InMux I__2328 (
            .O(N__16813),
            .I(N__16810));
    LocalMux I__2327 (
            .O(N__16810),
            .I(\tok.n6557 ));
    InMux I__2326 (
            .O(N__16807),
            .I(\tok.n4785 ));
    InMux I__2325 (
            .O(N__16804),
            .I(N__16801));
    LocalMux I__2324 (
            .O(N__16801),
            .I(\tok.n320 ));
    InMux I__2323 (
            .O(N__16798),
            .I(\tok.n4786 ));
    InMux I__2322 (
            .O(N__16795),
            .I(N__16789));
    InMux I__2321 (
            .O(N__16794),
            .I(N__16789));
    LocalMux I__2320 (
            .O(N__16789),
            .I(\tok.n12 ));
    CascadeMux I__2319 (
            .O(N__16786),
            .I(N__16783));
    InMux I__2318 (
            .O(N__16783),
            .I(N__16776));
    CascadeMux I__2317 (
            .O(N__16782),
            .I(N__16772));
    InMux I__2316 (
            .O(N__16781),
            .I(N__16766));
    InMux I__2315 (
            .O(N__16780),
            .I(N__16761));
    InMux I__2314 (
            .O(N__16779),
            .I(N__16761));
    LocalMux I__2313 (
            .O(N__16776),
            .I(N__16758));
    InMux I__2312 (
            .O(N__16775),
            .I(N__16755));
    InMux I__2311 (
            .O(N__16772),
            .I(N__16748));
    InMux I__2310 (
            .O(N__16771),
            .I(N__16748));
    InMux I__2309 (
            .O(N__16770),
            .I(N__16748));
    InMux I__2308 (
            .O(N__16769),
            .I(N__16745));
    LocalMux I__2307 (
            .O(N__16766),
            .I(N__16740));
    LocalMux I__2306 (
            .O(N__16761),
            .I(N__16740));
    Odrv4 I__2305 (
            .O(N__16758),
            .I(\tok.n796 ));
    LocalMux I__2304 (
            .O(N__16755),
            .I(\tok.n796 ));
    LocalMux I__2303 (
            .O(N__16748),
            .I(\tok.n796 ));
    LocalMux I__2302 (
            .O(N__16745),
            .I(\tok.n796 ));
    Odrv4 I__2301 (
            .O(N__16740),
            .I(\tok.n796 ));
    InMux I__2300 (
            .O(N__16729),
            .I(N__16720));
    InMux I__2299 (
            .O(N__16728),
            .I(N__16720));
    InMux I__2298 (
            .O(N__16727),
            .I(N__16720));
    LocalMux I__2297 (
            .O(N__16720),
            .I(\tok.n2702 ));
    InMux I__2296 (
            .O(N__16717),
            .I(N__16711));
    InMux I__2295 (
            .O(N__16716),
            .I(N__16704));
    InMux I__2294 (
            .O(N__16715),
            .I(N__16704));
    InMux I__2293 (
            .O(N__16714),
            .I(N__16704));
    LocalMux I__2292 (
            .O(N__16711),
            .I(\tok.uart_stall ));
    LocalMux I__2291 (
            .O(N__16704),
            .I(\tok.uart_stall ));
    InMux I__2290 (
            .O(N__16699),
            .I(N__16696));
    LocalMux I__2289 (
            .O(N__16696),
            .I(\tok.n6203 ));
    InMux I__2288 (
            .O(N__16693),
            .I(N__16690));
    LocalMux I__2287 (
            .O(N__16690),
            .I(\tok.search_clk_N_137 ));
    CascadeMux I__2286 (
            .O(N__16687),
            .I(\tok.n31_adj_637_cascade_ ));
    InMux I__2285 (
            .O(N__16684),
            .I(N__16681));
    LocalMux I__2284 (
            .O(N__16681),
            .I(\tok.n6170 ));
    InMux I__2283 (
            .O(N__16678),
            .I(N__16672));
    InMux I__2282 (
            .O(N__16677),
            .I(N__16672));
    LocalMux I__2281 (
            .O(N__16672),
            .I(N__16663));
    InMux I__2280 (
            .O(N__16671),
            .I(N__16660));
    InMux I__2279 (
            .O(N__16670),
            .I(N__16657));
    InMux I__2278 (
            .O(N__16669),
            .I(N__16648));
    InMux I__2277 (
            .O(N__16668),
            .I(N__16648));
    InMux I__2276 (
            .O(N__16667),
            .I(N__16648));
    InMux I__2275 (
            .O(N__16666),
            .I(N__16648));
    Span12Mux_s5_v I__2274 (
            .O(N__16663),
            .I(N__16643));
    LocalMux I__2273 (
            .O(N__16660),
            .I(N__16643));
    LocalMux I__2272 (
            .O(N__16657),
            .I(\tok.n30 ));
    LocalMux I__2271 (
            .O(N__16648),
            .I(\tok.n30 ));
    Odrv12 I__2270 (
            .O(N__16643),
            .I(\tok.n30 ));
    CascadeMux I__2269 (
            .O(N__16636),
            .I(\tok.n221_adj_753_cascade_ ));
    InMux I__2268 (
            .O(N__16633),
            .I(N__16630));
    LocalMux I__2267 (
            .O(N__16630),
            .I(N__16626));
    InMux I__2266 (
            .O(N__16629),
            .I(N__16623));
    Span4Mux_h I__2265 (
            .O(N__16626),
            .I(N__16620));
    LocalMux I__2264 (
            .O(N__16623),
            .I(\tok.key_rd_3 ));
    Odrv4 I__2263 (
            .O(N__16620),
            .I(\tok.key_rd_3 ));
    CascadeMux I__2262 (
            .O(N__16615),
            .I(N__16612));
    InMux I__2261 (
            .O(N__16612),
            .I(N__16609));
    LocalMux I__2260 (
            .O(N__16609),
            .I(N__16605));
    InMux I__2259 (
            .O(N__16608),
            .I(N__16602));
    Span4Mux_h I__2258 (
            .O(N__16605),
            .I(N__16599));
    LocalMux I__2257 (
            .O(N__16602),
            .I(\tok.key_rd_5 ));
    Odrv4 I__2256 (
            .O(N__16599),
            .I(\tok.key_rd_5 ));
    CascadeMux I__2255 (
            .O(N__16594),
            .I(\tok.n9_adj_651_cascade_ ));
    InMux I__2254 (
            .O(N__16591),
            .I(N__16588));
    LocalMux I__2253 (
            .O(N__16588),
            .I(N__16585));
    Odrv4 I__2252 (
            .O(N__16585),
            .I(\tok.n13 ));
    CascadeMux I__2251 (
            .O(N__16582),
            .I(n15_cascade_));
    CascadeMux I__2250 (
            .O(N__16579),
            .I(\tok.n6_adj_687_cascade_ ));
    InMux I__2249 (
            .O(N__16576),
            .I(N__16572));
    InMux I__2248 (
            .O(N__16575),
            .I(N__16569));
    LocalMux I__2247 (
            .O(N__16572),
            .I(N__16565));
    LocalMux I__2246 (
            .O(N__16569),
            .I(N__16562));
    InMux I__2245 (
            .O(N__16568),
            .I(N__16559));
    Odrv4 I__2244 (
            .O(N__16565),
            .I(\tok.n4_adj_641 ));
    Odrv4 I__2243 (
            .O(N__16562),
            .I(\tok.n4_adj_641 ));
    LocalMux I__2242 (
            .O(N__16559),
            .I(\tok.n4_adj_641 ));
    InMux I__2241 (
            .O(N__16552),
            .I(N__16549));
    LocalMux I__2240 (
            .O(N__16549),
            .I(\tok.n5 ));
    CascadeMux I__2239 (
            .O(N__16546),
            .I(\tok.n796_cascade_ ));
    CascadeMux I__2238 (
            .O(N__16543),
            .I(\tok.n80_cascade_ ));
    CascadeMux I__2237 (
            .O(N__16540),
            .I(\tok.n89_cascade_ ));
    CascadeMux I__2236 (
            .O(N__16537),
            .I(\tok.n83_adj_734_cascade_ ));
    InMux I__2235 (
            .O(N__16534),
            .I(N__16531));
    LocalMux I__2234 (
            .O(N__16531),
            .I(\tok.n6279 ));
    CascadeMux I__2233 (
            .O(N__16528),
            .I(N__16524));
    InMux I__2232 (
            .O(N__16527),
            .I(N__16519));
    InMux I__2231 (
            .O(N__16524),
            .I(N__16519));
    LocalMux I__2230 (
            .O(N__16519),
            .I(N__16516));
    Span4Mux_v I__2229 (
            .O(N__16516),
            .I(N__16513));
    Span4Mux_v I__2228 (
            .O(N__16513),
            .I(N__16510));
    Odrv4 I__2227 (
            .O(N__16510),
            .I(\tok.table_rd_0 ));
    InMux I__2226 (
            .O(N__16507),
            .I(N__16504));
    LocalMux I__2225 (
            .O(N__16504),
            .I(N__16501));
    Span4Mux_h I__2224 (
            .O(N__16501),
            .I(N__16498));
    Span4Mux_v I__2223 (
            .O(N__16498),
            .I(N__16495));
    Odrv4 I__2222 (
            .O(N__16495),
            .I(\tok.table_wr_data_14 ));
    InMux I__2221 (
            .O(N__16492),
            .I(N__16489));
    LocalMux I__2220 (
            .O(N__16489),
            .I(N__16486));
    Span4Mux_h I__2219 (
            .O(N__16486),
            .I(N__16483));
    Span4Mux_v I__2218 (
            .O(N__16483),
            .I(N__16480));
    Odrv4 I__2217 (
            .O(N__16480),
            .I(\tok.table_wr_data_11 ));
    InMux I__2216 (
            .O(N__16477),
            .I(N__16474));
    LocalMux I__2215 (
            .O(N__16474),
            .I(N__16471));
    Span4Mux_v I__2214 (
            .O(N__16471),
            .I(N__16468));
    Odrv4 I__2213 (
            .O(N__16468),
            .I(\tok.table_wr_data_12 ));
    InMux I__2212 (
            .O(N__16465),
            .I(N__16462));
    LocalMux I__2211 (
            .O(N__16462),
            .I(\tok.n2696 ));
    CascadeMux I__2210 (
            .O(N__16459),
            .I(\tok.ram.n6266_cascade_ ));
    CascadeMux I__2209 (
            .O(N__16456),
            .I(\tok.n1495_cascade_ ));
    InMux I__2208 (
            .O(N__16453),
            .I(N__16450));
    LocalMux I__2207 (
            .O(N__16450),
            .I(\tok.n13_adj_766 ));
    InMux I__2206 (
            .O(N__16447),
            .I(N__16444));
    LocalMux I__2205 (
            .O(N__16444),
            .I(n10_adj_907));
    CascadeMux I__2204 (
            .O(N__16441),
            .I(n10_adj_907_cascade_));
    CascadeMux I__2203 (
            .O(N__16438),
            .I(N__16435));
    InMux I__2202 (
            .O(N__16435),
            .I(N__16432));
    LocalMux I__2201 (
            .O(N__16432),
            .I(N__16429));
    Span4Mux_v I__2200 (
            .O(N__16429),
            .I(N__16426));
    Span4Mux_v I__2199 (
            .O(N__16426),
            .I(N__16423));
    Odrv4 I__2198 (
            .O(N__16423),
            .I(\tok.tc_6 ));
    CascadeMux I__2197 (
            .O(N__16420),
            .I(\tok.n83_adj_765_cascade_ ));
    InMux I__2196 (
            .O(N__16417),
            .I(N__16414));
    LocalMux I__2195 (
            .O(N__16414),
            .I(\tok.n6435 ));
    CascadeMux I__2194 (
            .O(N__16411),
            .I(\tok.n6283_cascade_ ));
    CascadeMux I__2193 (
            .O(N__16408),
            .I(N__16405));
    InMux I__2192 (
            .O(N__16405),
            .I(N__16399));
    InMux I__2191 (
            .O(N__16404),
            .I(N__16399));
    LocalMux I__2190 (
            .O(N__16399),
            .I(\tok.A_stk.tail_7 ));
    CascadeMux I__2189 (
            .O(N__16396),
            .I(N__16393));
    InMux I__2188 (
            .O(N__16393),
            .I(N__16390));
    LocalMux I__2187 (
            .O(N__16390),
            .I(N__16386));
    InMux I__2186 (
            .O(N__16389),
            .I(N__16383));
    Odrv4 I__2185 (
            .O(N__16386),
            .I(tail_97));
    LocalMux I__2184 (
            .O(N__16383),
            .I(tail_97));
    InMux I__2183 (
            .O(N__16378),
            .I(N__16374));
    InMux I__2182 (
            .O(N__16377),
            .I(N__16371));
    LocalMux I__2181 (
            .O(N__16374),
            .I(tail_113));
    LocalMux I__2180 (
            .O(N__16371),
            .I(tail_113));
    InMux I__2179 (
            .O(N__16366),
            .I(N__16362));
    InMux I__2178 (
            .O(N__16365),
            .I(N__16359));
    LocalMux I__2177 (
            .O(N__16362),
            .I(tail_108));
    LocalMux I__2176 (
            .O(N__16359),
            .I(tail_108));
    CascadeMux I__2175 (
            .O(N__16354),
            .I(N__16351));
    InMux I__2174 (
            .O(N__16351),
            .I(N__16347));
    InMux I__2173 (
            .O(N__16350),
            .I(N__16344));
    LocalMux I__2172 (
            .O(N__16347),
            .I(tail_124));
    LocalMux I__2171 (
            .O(N__16344),
            .I(tail_124));
    InMux I__2170 (
            .O(N__16339),
            .I(N__16336));
    LocalMux I__2169 (
            .O(N__16336),
            .I(N__16333));
    Span4Mux_v I__2168 (
            .O(N__16333),
            .I(N__16330));
    Span4Mux_v I__2167 (
            .O(N__16330),
            .I(N__16327));
    Odrv4 I__2166 (
            .O(N__16327),
            .I(\tok.table_wr_data_3 ));
    InMux I__2165 (
            .O(N__16324),
            .I(N__16321));
    LocalMux I__2164 (
            .O(N__16321),
            .I(N__16318));
    Span4Mux_v I__2163 (
            .O(N__16318),
            .I(N__16315));
    Span4Mux_v I__2162 (
            .O(N__16315),
            .I(N__16312));
    Odrv4 I__2161 (
            .O(N__16312),
            .I(table_wr_data_1));
    InMux I__2160 (
            .O(N__16309),
            .I(N__16306));
    LocalMux I__2159 (
            .O(N__16306),
            .I(N__16303));
    Span4Mux_v I__2158 (
            .O(N__16303),
            .I(N__16300));
    Span4Mux_v I__2157 (
            .O(N__16300),
            .I(N__16297));
    Odrv4 I__2156 (
            .O(N__16297),
            .I(\tok.table_wr_data_6 ));
    InMux I__2155 (
            .O(N__16294),
            .I(N__16291));
    LocalMux I__2154 (
            .O(N__16291),
            .I(N__16288));
    Span12Mux_v I__2153 (
            .O(N__16288),
            .I(N__16285));
    Odrv12 I__2152 (
            .O(N__16285),
            .I(\tok.table_wr_data_4 ));
    InMux I__2151 (
            .O(N__16282),
            .I(N__16279));
    LocalMux I__2150 (
            .O(N__16279),
            .I(N__16276));
    Span4Mux_v I__2149 (
            .O(N__16276),
            .I(N__16273));
    Span4Mux_v I__2148 (
            .O(N__16273),
            .I(N__16270));
    Odrv4 I__2147 (
            .O(N__16270),
            .I(\tok.table_wr_data_2 ));
    InMux I__2146 (
            .O(N__16267),
            .I(N__16264));
    LocalMux I__2145 (
            .O(N__16264),
            .I(\tok.n6412 ));
    InMux I__2144 (
            .O(N__16261),
            .I(N__16257));
    CascadeMux I__2143 (
            .O(N__16260),
            .I(N__16254));
    LocalMux I__2142 (
            .O(N__16257),
            .I(N__16251));
    InMux I__2141 (
            .O(N__16254),
            .I(N__16248));
    Odrv4 I__2140 (
            .O(N__16251),
            .I(tail_119));
    LocalMux I__2139 (
            .O(N__16248),
            .I(tail_119));
    InMux I__2138 (
            .O(N__16243),
            .I(N__16240));
    LocalMux I__2137 (
            .O(N__16240),
            .I(N__16236));
    InMux I__2136 (
            .O(N__16239),
            .I(N__16233));
    Odrv12 I__2135 (
            .O(N__16236),
            .I(tail_103));
    LocalMux I__2134 (
            .O(N__16233),
            .I(tail_103));
    InMux I__2133 (
            .O(N__16228),
            .I(N__16222));
    InMux I__2132 (
            .O(N__16227),
            .I(N__16222));
    LocalMux I__2131 (
            .O(N__16222),
            .I(\tok.A_stk.tail_87 ));
    InMux I__2130 (
            .O(N__16219),
            .I(N__16213));
    InMux I__2129 (
            .O(N__16218),
            .I(N__16213));
    LocalMux I__2128 (
            .O(N__16213),
            .I(\tok.A_stk.tail_71 ));
    InMux I__2127 (
            .O(N__16210),
            .I(N__16204));
    InMux I__2126 (
            .O(N__16209),
            .I(N__16204));
    LocalMux I__2125 (
            .O(N__16204),
            .I(\tok.A_stk.tail_55 ));
    InMux I__2124 (
            .O(N__16201),
            .I(N__16195));
    InMux I__2123 (
            .O(N__16200),
            .I(N__16195));
    LocalMux I__2122 (
            .O(N__16195),
            .I(\tok.A_stk.tail_39 ));
    InMux I__2121 (
            .O(N__16192),
            .I(N__16188));
    InMux I__2120 (
            .O(N__16191),
            .I(N__16185));
    LocalMux I__2119 (
            .O(N__16188),
            .I(\tok.A_stk.tail_23 ));
    LocalMux I__2118 (
            .O(N__16185),
            .I(\tok.A_stk.tail_23 ));
    InMux I__2117 (
            .O(N__16180),
            .I(N__16177));
    LocalMux I__2116 (
            .O(N__16177),
            .I(N__16174));
    Span4Mux_s3_v I__2115 (
            .O(N__16174),
            .I(N__16171));
    Odrv4 I__2114 (
            .O(N__16171),
            .I(\tok.table_rd_11 ));
    CascadeMux I__2113 (
            .O(N__16168),
            .I(\tok.n228_cascade_ ));
    CascadeMux I__2112 (
            .O(N__16165),
            .I(\tok.n203_adj_879_cascade_ ));
    InMux I__2111 (
            .O(N__16162),
            .I(N__16159));
    LocalMux I__2110 (
            .O(N__16159),
            .I(\tok.n228 ));
    CascadeMux I__2109 (
            .O(N__16156),
            .I(\tok.n212_adj_880_cascade_ ));
    InMux I__2108 (
            .O(N__16153),
            .I(N__16150));
    LocalMux I__2107 (
            .O(N__16150),
            .I(N__16147));
    Odrv4 I__2106 (
            .O(N__16147),
            .I(\tok.n6339 ));
    CascadeMux I__2105 (
            .O(N__16144),
            .I(\tok.n161_adj_692_cascade_ ));
    InMux I__2104 (
            .O(N__16141),
            .I(N__16138));
    LocalMux I__2103 (
            .O(N__16138),
            .I(N__16135));
    Odrv4 I__2102 (
            .O(N__16135),
            .I(\tok.n6356 ));
    InMux I__2101 (
            .O(N__16132),
            .I(N__16129));
    LocalMux I__2100 (
            .O(N__16129),
            .I(\tok.n6417 ));
    InMux I__2099 (
            .O(N__16126),
            .I(N__16123));
    LocalMux I__2098 (
            .O(N__16123),
            .I(\tok.n206_adj_881 ));
    InMux I__2097 (
            .O(N__16120),
            .I(N__16108));
    InMux I__2096 (
            .O(N__16119),
            .I(N__16108));
    InMux I__2095 (
            .O(N__16118),
            .I(N__16101));
    InMux I__2094 (
            .O(N__16117),
            .I(N__16101));
    InMux I__2093 (
            .O(N__16116),
            .I(N__16101));
    InMux I__2092 (
            .O(N__16115),
            .I(N__16094));
    InMux I__2091 (
            .O(N__16114),
            .I(N__16094));
    InMux I__2090 (
            .O(N__16113),
            .I(N__16094));
    LocalMux I__2089 (
            .O(N__16108),
            .I(\tok.n83 ));
    LocalMux I__2088 (
            .O(N__16101),
            .I(\tok.n83 ));
    LocalMux I__2087 (
            .O(N__16094),
            .I(\tok.n83 ));
    InMux I__2086 (
            .O(N__16087),
            .I(N__16084));
    LocalMux I__2085 (
            .O(N__16084),
            .I(N__16081));
    Span4Mux_v I__2084 (
            .O(N__16081),
            .I(N__16078));
    Odrv4 I__2083 (
            .O(N__16078),
            .I(\tok.n161_adj_836 ));
    CascadeMux I__2082 (
            .O(N__16075),
            .I(\tok.n197_adj_837_cascade_ ));
    InMux I__2081 (
            .O(N__16072),
            .I(N__16069));
    LocalMux I__2080 (
            .O(N__16069),
            .I(N__16066));
    Span4Mux_v I__2079 (
            .O(N__16066),
            .I(N__16063));
    Odrv4 I__2078 (
            .O(N__16063),
            .I(\tok.n248_adj_838 ));
    InMux I__2077 (
            .O(N__16060),
            .I(N__16057));
    LocalMux I__2076 (
            .O(N__16057),
            .I(N__16054));
    Span4Mux_v I__2075 (
            .O(N__16054),
            .I(N__16051));
    Odrv4 I__2074 (
            .O(N__16051),
            .I(\tok.n161_adj_650 ));
    CascadeMux I__2073 (
            .O(N__16048),
            .I(\tok.n6386_cascade_ ));
    CascadeMux I__2072 (
            .O(N__16045),
            .I(\tok.n197_adj_652_cascade_ ));
    InMux I__2071 (
            .O(N__16042),
            .I(\tok.n4807 ));
    InMux I__2070 (
            .O(N__16039),
            .I(\tok.n4808 ));
    CascadeMux I__2069 (
            .O(N__16036),
            .I(N__16033));
    InMux I__2068 (
            .O(N__16033),
            .I(N__16030));
    LocalMux I__2067 (
            .O(N__16030),
            .I(N__16027));
    Odrv12 I__2066 (
            .O(N__16027),
            .I(\tok.n6377 ));
    InMux I__2065 (
            .O(N__16024),
            .I(\tok.n4809 ));
    InMux I__2064 (
            .O(N__16021),
            .I(bfn_4_11_0_));
    InMux I__2063 (
            .O(N__16018),
            .I(\tok.n4811 ));
    InMux I__2062 (
            .O(N__16015),
            .I(N__16012));
    LocalMux I__2061 (
            .O(N__16012),
            .I(\tok.n6362 ));
    InMux I__2060 (
            .O(N__16009),
            .I(\tok.n4799 ));
    InMux I__2059 (
            .O(N__16006),
            .I(N__16003));
    LocalMux I__2058 (
            .O(N__16003),
            .I(\tok.n6556 ));
    InMux I__2057 (
            .O(N__16000),
            .I(\tok.n4800 ));
    InMux I__2056 (
            .O(N__15997),
            .I(\tok.n4801 ));
    InMux I__2055 (
            .O(N__15994),
            .I(\tok.n4802 ));
    InMux I__2054 (
            .O(N__15991),
            .I(bfn_4_10_0_));
    InMux I__2053 (
            .O(N__15988),
            .I(\tok.n4804 ));
    CascadeMux I__2052 (
            .O(N__15985),
            .I(N__15982));
    InMux I__2051 (
            .O(N__15982),
            .I(N__15979));
    LocalMux I__2050 (
            .O(N__15979),
            .I(N__15976));
    Odrv12 I__2049 (
            .O(N__15976),
            .I(\tok.n6437 ));
    InMux I__2048 (
            .O(N__15973),
            .I(\tok.n4805 ));
    InMux I__2047 (
            .O(N__15970),
            .I(\tok.n4806 ));
    CascadeMux I__2046 (
            .O(N__15967),
            .I(N__15964));
    InMux I__2045 (
            .O(N__15964),
            .I(N__15958));
    InMux I__2044 (
            .O(N__15963),
            .I(N__15958));
    LocalMux I__2043 (
            .O(N__15958),
            .I(\tok.key_rd_6 ));
    InMux I__2042 (
            .O(N__15955),
            .I(N__15949));
    InMux I__2041 (
            .O(N__15954),
            .I(N__15949));
    LocalMux I__2040 (
            .O(N__15949),
            .I(\tok.key_rd_0 ));
    InMux I__2039 (
            .O(N__15946),
            .I(N__15943));
    LocalMux I__2038 (
            .O(N__15943),
            .I(N__15940));
    Odrv4 I__2037 (
            .O(N__15940),
            .I(\tok.n25 ));
    CascadeMux I__2036 (
            .O(N__15937),
            .I(N__15934));
    InMux I__2035 (
            .O(N__15934),
            .I(N__15928));
    InMux I__2034 (
            .O(N__15933),
            .I(N__15928));
    LocalMux I__2033 (
            .O(N__15928),
            .I(\tok.key_rd_4 ));
    InMux I__2032 (
            .O(N__15925),
            .I(N__15919));
    InMux I__2031 (
            .O(N__15924),
            .I(N__15919));
    LocalMux I__2030 (
            .O(N__15919),
            .I(\tok.key_rd_1 ));
    InMux I__2029 (
            .O(N__15916),
            .I(N__15913));
    LocalMux I__2028 (
            .O(N__15913),
            .I(N__15910));
    Span4Mux_h I__2027 (
            .O(N__15910),
            .I(N__15907));
    Odrv4 I__2026 (
            .O(N__15907),
            .I(\tok.n18 ));
    CascadeMux I__2025 (
            .O(N__15904),
            .I(\tok.n6575_cascade_ ));
    InMux I__2024 (
            .O(N__15901),
            .I(N__15898));
    LocalMux I__2023 (
            .O(N__15898),
            .I(\tok.n177 ));
    InMux I__2022 (
            .O(N__15895),
            .I(\tok.n4797 ));
    InMux I__2021 (
            .O(N__15892),
            .I(\tok.n4798 ));
    InMux I__2020 (
            .O(N__15889),
            .I(N__15886));
    LocalMux I__2019 (
            .O(N__15886),
            .I(N__15883));
    Odrv4 I__2018 (
            .O(N__15883),
            .I(\tok.n33 ));
    InMux I__2017 (
            .O(N__15880),
            .I(N__15877));
    LocalMux I__2016 (
            .O(N__15877),
            .I(\tok.n27_adj_707 ));
    InMux I__2015 (
            .O(N__15874),
            .I(N__15871));
    LocalMux I__2014 (
            .O(N__15871),
            .I(N__15868));
    Odrv12 I__2013 (
            .O(N__15868),
            .I(\tok.n33_adj_663 ));
    CascadeMux I__2012 (
            .O(N__15865),
            .I(\tok.n27_adj_708_cascade_ ));
    CascadeMux I__2011 (
            .O(N__15862),
            .I(N__15858));
    CascadeMux I__2010 (
            .O(N__15861),
            .I(N__15855));
    CascadeBuf I__2009 (
            .O(N__15858),
            .I(N__15852));
    CascadeBuf I__2008 (
            .O(N__15855),
            .I(N__15849));
    CascadeMux I__2007 (
            .O(N__15852),
            .I(N__15846));
    CascadeMux I__2006 (
            .O(N__15849),
            .I(N__15841));
    InMux I__2005 (
            .O(N__15846),
            .I(N__15837));
    InMux I__2004 (
            .O(N__15845),
            .I(N__15834));
    InMux I__2003 (
            .O(N__15844),
            .I(N__15831));
    InMux I__2002 (
            .O(N__15841),
            .I(N__15828));
    InMux I__2001 (
            .O(N__15840),
            .I(N__15825));
    LocalMux I__2000 (
            .O(N__15837),
            .I(N__15822));
    LocalMux I__1999 (
            .O(N__15834),
            .I(N__15817));
    LocalMux I__1998 (
            .O(N__15831),
            .I(N__15817));
    LocalMux I__1997 (
            .O(N__15828),
            .I(N__15814));
    LocalMux I__1996 (
            .O(N__15825),
            .I(N__15809));
    Span4Mux_h I__1995 (
            .O(N__15822),
            .I(N__15809));
    Odrv4 I__1994 (
            .O(N__15817),
            .I(\tok.n29 ));
    Odrv4 I__1993 (
            .O(N__15814),
            .I(\tok.n29 ));
    Odrv4 I__1992 (
            .O(N__15809),
            .I(\tok.n29 ));
    CascadeMux I__1991 (
            .O(N__15802),
            .I(N__15798));
    InMux I__1990 (
            .O(N__15801),
            .I(N__15789));
    InMux I__1989 (
            .O(N__15798),
            .I(N__15789));
    InMux I__1988 (
            .O(N__15797),
            .I(N__15789));
    CascadeMux I__1987 (
            .O(N__15796),
            .I(N__15784));
    LocalMux I__1986 (
            .O(N__15789),
            .I(N__15780));
    InMux I__1985 (
            .O(N__15788),
            .I(N__15773));
    InMux I__1984 (
            .O(N__15787),
            .I(N__15773));
    InMux I__1983 (
            .O(N__15784),
            .I(N__15773));
    CascadeMux I__1982 (
            .O(N__15783),
            .I(N__15768));
    Span4Mux_h I__1981 (
            .O(N__15780),
            .I(N__15763));
    LocalMux I__1980 (
            .O(N__15773),
            .I(N__15760));
    InMux I__1979 (
            .O(N__15772),
            .I(N__15749));
    InMux I__1978 (
            .O(N__15771),
            .I(N__15749));
    InMux I__1977 (
            .O(N__15768),
            .I(N__15749));
    InMux I__1976 (
            .O(N__15767),
            .I(N__15749));
    InMux I__1975 (
            .O(N__15766),
            .I(N__15749));
    Odrv4 I__1974 (
            .O(N__15763),
            .I(\tok.search_clk ));
    Odrv4 I__1973 (
            .O(N__15760),
            .I(\tok.search_clk ));
    LocalMux I__1972 (
            .O(N__15749),
            .I(\tok.search_clk ));
    CascadeMux I__1971 (
            .O(N__15742),
            .I(N__15736));
    CascadeMux I__1970 (
            .O(N__15741),
            .I(N__15733));
    CascadeMux I__1969 (
            .O(N__15740),
            .I(N__15730));
    CascadeMux I__1968 (
            .O(N__15739),
            .I(N__15727));
    InMux I__1967 (
            .O(N__15736),
            .I(N__15714));
    InMux I__1966 (
            .O(N__15733),
            .I(N__15714));
    InMux I__1965 (
            .O(N__15730),
            .I(N__15714));
    InMux I__1964 (
            .O(N__15727),
            .I(N__15714));
    CascadeMux I__1963 (
            .O(N__15726),
            .I(N__15710));
    CascadeMux I__1962 (
            .O(N__15725),
            .I(N__15707));
    CascadeMux I__1961 (
            .O(N__15724),
            .I(N__15704));
    CascadeMux I__1960 (
            .O(N__15723),
            .I(N__15701));
    LocalMux I__1959 (
            .O(N__15714),
            .I(N__15698));
    InMux I__1958 (
            .O(N__15713),
            .I(N__15695));
    InMux I__1957 (
            .O(N__15710),
            .I(N__15686));
    InMux I__1956 (
            .O(N__15707),
            .I(N__15686));
    InMux I__1955 (
            .O(N__15704),
            .I(N__15686));
    InMux I__1954 (
            .O(N__15701),
            .I(N__15686));
    Span4Mux_s2_h I__1953 (
            .O(N__15698),
            .I(N__15681));
    LocalMux I__1952 (
            .O(N__15695),
            .I(N__15681));
    LocalMux I__1951 (
            .O(N__15686),
            .I(\tok.found_slot ));
    Odrv4 I__1950 (
            .O(N__15681),
            .I(\tok.found_slot ));
    InMux I__1949 (
            .O(N__15676),
            .I(N__15673));
    LocalMux I__1948 (
            .O(N__15673),
            .I(N__15670));
    Span4Mux_v I__1947 (
            .O(N__15670),
            .I(N__15667));
    Span4Mux_s2_h I__1946 (
            .O(N__15667),
            .I(N__15664));
    Odrv4 I__1945 (
            .O(N__15664),
            .I(\tok.n6670 ));
    InMux I__1944 (
            .O(N__15661),
            .I(N__15658));
    LocalMux I__1943 (
            .O(N__15658),
            .I(N__15655));
    Span4Mux_h I__1942 (
            .O(N__15655),
            .I(N__15652));
    Odrv4 I__1941 (
            .O(N__15652),
            .I(\tok.n33_adj_633 ));
    CascadeMux I__1940 (
            .O(N__15649),
            .I(\tok.n27_adj_704_cascade_ ));
    CascadeMux I__1939 (
            .O(N__15646),
            .I(N__15642));
    CascadeMux I__1938 (
            .O(N__15645),
            .I(N__15639));
    CascadeBuf I__1937 (
            .O(N__15642),
            .I(N__15636));
    CascadeBuf I__1936 (
            .O(N__15639),
            .I(N__15633));
    CascadeMux I__1935 (
            .O(N__15636),
            .I(N__15628));
    CascadeMux I__1934 (
            .O(N__15633),
            .I(N__15625));
    InMux I__1933 (
            .O(N__15632),
            .I(N__15622));
    InMux I__1932 (
            .O(N__15631),
            .I(N__15619));
    InMux I__1931 (
            .O(N__15628),
            .I(N__15616));
    InMux I__1930 (
            .O(N__15625),
            .I(N__15613));
    LocalMux I__1929 (
            .O(N__15622),
            .I(N__15608));
    LocalMux I__1928 (
            .O(N__15619),
            .I(N__15608));
    LocalMux I__1927 (
            .O(N__15616),
            .I(N__15603));
    LocalMux I__1926 (
            .O(N__15613),
            .I(N__15603));
    Span4Mux_h I__1925 (
            .O(N__15608),
            .I(N__15599));
    Span4Mux_v I__1924 (
            .O(N__15603),
            .I(N__15596));
    InMux I__1923 (
            .O(N__15602),
            .I(N__15593));
    Span4Mux_h I__1922 (
            .O(N__15599),
            .I(N__15590));
    Span4Mux_s3_h I__1921 (
            .O(N__15596),
            .I(N__15587));
    LocalMux I__1920 (
            .O(N__15593),
            .I(\tok.n38 ));
    Odrv4 I__1919 (
            .O(N__15590),
            .I(\tok.n38 ));
    Odrv4 I__1918 (
            .O(N__15587),
            .I(\tok.n38 ));
    InMux I__1917 (
            .O(N__15580),
            .I(N__15577));
    LocalMux I__1916 (
            .O(N__15577),
            .I(N__15574));
    Span4Mux_v I__1915 (
            .O(N__15574),
            .I(N__15571));
    Odrv4 I__1914 (
            .O(N__15571),
            .I(\tok.n33_adj_632 ));
    CascadeMux I__1913 (
            .O(N__15568),
            .I(N__15565));
    InMux I__1912 (
            .O(N__15565),
            .I(N__15562));
    LocalMux I__1911 (
            .O(N__15562),
            .I(N__15559));
    Span4Mux_h I__1910 (
            .O(N__15559),
            .I(N__15556));
    Odrv4 I__1909 (
            .O(N__15556),
            .I(\tok.n33_adj_661 ));
    CascadeMux I__1908 (
            .O(N__15553),
            .I(\tok.n27_adj_705_cascade_ ));
    CascadeMux I__1907 (
            .O(N__15550),
            .I(N__15546));
    CascadeMux I__1906 (
            .O(N__15549),
            .I(N__15543));
    CascadeBuf I__1905 (
            .O(N__15546),
            .I(N__15539));
    CascadeBuf I__1904 (
            .O(N__15543),
            .I(N__15536));
    InMux I__1903 (
            .O(N__15542),
            .I(N__15533));
    CascadeMux I__1902 (
            .O(N__15539),
            .I(N__15529));
    CascadeMux I__1901 (
            .O(N__15536),
            .I(N__15526));
    LocalMux I__1900 (
            .O(N__15533),
            .I(N__15523));
    InMux I__1899 (
            .O(N__15532),
            .I(N__15520));
    InMux I__1898 (
            .O(N__15529),
            .I(N__15517));
    InMux I__1897 (
            .O(N__15526),
            .I(N__15514));
    Span4Mux_v I__1896 (
            .O(N__15523),
            .I(N__15510));
    LocalMux I__1895 (
            .O(N__15520),
            .I(N__15507));
    LocalMux I__1894 (
            .O(N__15517),
            .I(N__15502));
    LocalMux I__1893 (
            .O(N__15514),
            .I(N__15502));
    InMux I__1892 (
            .O(N__15513),
            .I(N__15499));
    Span4Mux_s1_h I__1891 (
            .O(N__15510),
            .I(N__15494));
    Span4Mux_v I__1890 (
            .O(N__15507),
            .I(N__15494));
    Span4Mux_v I__1889 (
            .O(N__15502),
            .I(N__15491));
    LocalMux I__1888 (
            .O(N__15499),
            .I(\tok.n36 ));
    Odrv4 I__1887 (
            .O(N__15494),
            .I(\tok.n36 ));
    Odrv4 I__1886 (
            .O(N__15491),
            .I(\tok.n36 ));
    InMux I__1885 (
            .O(N__15484),
            .I(N__15481));
    LocalMux I__1884 (
            .O(N__15481),
            .I(\tok.n27_adj_703 ));
    CascadeMux I__1883 (
            .O(N__15478),
            .I(N__15474));
    CascadeMux I__1882 (
            .O(N__15477),
            .I(N__15471));
    CascadeBuf I__1881 (
            .O(N__15474),
            .I(N__15468));
    CascadeBuf I__1880 (
            .O(N__15471),
            .I(N__15465));
    CascadeMux I__1879 (
            .O(N__15468),
            .I(N__15462));
    CascadeMux I__1878 (
            .O(N__15465),
            .I(N__15457));
    InMux I__1877 (
            .O(N__15462),
            .I(N__15454));
    InMux I__1876 (
            .O(N__15461),
            .I(N__15451));
    InMux I__1875 (
            .O(N__15460),
            .I(N__15448));
    InMux I__1874 (
            .O(N__15457),
            .I(N__15445));
    LocalMux I__1873 (
            .O(N__15454),
            .I(N__15442));
    LocalMux I__1872 (
            .O(N__15451),
            .I(N__15436));
    LocalMux I__1871 (
            .O(N__15448),
            .I(N__15436));
    LocalMux I__1870 (
            .O(N__15445),
            .I(N__15433));
    Span4Mux_h I__1869 (
            .O(N__15442),
            .I(N__15430));
    InMux I__1868 (
            .O(N__15441),
            .I(N__15427));
    Span4Mux_h I__1867 (
            .O(N__15436),
            .I(N__15424));
    Span4Mux_v I__1866 (
            .O(N__15433),
            .I(N__15419));
    Span4Mux_v I__1865 (
            .O(N__15430),
            .I(N__15419));
    LocalMux I__1864 (
            .O(N__15427),
            .I(\tok.n40 ));
    Odrv4 I__1863 (
            .O(N__15424),
            .I(\tok.n40 ));
    Odrv4 I__1862 (
            .O(N__15419),
            .I(\tok.n40 ));
    CascadeMux I__1861 (
            .O(N__15412),
            .I(N__15408));
    CascadeMux I__1860 (
            .O(N__15411),
            .I(N__15405));
    CascadeBuf I__1859 (
            .O(N__15408),
            .I(N__15402));
    CascadeBuf I__1858 (
            .O(N__15405),
            .I(N__15399));
    CascadeMux I__1857 (
            .O(N__15402),
            .I(N__15394));
    CascadeMux I__1856 (
            .O(N__15399),
            .I(N__15391));
    InMux I__1855 (
            .O(N__15398),
            .I(N__15388));
    InMux I__1854 (
            .O(N__15397),
            .I(N__15385));
    InMux I__1853 (
            .O(N__15394),
            .I(N__15382));
    InMux I__1852 (
            .O(N__15391),
            .I(N__15379));
    LocalMux I__1851 (
            .O(N__15388),
            .I(N__15373));
    LocalMux I__1850 (
            .O(N__15385),
            .I(N__15373));
    LocalMux I__1849 (
            .O(N__15382),
            .I(N__15368));
    LocalMux I__1848 (
            .O(N__15379),
            .I(N__15368));
    InMux I__1847 (
            .O(N__15378),
            .I(N__15365));
    Span12Mux_s8_v I__1846 (
            .O(N__15373),
            .I(N__15362));
    Sp12to4 I__1845 (
            .O(N__15368),
            .I(N__15359));
    LocalMux I__1844 (
            .O(N__15365),
            .I(\tok.n32 ));
    Odrv12 I__1843 (
            .O(N__15362),
            .I(\tok.n32 ));
    Odrv12 I__1842 (
            .O(N__15359),
            .I(\tok.n32 ));
    InMux I__1841 (
            .O(N__15352),
            .I(N__15346));
    InMux I__1840 (
            .O(N__15351),
            .I(N__15346));
    LocalMux I__1839 (
            .O(N__15346),
            .I(\tok.A_stk.tail_19 ));
    CascadeMux I__1838 (
            .O(N__15343),
            .I(N__15340));
    InMux I__1837 (
            .O(N__15340),
            .I(N__15334));
    InMux I__1836 (
            .O(N__15339),
            .I(N__15334));
    LocalMux I__1835 (
            .O(N__15334),
            .I(\tok.A_stk.tail_3 ));
    CascadeMux I__1834 (
            .O(N__15331),
            .I(\tok.n4_cascade_ ));
    InMux I__1833 (
            .O(N__15328),
            .I(N__15325));
    LocalMux I__1832 (
            .O(N__15325),
            .I(N__15322));
    Odrv4 I__1831 (
            .O(N__15322),
            .I(\tok.n6273 ));
    InMux I__1830 (
            .O(N__15319),
            .I(N__15316));
    LocalMux I__1829 (
            .O(N__15316),
            .I(N__15313));
    Span4Mux_v I__1828 (
            .O(N__15313),
            .I(N__15310));
    Odrv4 I__1827 (
            .O(N__15310),
            .I(\tok.table_wr_data_9 ));
    CascadeMux I__1826 (
            .O(N__15307),
            .I(N__15304));
    InMux I__1825 (
            .O(N__15304),
            .I(N__15301));
    LocalMux I__1824 (
            .O(N__15301),
            .I(\tok.n4 ));
    InMux I__1823 (
            .O(N__15298),
            .I(N__15295));
    LocalMux I__1822 (
            .O(N__15295),
            .I(N__15292));
    Odrv4 I__1821 (
            .O(N__15292),
            .I(\tok.n6252 ));
    CascadeMux I__1820 (
            .O(N__15289),
            .I(\tok.n6253_cascade_ ));
    InMux I__1819 (
            .O(N__15286),
            .I(N__15282));
    InMux I__1818 (
            .O(N__15285),
            .I(N__15279));
    LocalMux I__1817 (
            .O(N__15282),
            .I(tail_99));
    LocalMux I__1816 (
            .O(N__15279),
            .I(tail_99));
    CascadeMux I__1815 (
            .O(N__15274),
            .I(N__15270));
    InMux I__1814 (
            .O(N__15273),
            .I(N__15267));
    InMux I__1813 (
            .O(N__15270),
            .I(N__15264));
    LocalMux I__1812 (
            .O(N__15267),
            .I(tail_115));
    LocalMux I__1811 (
            .O(N__15264),
            .I(tail_115));
    InMux I__1810 (
            .O(N__15259),
            .I(N__15255));
    InMux I__1809 (
            .O(N__15258),
            .I(N__15252));
    LocalMux I__1808 (
            .O(N__15255),
            .I(\tok.A_stk.tail_92 ));
    LocalMux I__1807 (
            .O(N__15252),
            .I(\tok.A_stk.tail_92 ));
    InMux I__1806 (
            .O(N__15247),
            .I(N__15241));
    InMux I__1805 (
            .O(N__15246),
            .I(N__15241));
    LocalMux I__1804 (
            .O(N__15241),
            .I(\tok.A_stk.tail_60 ));
    InMux I__1803 (
            .O(N__15238),
            .I(N__15234));
    InMux I__1802 (
            .O(N__15237),
            .I(N__15231));
    LocalMux I__1801 (
            .O(N__15234),
            .I(\tok.A_stk.tail_76 ));
    LocalMux I__1800 (
            .O(N__15231),
            .I(\tok.A_stk.tail_76 ));
    InMux I__1799 (
            .O(N__15226),
            .I(N__15222));
    InMux I__1798 (
            .O(N__15225),
            .I(N__15219));
    LocalMux I__1797 (
            .O(N__15222),
            .I(\tok.A_stk.tail_6 ));
    LocalMux I__1796 (
            .O(N__15219),
            .I(\tok.A_stk.tail_6 ));
    InMux I__1795 (
            .O(N__15214),
            .I(N__15210));
    InMux I__1794 (
            .O(N__15213),
            .I(N__15207));
    LocalMux I__1793 (
            .O(N__15210),
            .I(\tok.A_stk.tail_12 ));
    LocalMux I__1792 (
            .O(N__15207),
            .I(\tok.A_stk.tail_12 ));
    InMux I__1791 (
            .O(N__15202),
            .I(N__15198));
    InMux I__1790 (
            .O(N__15201),
            .I(N__15195));
    LocalMux I__1789 (
            .O(N__15198),
            .I(N__15192));
    LocalMux I__1788 (
            .O(N__15195),
            .I(N__15189));
    Span4Mux_v I__1787 (
            .O(N__15192),
            .I(N__15184));
    Span4Mux_h I__1786 (
            .O(N__15189),
            .I(N__15184));
    Odrv4 I__1785 (
            .O(N__15184),
            .I(\tok.A_stk.tail_10 ));
    InMux I__1784 (
            .O(N__15181),
            .I(N__15175));
    InMux I__1783 (
            .O(N__15180),
            .I(N__15175));
    LocalMux I__1782 (
            .O(N__15175),
            .I(\tok.A_stk.tail_83 ));
    InMux I__1781 (
            .O(N__15172),
            .I(N__15166));
    InMux I__1780 (
            .O(N__15171),
            .I(N__15166));
    LocalMux I__1779 (
            .O(N__15166),
            .I(\tok.A_stk.tail_67 ));
    InMux I__1778 (
            .O(N__15163),
            .I(N__15157));
    InMux I__1777 (
            .O(N__15162),
            .I(N__15157));
    LocalMux I__1776 (
            .O(N__15157),
            .I(\tok.A_stk.tail_51 ));
    InMux I__1775 (
            .O(N__15154),
            .I(N__15148));
    InMux I__1774 (
            .O(N__15153),
            .I(N__15148));
    LocalMux I__1773 (
            .O(N__15148),
            .I(\tok.A_stk.tail_35 ));
    InMux I__1772 (
            .O(N__15145),
            .I(N__15139));
    InMux I__1771 (
            .O(N__15144),
            .I(N__15139));
    LocalMux I__1770 (
            .O(N__15139),
            .I(\tok.A_stk.tail_70 ));
    InMux I__1769 (
            .O(N__15136),
            .I(N__15130));
    InMux I__1768 (
            .O(N__15135),
            .I(N__15130));
    LocalMux I__1767 (
            .O(N__15130),
            .I(\tok.A_stk.tail_54 ));
    InMux I__1766 (
            .O(N__15127),
            .I(N__15121));
    InMux I__1765 (
            .O(N__15126),
            .I(N__15121));
    LocalMux I__1764 (
            .O(N__15121),
            .I(\tok.A_stk.tail_38 ));
    InMux I__1763 (
            .O(N__15118),
            .I(N__15114));
    InMux I__1762 (
            .O(N__15117),
            .I(N__15111));
    LocalMux I__1761 (
            .O(N__15114),
            .I(\tok.A_stk.tail_22 ));
    LocalMux I__1760 (
            .O(N__15111),
            .I(\tok.A_stk.tail_22 ));
    InMux I__1759 (
            .O(N__15106),
            .I(N__15100));
    InMux I__1758 (
            .O(N__15105),
            .I(N__15100));
    LocalMux I__1757 (
            .O(N__15100),
            .I(\tok.A_stk.tail_28 ));
    InMux I__1756 (
            .O(N__15097),
            .I(N__15091));
    InMux I__1755 (
            .O(N__15096),
            .I(N__15091));
    LocalMux I__1754 (
            .O(N__15091),
            .I(\tok.A_stk.tail_44 ));
    InMux I__1753 (
            .O(N__15088),
            .I(N__15082));
    InMux I__1752 (
            .O(N__15087),
            .I(N__15082));
    LocalMux I__1751 (
            .O(N__15082),
            .I(\tok.A_stk.tail_65 ));
    InMux I__1750 (
            .O(N__15079),
            .I(N__15073));
    InMux I__1749 (
            .O(N__15078),
            .I(N__15073));
    LocalMux I__1748 (
            .O(N__15073),
            .I(tail_49));
    InMux I__1747 (
            .O(N__15070),
            .I(N__15064));
    InMux I__1746 (
            .O(N__15069),
            .I(N__15064));
    LocalMux I__1745 (
            .O(N__15064),
            .I(tail_81));
    InMux I__1744 (
            .O(N__15061),
            .I(N__15055));
    InMux I__1743 (
            .O(N__15060),
            .I(N__15055));
    LocalMux I__1742 (
            .O(N__15055),
            .I(\tok.A_stk.tail_33 ));
    CascadeMux I__1741 (
            .O(N__15052),
            .I(N__15049));
    InMux I__1740 (
            .O(N__15049),
            .I(N__15043));
    InMux I__1739 (
            .O(N__15048),
            .I(N__15043));
    LocalMux I__1738 (
            .O(N__15043),
            .I(tail_17));
    InMux I__1737 (
            .O(N__15040),
            .I(N__15034));
    InMux I__1736 (
            .O(N__15039),
            .I(N__15034));
    LocalMux I__1735 (
            .O(N__15034),
            .I(\tok.A_stk.tail_1 ));
    InMux I__1734 (
            .O(N__15031),
            .I(N__15027));
    InMux I__1733 (
            .O(N__15030),
            .I(N__15024));
    LocalMux I__1732 (
            .O(N__15027),
            .I(N__15021));
    LocalMux I__1731 (
            .O(N__15024),
            .I(tail_102));
    Odrv12 I__1730 (
            .O(N__15021),
            .I(tail_102));
    InMux I__1729 (
            .O(N__15016),
            .I(N__15012));
    InMux I__1728 (
            .O(N__15015),
            .I(N__15009));
    LocalMux I__1727 (
            .O(N__15012),
            .I(N__15006));
    LocalMux I__1726 (
            .O(N__15009),
            .I(\tok.A_stk.tail_86 ));
    Odrv12 I__1725 (
            .O(N__15006),
            .I(\tok.A_stk.tail_86 ));
    CascadeMux I__1724 (
            .O(N__15001),
            .I(\tok.n281_cascade_ ));
    CascadeMux I__1723 (
            .O(N__14998),
            .I(\tok.n236_adj_864_cascade_ ));
    CascadeMux I__1722 (
            .O(N__14995),
            .I(\tok.n2648_cascade_ ));
    InMux I__1721 (
            .O(N__14992),
            .I(N__14989));
    LocalMux I__1720 (
            .O(N__14989),
            .I(\tok.n226_adj_865 ));
    InMux I__1719 (
            .O(N__14986),
            .I(N__14983));
    LocalMux I__1718 (
            .O(N__14983),
            .I(\tok.n6334 ));
    InMux I__1717 (
            .O(N__14980),
            .I(N__14977));
    LocalMux I__1716 (
            .O(N__14977),
            .I(\tok.n4_adj_762 ));
    InMux I__1715 (
            .O(N__14974),
            .I(N__14971));
    LocalMux I__1714 (
            .O(N__14971),
            .I(\tok.n6316 ));
    InMux I__1713 (
            .O(N__14968),
            .I(N__14965));
    LocalMux I__1712 (
            .O(N__14965),
            .I(N__14961));
    InMux I__1711 (
            .O(N__14964),
            .I(N__14958));
    Odrv4 I__1710 (
            .O(N__14961),
            .I(sender_1));
    LocalMux I__1709 (
            .O(N__14958),
            .I(sender_1));
    IoInMux I__1708 (
            .O(N__14953),
            .I(N__14950));
    LocalMux I__1707 (
            .O(N__14950),
            .I(N__14947));
    Span4Mux_s0_v I__1706 (
            .O(N__14947),
            .I(N__14944));
    Odrv4 I__1705 (
            .O(N__14944),
            .I(tx_c));
    InMux I__1704 (
            .O(N__14941),
            .I(N__14938));
    LocalMux I__1703 (
            .O(N__14938),
            .I(N__14935));
    Span4Mux_v I__1702 (
            .O(N__14935),
            .I(N__14932));
    Odrv4 I__1701 (
            .O(N__14932),
            .I(\tok.table_rd_14 ));
    CascadeMux I__1700 (
            .O(N__14929),
            .I(\tok.n225_cascade_ ));
    CascadeMux I__1699 (
            .O(N__14926),
            .I(\tok.n203_adj_664_cascade_ ));
    InMux I__1698 (
            .O(N__14923),
            .I(N__14920));
    LocalMux I__1697 (
            .O(N__14920),
            .I(\tok.n225 ));
    InMux I__1696 (
            .O(N__14917),
            .I(N__14914));
    LocalMux I__1695 (
            .O(N__14914),
            .I(\tok.n224 ));
    InMux I__1694 (
            .O(N__14911),
            .I(N__14908));
    LocalMux I__1693 (
            .O(N__14908),
            .I(N__14905));
    Span4Mux_s3_v I__1692 (
            .O(N__14905),
            .I(N__14902));
    Odrv4 I__1691 (
            .O(N__14902),
            .I(\tok.table_rd_15 ));
    CascadeMux I__1690 (
            .O(N__14899),
            .I(\tok.n224_cascade_ ));
    InMux I__1689 (
            .O(N__14896),
            .I(N__14893));
    LocalMux I__1688 (
            .O(N__14893),
            .I(\tok.n203_adj_688 ));
    CascadeMux I__1687 (
            .O(N__14890),
            .I(\tok.n6373_cascade_ ));
    CascadeMux I__1686 (
            .O(N__14887),
            .I(\tok.n206_adj_666_cascade_ ));
    InMux I__1685 (
            .O(N__14884),
            .I(N__14881));
    LocalMux I__1684 (
            .O(N__14881),
            .I(\tok.n212_adj_665 ));
    InMux I__1683 (
            .O(N__14878),
            .I(\tok.n4779 ));
    InMux I__1682 (
            .O(N__14875),
            .I(\tok.n4780 ));
    InMux I__1681 (
            .O(N__14872),
            .I(bfn_2_11_0_));
    CascadeMux I__1680 (
            .O(N__14869),
            .I(\tok.n214_cascade_ ));
    InMux I__1679 (
            .O(N__14866),
            .I(N__14863));
    LocalMux I__1678 (
            .O(N__14863),
            .I(N__14860));
    Span4Mux_v I__1677 (
            .O(N__14860),
            .I(N__14857));
    Odrv4 I__1676 (
            .O(N__14857),
            .I(\tok.n6358 ));
    InMux I__1675 (
            .O(N__14854),
            .I(N__14851));
    LocalMux I__1674 (
            .O(N__14851),
            .I(N__14848));
    Odrv4 I__1673 (
            .O(N__14848),
            .I(\tok.n6402 ));
    InMux I__1672 (
            .O(N__14845),
            .I(N__14842));
    LocalMux I__1671 (
            .O(N__14842),
            .I(N__14839));
    Odrv4 I__1670 (
            .O(N__14839),
            .I(\tok.table_rd_12 ));
    InMux I__1669 (
            .O(N__14836),
            .I(N__14830));
    InMux I__1668 (
            .O(N__14835),
            .I(N__14830));
    LocalMux I__1667 (
            .O(N__14830),
            .I(\tok.n227 ));
    CascadeMux I__1666 (
            .O(N__14827),
            .I(\tok.n203_cascade_ ));
    CascadeMux I__1665 (
            .O(N__14824),
            .I(\tok.n212_cascade_ ));
    InMux I__1664 (
            .O(N__14821),
            .I(N__14818));
    LocalMux I__1663 (
            .O(N__14818),
            .I(\tok.n206 ));
    InMux I__1662 (
            .O(N__14815),
            .I(\tok.n4774 ));
    InMux I__1661 (
            .O(N__14812),
            .I(\tok.n4775 ));
    InMux I__1660 (
            .O(N__14809),
            .I(\tok.n4776 ));
    InMux I__1659 (
            .O(N__14806),
            .I(\tok.n4777 ));
    InMux I__1658 (
            .O(N__14803),
            .I(\tok.n4778 ));
    InMux I__1657 (
            .O(N__14800),
            .I(N__14794));
    InMux I__1656 (
            .O(N__14799),
            .I(N__14794));
    LocalMux I__1655 (
            .O(N__14794),
            .I(\tok.key_rd_10 ));
    CascadeMux I__1654 (
            .O(N__14791),
            .I(N__14787));
    CascadeMux I__1653 (
            .O(N__14790),
            .I(N__14784));
    InMux I__1652 (
            .O(N__14787),
            .I(N__14779));
    InMux I__1651 (
            .O(N__14784),
            .I(N__14779));
    LocalMux I__1650 (
            .O(N__14779),
            .I(\tok.key_rd_12 ));
    InMux I__1649 (
            .O(N__14776),
            .I(N__14773));
    LocalMux I__1648 (
            .O(N__14773),
            .I(\tok.n26 ));
    CascadeMux I__1647 (
            .O(N__14770),
            .I(\tok.n27_adj_639_cascade_ ));
    InMux I__1646 (
            .O(N__14767),
            .I(N__14764));
    LocalMux I__1645 (
            .O(N__14764),
            .I(\tok.found_slot_N_144 ));
    InMux I__1644 (
            .O(N__14761),
            .I(N__14758));
    LocalMux I__1643 (
            .O(N__14758),
            .I(\tok.n6322 ));
    CascadeMux I__1642 (
            .O(N__14755),
            .I(\tok.n313_cascade_ ));
    InMux I__1641 (
            .O(N__14752),
            .I(N__14748));
    InMux I__1640 (
            .O(N__14751),
            .I(N__14745));
    LocalMux I__1639 (
            .O(N__14748),
            .I(\tok.key_rd_2 ));
    LocalMux I__1638 (
            .O(N__14745),
            .I(\tok.key_rd_2 ));
    CascadeMux I__1637 (
            .O(N__14740),
            .I(N__14736));
    InMux I__1636 (
            .O(N__14739),
            .I(N__14733));
    InMux I__1635 (
            .O(N__14736),
            .I(N__14730));
    LocalMux I__1634 (
            .O(N__14733),
            .I(\tok.key_rd_7 ));
    LocalMux I__1633 (
            .O(N__14730),
            .I(\tok.key_rd_7 ));
    InMux I__1632 (
            .O(N__14725),
            .I(N__14722));
    LocalMux I__1631 (
            .O(N__14722),
            .I(\tok.n22 ));
    InMux I__1630 (
            .O(N__14719),
            .I(N__14716));
    LocalMux I__1629 (
            .O(N__14716),
            .I(\tok.n33_adj_634 ));
    CascadeMux I__1628 (
            .O(N__14713),
            .I(\tok.n27_adj_706_cascade_ ));
    CascadeMux I__1627 (
            .O(N__14710),
            .I(N__14706));
    CascadeMux I__1626 (
            .O(N__14709),
            .I(N__14703));
    CascadeBuf I__1625 (
            .O(N__14706),
            .I(N__14700));
    CascadeBuf I__1624 (
            .O(N__14703),
            .I(N__14697));
    CascadeMux I__1623 (
            .O(N__14700),
            .I(N__14694));
    CascadeMux I__1622 (
            .O(N__14697),
            .I(N__14691));
    InMux I__1621 (
            .O(N__14694),
            .I(N__14688));
    InMux I__1620 (
            .O(N__14691),
            .I(N__14685));
    LocalMux I__1619 (
            .O(N__14688),
            .I(N__14677));
    LocalMux I__1618 (
            .O(N__14685),
            .I(N__14677));
    InMux I__1617 (
            .O(N__14684),
            .I(N__14674));
    InMux I__1616 (
            .O(N__14683),
            .I(N__14671));
    InMux I__1615 (
            .O(N__14682),
            .I(N__14668));
    Span12Mux_s8_v I__1614 (
            .O(N__14677),
            .I(N__14665));
    LocalMux I__1613 (
            .O(N__14674),
            .I(\tok.n35 ));
    LocalMux I__1612 (
            .O(N__14671),
            .I(\tok.n35 ));
    LocalMux I__1611 (
            .O(N__14668),
            .I(\tok.n35 ));
    Odrv12 I__1610 (
            .O(N__14665),
            .I(\tok.n35 ));
    CascadeMux I__1609 (
            .O(N__14656),
            .I(\tok.n6667_cascade_ ));
    InMux I__1608 (
            .O(N__14653),
            .I(N__14650));
    LocalMux I__1607 (
            .O(N__14650),
            .I(N__14647));
    Odrv4 I__1606 (
            .O(N__14647),
            .I(\tok.n2532 ));
    InMux I__1605 (
            .O(N__14644),
            .I(N__14641));
    LocalMux I__1604 (
            .O(N__14641),
            .I(N__14638));
    Odrv4 I__1603 (
            .O(N__14638),
            .I(\tok.n4_adj_642 ));
    CascadeMux I__1602 (
            .O(N__14635),
            .I(\tok.found_slot_cascade_ ));
    SRMux I__1601 (
            .O(N__14632),
            .I(N__14628));
    SRMux I__1600 (
            .O(N__14631),
            .I(N__14625));
    LocalMux I__1599 (
            .O(N__14628),
            .I(N__14622));
    LocalMux I__1598 (
            .O(N__14625),
            .I(N__14619));
    Span4Mux_h I__1597 (
            .O(N__14622),
            .I(N__14616));
    Span4Mux_h I__1596 (
            .O(N__14619),
            .I(N__14613));
    Span4Mux_s2_h I__1595 (
            .O(N__14616),
            .I(N__14610));
    Odrv4 I__1594 (
            .O(N__14613),
            .I(\tok.write_slot ));
    Odrv4 I__1593 (
            .O(N__14610),
            .I(\tok.write_slot ));
    CascadeMux I__1592 (
            .O(N__14605),
            .I(\tok.n21_cascade_ ));
    CascadeMux I__1591 (
            .O(N__14602),
            .I(N__14599));
    InMux I__1590 (
            .O(N__14599),
            .I(N__14596));
    LocalMux I__1589 (
            .O(N__14596),
            .I(\tok.n30_adj_647 ));
    CascadeMux I__1588 (
            .O(N__14593),
            .I(\tok.n4_adj_642_cascade_ ));
    InMux I__1587 (
            .O(N__14590),
            .I(N__14587));
    LocalMux I__1586 (
            .O(N__14587),
            .I(N__14584));
    Span4Mux_v I__1585 (
            .O(N__14584),
            .I(N__14581));
    Odrv4 I__1584 (
            .O(N__14581),
            .I(\tok.table_wr_data_13 ));
    InMux I__1583 (
            .O(N__14578),
            .I(N__14575));
    LocalMux I__1582 (
            .O(N__14575),
            .I(N__14572));
    Span4Mux_h I__1581 (
            .O(N__14572),
            .I(N__14569));
    Span4Mux_v I__1580 (
            .O(N__14569),
            .I(N__14566));
    Odrv4 I__1579 (
            .O(N__14566),
            .I(\tok.table_wr_data_10 ));
    InMux I__1578 (
            .O(N__14563),
            .I(N__14560));
    LocalMux I__1577 (
            .O(N__14560),
            .I(N__14557));
    Span4Mux_v I__1576 (
            .O(N__14557),
            .I(N__14554));
    Odrv4 I__1575 (
            .O(N__14554),
            .I(\tok.table_wr_data_15 ));
    InMux I__1574 (
            .O(N__14551),
            .I(N__14548));
    LocalMux I__1573 (
            .O(N__14548),
            .I(\tok.n33_adj_631 ));
    CascadeMux I__1572 (
            .O(N__14545),
            .I(\tok.n27_cascade_ ));
    CascadeMux I__1571 (
            .O(N__14542),
            .I(N__14538));
    CascadeMux I__1570 (
            .O(N__14541),
            .I(N__14535));
    CascadeBuf I__1569 (
            .O(N__14538),
            .I(N__14532));
    CascadeBuf I__1568 (
            .O(N__14535),
            .I(N__14529));
    CascadeMux I__1567 (
            .O(N__14532),
            .I(N__14526));
    CascadeMux I__1566 (
            .O(N__14529),
            .I(N__14523));
    InMux I__1565 (
            .O(N__14526),
            .I(N__14520));
    InMux I__1564 (
            .O(N__14523),
            .I(N__14517));
    LocalMux I__1563 (
            .O(N__14520),
            .I(N__14509));
    LocalMux I__1562 (
            .O(N__14517),
            .I(N__14509));
    InMux I__1561 (
            .O(N__14516),
            .I(N__14506));
    InMux I__1560 (
            .O(N__14515),
            .I(N__14503));
    InMux I__1559 (
            .O(N__14514),
            .I(N__14500));
    Span4Mux_v I__1558 (
            .O(N__14509),
            .I(N__14497));
    LocalMux I__1557 (
            .O(N__14506),
            .I(\tok.n41 ));
    LocalMux I__1556 (
            .O(N__14503),
            .I(\tok.n41 ));
    LocalMux I__1555 (
            .O(N__14500),
            .I(\tok.n41 ));
    Odrv4 I__1554 (
            .O(N__14497),
            .I(\tok.n41 ));
    InMux I__1553 (
            .O(N__14488),
            .I(N__14485));
    LocalMux I__1552 (
            .O(N__14485),
            .I(\tok.n33_adj_662 ));
    CascadeMux I__1551 (
            .O(N__14482),
            .I(\tok.n27_adj_709_cascade_ ));
    CascadeMux I__1550 (
            .O(N__14479),
            .I(N__14475));
    CascadeMux I__1549 (
            .O(N__14478),
            .I(N__14472));
    CascadeBuf I__1548 (
            .O(N__14475),
            .I(N__14469));
    CascadeBuf I__1547 (
            .O(N__14472),
            .I(N__14466));
    CascadeMux I__1546 (
            .O(N__14469),
            .I(N__14463));
    CascadeMux I__1545 (
            .O(N__14466),
            .I(N__14460));
    InMux I__1544 (
            .O(N__14463),
            .I(N__14457));
    InMux I__1543 (
            .O(N__14460),
            .I(N__14454));
    LocalMux I__1542 (
            .O(N__14457),
            .I(N__14446));
    LocalMux I__1541 (
            .O(N__14454),
            .I(N__14446));
    InMux I__1540 (
            .O(N__14453),
            .I(N__14443));
    InMux I__1539 (
            .O(N__14452),
            .I(N__14440));
    InMux I__1538 (
            .O(N__14451),
            .I(N__14437));
    Span4Mux_v I__1537 (
            .O(N__14446),
            .I(N__14434));
    LocalMux I__1536 (
            .O(N__14443),
            .I(\tok.n19 ));
    LocalMux I__1535 (
            .O(N__14440),
            .I(\tok.n19 ));
    LocalMux I__1534 (
            .O(N__14437),
            .I(\tok.n19 ));
    Odrv4 I__1533 (
            .O(N__14434),
            .I(\tok.n19 ));
    InMux I__1532 (
            .O(N__14425),
            .I(N__14419));
    InMux I__1531 (
            .O(N__14424),
            .I(N__14419));
    LocalMux I__1530 (
            .O(N__14419),
            .I(\tok.A_stk.tail_34 ));
    InMux I__1529 (
            .O(N__14416),
            .I(N__14410));
    InMux I__1528 (
            .O(N__14415),
            .I(N__14410));
    LocalMux I__1527 (
            .O(N__14410),
            .I(\tok.A_stk.tail_50 ));
    InMux I__1526 (
            .O(N__14407),
            .I(N__14401));
    InMux I__1525 (
            .O(N__14406),
            .I(N__14401));
    LocalMux I__1524 (
            .O(N__14401),
            .I(\tok.A_stk.tail_66 ));
    InMux I__1523 (
            .O(N__14398),
            .I(N__14392));
    InMux I__1522 (
            .O(N__14397),
            .I(N__14392));
    LocalMux I__1521 (
            .O(N__14392),
            .I(\tok.A_stk.tail_82 ));
    InMux I__1520 (
            .O(N__14389),
            .I(N__14386));
    LocalMux I__1519 (
            .O(N__14386),
            .I(N__14383));
    Span4Mux_v I__1518 (
            .O(N__14383),
            .I(N__14380));
    Odrv4 I__1517 (
            .O(N__14380),
            .I(table_wr_data_0));
    InMux I__1516 (
            .O(N__14377),
            .I(N__14373));
    InMux I__1515 (
            .O(N__14376),
            .I(N__14370));
    LocalMux I__1514 (
            .O(N__14373),
            .I(tail_98));
    LocalMux I__1513 (
            .O(N__14370),
            .I(tail_98));
    CascadeMux I__1512 (
            .O(N__14365),
            .I(N__14361));
    InMux I__1511 (
            .O(N__14364),
            .I(N__14358));
    InMux I__1510 (
            .O(N__14361),
            .I(N__14355));
    LocalMux I__1509 (
            .O(N__14358),
            .I(tail_114));
    LocalMux I__1508 (
            .O(N__14355),
            .I(tail_114));
    InMux I__1507 (
            .O(N__14350),
            .I(N__14347));
    LocalMux I__1506 (
            .O(N__14347),
            .I(N__14343));
    InMux I__1505 (
            .O(N__14346),
            .I(N__14340));
    Odrv4 I__1504 (
            .O(N__14343),
            .I(\tok.A_stk.tail_26 ));
    LocalMux I__1503 (
            .O(N__14340),
            .I(\tok.A_stk.tail_26 ));
    InMux I__1502 (
            .O(N__14335),
            .I(N__14332));
    LocalMux I__1501 (
            .O(N__14332),
            .I(N__14328));
    InMux I__1500 (
            .O(N__14331),
            .I(N__14325));
    Odrv4 I__1499 (
            .O(N__14328),
            .I(tail_126));
    LocalMux I__1498 (
            .O(N__14325),
            .I(tail_126));
    InMux I__1497 (
            .O(N__14320),
            .I(N__14317));
    LocalMux I__1496 (
            .O(N__14317),
            .I(N__14314));
    Span4Mux_s2_h I__1495 (
            .O(N__14314),
            .I(N__14310));
    InMux I__1494 (
            .O(N__14313),
            .I(N__14307));
    Odrv4 I__1493 (
            .O(N__14310),
            .I(tail_110));
    LocalMux I__1492 (
            .O(N__14307),
            .I(tail_110));
    InMux I__1491 (
            .O(N__14302),
            .I(N__14298));
    InMux I__1490 (
            .O(N__14301),
            .I(N__14295));
    LocalMux I__1489 (
            .O(N__14298),
            .I(\tok.A_stk.tail_94 ));
    LocalMux I__1488 (
            .O(N__14295),
            .I(\tok.A_stk.tail_94 ));
    InMux I__1487 (
            .O(N__14290),
            .I(N__14284));
    InMux I__1486 (
            .O(N__14289),
            .I(N__14284));
    LocalMux I__1485 (
            .O(N__14284),
            .I(\tok.A_stk.tail_78 ));
    CascadeMux I__1484 (
            .O(N__14281),
            .I(N__14278));
    InMux I__1483 (
            .O(N__14278),
            .I(N__14272));
    InMux I__1482 (
            .O(N__14277),
            .I(N__14272));
    LocalMux I__1481 (
            .O(N__14272),
            .I(\tok.A_stk.tail_62 ));
    CascadeMux I__1480 (
            .O(N__14269),
            .I(N__14266));
    InMux I__1479 (
            .O(N__14266),
            .I(N__14260));
    InMux I__1478 (
            .O(N__14265),
            .I(N__14260));
    LocalMux I__1477 (
            .O(N__14260),
            .I(\tok.A_stk.tail_46 ));
    InMux I__1476 (
            .O(N__14257),
            .I(N__14251));
    InMux I__1475 (
            .O(N__14256),
            .I(N__14251));
    LocalMux I__1474 (
            .O(N__14251),
            .I(\tok.A_stk.tail_30 ));
    InMux I__1473 (
            .O(N__14248),
            .I(N__14244));
    InMux I__1472 (
            .O(N__14247),
            .I(N__14241));
    LocalMux I__1471 (
            .O(N__14244),
            .I(\tok.A_stk.tail_14 ));
    LocalMux I__1470 (
            .O(N__14241),
            .I(\tok.A_stk.tail_14 ));
    InMux I__1469 (
            .O(N__14236),
            .I(N__14232));
    InMux I__1468 (
            .O(N__14235),
            .I(N__14229));
    LocalMux I__1467 (
            .O(N__14232),
            .I(tail_127));
    LocalMux I__1466 (
            .O(N__14229),
            .I(tail_127));
    InMux I__1465 (
            .O(N__14224),
            .I(N__14220));
    InMux I__1464 (
            .O(N__14223),
            .I(N__14217));
    LocalMux I__1463 (
            .O(N__14220),
            .I(tail_111));
    LocalMux I__1462 (
            .O(N__14217),
            .I(tail_111));
    InMux I__1461 (
            .O(N__14212),
            .I(N__14206));
    InMux I__1460 (
            .O(N__14211),
            .I(N__14206));
    LocalMux I__1459 (
            .O(N__14206),
            .I(\tok.A_stk.tail_95 ));
    InMux I__1458 (
            .O(N__14203),
            .I(N__14197));
    InMux I__1457 (
            .O(N__14202),
            .I(N__14197));
    LocalMux I__1456 (
            .O(N__14197),
            .I(\tok.A_stk.tail_79 ));
    InMux I__1455 (
            .O(N__14194),
            .I(N__14188));
    InMux I__1454 (
            .O(N__14193),
            .I(N__14188));
    LocalMux I__1453 (
            .O(N__14188),
            .I(\tok.A_stk.tail_63 ));
    InMux I__1452 (
            .O(N__14185),
            .I(N__14179));
    InMux I__1451 (
            .O(N__14184),
            .I(N__14179));
    LocalMux I__1450 (
            .O(N__14179),
            .I(\tok.A_stk.tail_47 ));
    InMux I__1449 (
            .O(N__14176),
            .I(N__14170));
    InMux I__1448 (
            .O(N__14175),
            .I(N__14170));
    LocalMux I__1447 (
            .O(N__14170),
            .I(\tok.A_stk.tail_31 ));
    CascadeMux I__1446 (
            .O(N__14167),
            .I(N__14164));
    InMux I__1445 (
            .O(N__14164),
            .I(N__14161));
    LocalMux I__1444 (
            .O(N__14161),
            .I(N__14158));
    Span12Mux_s2_h I__1443 (
            .O(N__14158),
            .I(N__14154));
    InMux I__1442 (
            .O(N__14157),
            .I(N__14151));
    Odrv12 I__1441 (
            .O(N__14154),
            .I(\tok.A_stk.tail_15 ));
    LocalMux I__1440 (
            .O(N__14151),
            .I(\tok.A_stk.tail_15 ));
    InMux I__1439 (
            .O(N__14146),
            .I(N__14142));
    InMux I__1438 (
            .O(N__14145),
            .I(N__14139));
    LocalMux I__1437 (
            .O(N__14142),
            .I(\tok.uart.txclkcounter_1 ));
    LocalMux I__1436 (
            .O(N__14139),
            .I(\tok.uart.txclkcounter_1 ));
    InMux I__1435 (
            .O(N__14134),
            .I(\tok.uart.n4830 ));
    InMux I__1434 (
            .O(N__14131),
            .I(N__14127));
    InMux I__1433 (
            .O(N__14130),
            .I(N__14124));
    LocalMux I__1432 (
            .O(N__14127),
            .I(\tok.uart.txclkcounter_2 ));
    LocalMux I__1431 (
            .O(N__14124),
            .I(\tok.uart.txclkcounter_2 ));
    InMux I__1430 (
            .O(N__14119),
            .I(\tok.uart.n4831 ));
    InMux I__1429 (
            .O(N__14116),
            .I(N__14112));
    InMux I__1428 (
            .O(N__14115),
            .I(N__14109));
    LocalMux I__1427 (
            .O(N__14112),
            .I(\tok.uart.txclkcounter_3 ));
    LocalMux I__1426 (
            .O(N__14109),
            .I(\tok.uart.txclkcounter_3 ));
    InMux I__1425 (
            .O(N__14104),
            .I(\tok.uart.n4832 ));
    InMux I__1424 (
            .O(N__14101),
            .I(N__14097));
    InMux I__1423 (
            .O(N__14100),
            .I(N__14094));
    LocalMux I__1422 (
            .O(N__14097),
            .I(\tok.uart.txclkcounter_4 ));
    LocalMux I__1421 (
            .O(N__14094),
            .I(\tok.uart.txclkcounter_4 ));
    InMux I__1420 (
            .O(N__14089),
            .I(\tok.uart.n4833 ));
    InMux I__1419 (
            .O(N__14086),
            .I(N__14082));
    InMux I__1418 (
            .O(N__14085),
            .I(N__14079));
    LocalMux I__1417 (
            .O(N__14082),
            .I(\tok.uart.txclkcounter_5 ));
    LocalMux I__1416 (
            .O(N__14079),
            .I(\tok.uart.txclkcounter_5 ));
    InMux I__1415 (
            .O(N__14074),
            .I(\tok.uart.n4834 ));
    InMux I__1414 (
            .O(N__14071),
            .I(N__14067));
    InMux I__1413 (
            .O(N__14070),
            .I(N__14064));
    LocalMux I__1412 (
            .O(N__14067),
            .I(\tok.uart.txclkcounter_6 ));
    LocalMux I__1411 (
            .O(N__14064),
            .I(\tok.uart.txclkcounter_6 ));
    InMux I__1410 (
            .O(N__14059),
            .I(\tok.uart.n4835 ));
    InMux I__1409 (
            .O(N__14056),
            .I(N__14052));
    InMux I__1408 (
            .O(N__14055),
            .I(N__14049));
    LocalMux I__1407 (
            .O(N__14052),
            .I(\tok.uart.txclkcounter_7 ));
    LocalMux I__1406 (
            .O(N__14049),
            .I(\tok.uart.txclkcounter_7 ));
    InMux I__1405 (
            .O(N__14044),
            .I(\tok.uart.n4836 ));
    InMux I__1404 (
            .O(N__14041),
            .I(bfn_1_14_0_));
    InMux I__1403 (
            .O(N__14038),
            .I(N__14034));
    InMux I__1402 (
            .O(N__14037),
            .I(N__14031));
    LocalMux I__1401 (
            .O(N__14034),
            .I(N__14028));
    LocalMux I__1400 (
            .O(N__14031),
            .I(\tok.uart.txclkcounter_8 ));
    Odrv4 I__1399 (
            .O(N__14028),
            .I(\tok.uart.txclkcounter_8 ));
    InMux I__1398 (
            .O(N__14023),
            .I(N__14020));
    LocalMux I__1397 (
            .O(N__14020),
            .I(\tok.n206_adj_691 ));
    CascadeMux I__1396 (
            .O(N__14017),
            .I(\tok.n212_adj_689_cascade_ ));
    InMux I__1395 (
            .O(N__14014),
            .I(N__14008));
    InMux I__1394 (
            .O(N__14013),
            .I(N__14008));
    LocalMux I__1393 (
            .O(N__14008),
            .I(\tok.n229_adj_863 ));
    CascadeMux I__1392 (
            .O(N__14005),
            .I(\tok.uart.n6223_cascade_ ));
    CascadeMux I__1391 (
            .O(N__14002),
            .I(txtick_cascade_));
    InMux I__1390 (
            .O(N__13999),
            .I(N__13996));
    LocalMux I__1389 (
            .O(N__13996),
            .I(\tok.uart.n12 ));
    CascadeMux I__1388 (
            .O(N__13993),
            .I(N__13989));
    InMux I__1387 (
            .O(N__13992),
            .I(N__13986));
    InMux I__1386 (
            .O(N__13989),
            .I(N__13983));
    LocalMux I__1385 (
            .O(N__13986),
            .I(\tok.uart.txclkcounter_0 ));
    LocalMux I__1384 (
            .O(N__13983),
            .I(\tok.uart.txclkcounter_0 ));
    InMux I__1383 (
            .O(N__13978),
            .I(bfn_1_13_0_));
    CascadeMux I__1382 (
            .O(N__13975),
            .I(\tok.n203_adj_833_cascade_ ));
    CascadeMux I__1381 (
            .O(N__13972),
            .I(\tok.n212_adj_835_cascade_ ));
    InMux I__1380 (
            .O(N__13969),
            .I(N__13966));
    LocalMux I__1379 (
            .O(N__13966),
            .I(\tok.n206_adj_834 ));
    CascadeMux I__1378 (
            .O(N__13963),
            .I(\tok.n6443_cascade_ ));
    CascadeMux I__1377 (
            .O(N__13960),
            .I(\tok.n242_adj_839_cascade_ ));
    InMux I__1376 (
            .O(N__13957),
            .I(N__13951));
    InMux I__1375 (
            .O(N__13956),
            .I(N__13951));
    LocalMux I__1374 (
            .O(N__13951),
            .I(\tok.n230 ));
    InMux I__1373 (
            .O(N__13948),
            .I(N__13945));
    LocalMux I__1372 (
            .O(N__13945),
            .I(\tok.n242_adj_874 ));
    CascadeMux I__1371 (
            .O(N__13942),
            .I(\tok.n6431_cascade_ ));
    InMux I__1370 (
            .O(N__13939),
            .I(N__13936));
    LocalMux I__1369 (
            .O(N__13936),
            .I(\tok.n206_adj_869 ));
    InMux I__1368 (
            .O(N__13933),
            .I(N__13930));
    LocalMux I__1367 (
            .O(N__13930),
            .I(N__13927));
    Odrv4 I__1366 (
            .O(N__13927),
            .I(\tok.table_rd_13 ));
    CascadeMux I__1365 (
            .O(N__13924),
            .I(\tok.n226_cascade_ ));
    CascadeMux I__1364 (
            .O(N__13921),
            .I(\tok.n203_adj_643_cascade_ ));
    InMux I__1363 (
            .O(N__13918),
            .I(N__13915));
    LocalMux I__1362 (
            .O(N__13915),
            .I(\tok.n226 ));
    CascadeMux I__1361 (
            .O(N__13912),
            .I(\tok.n212_adj_646_cascade_ ));
    CascadeMux I__1360 (
            .O(N__13909),
            .I(\tok.n6448_cascade_ ));
    InMux I__1359 (
            .O(N__13906),
            .I(N__13903));
    LocalMux I__1358 (
            .O(N__13903),
            .I(\tok.n6388 ));
    InMux I__1357 (
            .O(N__13900),
            .I(N__13897));
    LocalMux I__1356 (
            .O(N__13897),
            .I(\tok.n206_adj_649 ));
    InMux I__1355 (
            .O(N__13894),
            .I(N__13891));
    LocalMux I__1354 (
            .O(N__13891),
            .I(N__13888));
    Span4Mux_v I__1353 (
            .O(N__13888),
            .I(N__13885));
    Odrv4 I__1352 (
            .O(N__13885),
            .I(\tok.table_rd_9 ));
    InMux I__1351 (
            .O(N__13882),
            .I(\tok.n4773 ));
    CascadeMux I__1350 (
            .O(N__13879),
            .I(N__13875));
    InMux I__1349 (
            .O(N__13878),
            .I(N__13872));
    InMux I__1348 (
            .O(N__13875),
            .I(N__13869));
    LocalMux I__1347 (
            .O(N__13872),
            .I(tail_120));
    LocalMux I__1346 (
            .O(N__13869),
            .I(tail_120));
    InMux I__1345 (
            .O(N__13864),
            .I(N__13860));
    InMux I__1344 (
            .O(N__13863),
            .I(N__13857));
    LocalMux I__1343 (
            .O(N__13860),
            .I(tail_104));
    LocalMux I__1342 (
            .O(N__13857),
            .I(tail_104));
    InMux I__1341 (
            .O(N__13852),
            .I(N__13848));
    InMux I__1340 (
            .O(N__13851),
            .I(N__13845));
    LocalMux I__1339 (
            .O(N__13848),
            .I(\tok.A_stk.tail_88 ));
    LocalMux I__1338 (
            .O(N__13845),
            .I(\tok.A_stk.tail_88 ));
    InMux I__1337 (
            .O(N__13840),
            .I(N__13834));
    InMux I__1336 (
            .O(N__13839),
            .I(N__13834));
    LocalMux I__1335 (
            .O(N__13834),
            .I(\tok.A_stk.tail_72 ));
    InMux I__1334 (
            .O(N__13831),
            .I(N__13825));
    InMux I__1333 (
            .O(N__13830),
            .I(N__13825));
    LocalMux I__1332 (
            .O(N__13825),
            .I(\tok.A_stk.tail_56 ));
    InMux I__1331 (
            .O(N__13822),
            .I(N__13816));
    InMux I__1330 (
            .O(N__13821),
            .I(N__13816));
    LocalMux I__1329 (
            .O(N__13816),
            .I(\tok.A_stk.tail_40 ));
    InMux I__1328 (
            .O(N__13813),
            .I(N__13807));
    InMux I__1327 (
            .O(N__13812),
            .I(N__13807));
    LocalMux I__1326 (
            .O(N__13807),
            .I(\tok.A_stk.tail_24 ));
    CascadeMux I__1325 (
            .O(N__13804),
            .I(N__13801));
    InMux I__1324 (
            .O(N__13801),
            .I(N__13795));
    InMux I__1323 (
            .O(N__13800),
            .I(N__13795));
    LocalMux I__1322 (
            .O(N__13795),
            .I(\tok.A_stk.tail_8 ));
    InMux I__1321 (
            .O(N__13792),
            .I(N__13789));
    LocalMux I__1320 (
            .O(N__13789),
            .I(N__13785));
    InMux I__1319 (
            .O(N__13788),
            .I(N__13782));
    Odrv12 I__1318 (
            .O(N__13785),
            .I(\tok.A_stk.tail_0 ));
    LocalMux I__1317 (
            .O(N__13782),
            .I(\tok.A_stk.tail_0 ));
    InMux I__1316 (
            .O(N__13777),
            .I(N__13771));
    InMux I__1315 (
            .O(N__13776),
            .I(N__13771));
    LocalMux I__1314 (
            .O(N__13771),
            .I(\tok.A_stk.tail_4 ));
    InMux I__1313 (
            .O(N__13768),
            .I(bfn_1_7_0_));
    InMux I__1312 (
            .O(N__13765),
            .I(\tok.n4767 ));
    InMux I__1311 (
            .O(N__13762),
            .I(\tok.n4768 ));
    InMux I__1310 (
            .O(N__13759),
            .I(\tok.n4769 ));
    InMux I__1309 (
            .O(N__13756),
            .I(\tok.n4770 ));
    InMux I__1308 (
            .O(N__13753),
            .I(\tok.n4771 ));
    InMux I__1307 (
            .O(N__13750),
            .I(\tok.n4772 ));
    InMux I__1306 (
            .O(N__13747),
            .I(N__13744));
    LocalMux I__1305 (
            .O(N__13744),
            .I(N__13741));
    Span4Mux_h I__1304 (
            .O(N__13741),
            .I(N__13737));
    InMux I__1303 (
            .O(N__13740),
            .I(N__13734));
    Odrv4 I__1302 (
            .O(N__13737),
            .I(tail_101));
    LocalMux I__1301 (
            .O(N__13734),
            .I(tail_101));
    InMux I__1300 (
            .O(N__13729),
            .I(N__13726));
    LocalMux I__1299 (
            .O(N__13726),
            .I(N__13722));
    CascadeMux I__1298 (
            .O(N__13725),
            .I(N__13719));
    Span4Mux_s2_h I__1297 (
            .O(N__13722),
            .I(N__13716));
    InMux I__1296 (
            .O(N__13719),
            .I(N__13713));
    Odrv4 I__1295 (
            .O(N__13716),
            .I(tail_117));
    LocalMux I__1294 (
            .O(N__13713),
            .I(tail_117));
    CascadeMux I__1293 (
            .O(N__13708),
            .I(N__13705));
    InMux I__1292 (
            .O(N__13705),
            .I(N__13702));
    LocalMux I__1291 (
            .O(N__13702),
            .I(\tok.n34 ));
    InMux I__1290 (
            .O(N__13699),
            .I(N__13696));
    LocalMux I__1289 (
            .O(N__13696),
            .I(N__13692));
    InMux I__1288 (
            .O(N__13695),
            .I(N__13689));
    Span4Mux_v I__1287 (
            .O(N__13692),
            .I(N__13686));
    LocalMux I__1286 (
            .O(N__13689),
            .I(tail_100));
    Odrv4 I__1285 (
            .O(N__13686),
            .I(tail_100));
    CascadeMux I__1284 (
            .O(N__13681),
            .I(rd_15__N_300_cascade_));
    InMux I__1283 (
            .O(N__13678),
            .I(N__13674));
    InMux I__1282 (
            .O(N__13677),
            .I(N__13671));
    LocalMux I__1281 (
            .O(N__13674),
            .I(tail_116));
    LocalMux I__1280 (
            .O(N__13671),
            .I(tail_116));
    InMux I__1279 (
            .O(N__13666),
            .I(N__13662));
    InMux I__1278 (
            .O(N__13665),
            .I(N__13659));
    LocalMux I__1277 (
            .O(N__13662),
            .I(\tok.A_stk.tail_91 ));
    LocalMux I__1276 (
            .O(N__13659),
            .I(\tok.A_stk.tail_91 ));
    InMux I__1275 (
            .O(N__13654),
            .I(N__13650));
    InMux I__1274 (
            .O(N__13653),
            .I(N__13647));
    LocalMux I__1273 (
            .O(N__13650),
            .I(tail_123));
    LocalMux I__1272 (
            .O(N__13647),
            .I(tail_123));
    InMux I__1271 (
            .O(N__13642),
            .I(N__13638));
    InMux I__1270 (
            .O(N__13641),
            .I(N__13635));
    LocalMux I__1269 (
            .O(N__13638),
            .I(tail_107));
    LocalMux I__1268 (
            .O(N__13635),
            .I(tail_107));
    InMux I__1267 (
            .O(N__13630),
            .I(N__13626));
    InMux I__1266 (
            .O(N__13629),
            .I(N__13623));
    LocalMux I__1265 (
            .O(N__13626),
            .I(N__13620));
    LocalMux I__1264 (
            .O(N__13623),
            .I(N__13617));
    Span4Mux_h I__1263 (
            .O(N__13620),
            .I(N__13614));
    Odrv4 I__1262 (
            .O(N__13617),
            .I(\tok.A_stk.tail_84 ));
    Odrv4 I__1261 (
            .O(N__13614),
            .I(\tok.A_stk.tail_84 ));
    CascadeMux I__1260 (
            .O(N__13609),
            .I(N__13605));
    InMux I__1259 (
            .O(N__13608),
            .I(N__13602));
    InMux I__1258 (
            .O(N__13605),
            .I(N__13599));
    LocalMux I__1257 (
            .O(N__13602),
            .I(\tok.A_stk.tail_68 ));
    LocalMux I__1256 (
            .O(N__13599),
            .I(\tok.A_stk.tail_68 ));
    InMux I__1255 (
            .O(N__13594),
            .I(N__13588));
    InMux I__1254 (
            .O(N__13593),
            .I(N__13588));
    LocalMux I__1253 (
            .O(N__13588),
            .I(\tok.A_stk.tail_52 ));
    InMux I__1252 (
            .O(N__13585),
            .I(N__13579));
    InMux I__1251 (
            .O(N__13584),
            .I(N__13579));
    LocalMux I__1250 (
            .O(N__13579),
            .I(\tok.A_stk.tail_36 ));
    CascadeMux I__1249 (
            .O(N__13576),
            .I(N__13573));
    InMux I__1248 (
            .O(N__13573),
            .I(N__13567));
    InMux I__1247 (
            .O(N__13572),
            .I(N__13567));
    LocalMux I__1246 (
            .O(N__13567),
            .I(\tok.A_stk.tail_20 ));
    InMux I__1245 (
            .O(N__13564),
            .I(N__13560));
    InMux I__1244 (
            .O(N__13563),
            .I(N__13557));
    LocalMux I__1243 (
            .O(N__13560),
            .I(N__13554));
    LocalMux I__1242 (
            .O(N__13557),
            .I(tail_106));
    Odrv4 I__1241 (
            .O(N__13554),
            .I(tail_106));
    InMux I__1240 (
            .O(N__13549),
            .I(N__13543));
    InMux I__1239 (
            .O(N__13548),
            .I(N__13543));
    LocalMux I__1238 (
            .O(N__13543),
            .I(\tok.A_stk.tail_90 ));
    InMux I__1237 (
            .O(N__13540),
            .I(N__13536));
    InMux I__1236 (
            .O(N__13539),
            .I(N__13533));
    LocalMux I__1235 (
            .O(N__13536),
            .I(\tok.A_stk.tail_74 ));
    LocalMux I__1234 (
            .O(N__13533),
            .I(\tok.A_stk.tail_74 ));
    InMux I__1233 (
            .O(N__13528),
            .I(N__13522));
    InMux I__1232 (
            .O(N__13527),
            .I(N__13522));
    LocalMux I__1231 (
            .O(N__13522),
            .I(\tok.A_stk.tail_58 ));
    CascadeMux I__1230 (
            .O(N__13519),
            .I(N__13516));
    InMux I__1229 (
            .O(N__13516),
            .I(N__13510));
    InMux I__1228 (
            .O(N__13515),
            .I(N__13510));
    LocalMux I__1227 (
            .O(N__13510),
            .I(\tok.A_stk.tail_42 ));
    InMux I__1226 (
            .O(N__13507),
            .I(N__13503));
    InMux I__1225 (
            .O(N__13506),
            .I(N__13500));
    LocalMux I__1224 (
            .O(N__13503),
            .I(tail_109));
    LocalMux I__1223 (
            .O(N__13500),
            .I(tail_109));
    InMux I__1222 (
            .O(N__13495),
            .I(N__13491));
    InMux I__1221 (
            .O(N__13494),
            .I(N__13488));
    LocalMux I__1220 (
            .O(N__13491),
            .I(tail_125));
    LocalMux I__1219 (
            .O(N__13488),
            .I(tail_125));
    CascadeMux I__1218 (
            .O(N__13483),
            .I(N__13480));
    InMux I__1217 (
            .O(N__13480),
            .I(N__13477));
    LocalMux I__1216 (
            .O(N__13477),
            .I(N__13474));
    Odrv4 I__1215 (
            .O(N__13474),
            .I(\tok.n6274 ));
    CascadeMux I__1214 (
            .O(N__13471),
            .I(\tok.n34_cascade_ ));
    CascadeMux I__1213 (
            .O(N__13468),
            .I(A_stk_delta_1_cascade_));
    InMux I__1212 (
            .O(N__13465),
            .I(N__13461));
    InMux I__1211 (
            .O(N__13464),
            .I(N__13458));
    LocalMux I__1210 (
            .O(N__13461),
            .I(N__13455));
    LocalMux I__1209 (
            .O(N__13458),
            .I(N__13452));
    Odrv4 I__1208 (
            .O(N__13455),
            .I(tail_105));
    Odrv4 I__1207 (
            .O(N__13452),
            .I(tail_105));
    InMux I__1206 (
            .O(N__13447),
            .I(N__13444));
    LocalMux I__1205 (
            .O(N__13444),
            .I(N__13440));
    InMux I__1204 (
            .O(N__13443),
            .I(N__13437));
    Odrv4 I__1203 (
            .O(N__13440),
            .I(tail_121));
    LocalMux I__1202 (
            .O(N__13437),
            .I(tail_121));
    InMux I__1201 (
            .O(N__13432),
            .I(N__13428));
    InMux I__1200 (
            .O(N__13431),
            .I(N__13425));
    LocalMux I__1199 (
            .O(N__13428),
            .I(tail_96));
    LocalMux I__1198 (
            .O(N__13425),
            .I(tail_96));
    CascadeMux I__1197 (
            .O(N__13420),
            .I(N__13416));
    CascadeMux I__1196 (
            .O(N__13419),
            .I(N__13413));
    InMux I__1195 (
            .O(N__13416),
            .I(N__13410));
    InMux I__1194 (
            .O(N__13413),
            .I(N__13407));
    LocalMux I__1193 (
            .O(N__13410),
            .I(tail_112));
    LocalMux I__1192 (
            .O(N__13407),
            .I(tail_112));
    InMux I__1191 (
            .O(N__13402),
            .I(N__13398));
    InMux I__1190 (
            .O(N__13401),
            .I(N__13395));
    LocalMux I__1189 (
            .O(N__13398),
            .I(N__13392));
    LocalMux I__1188 (
            .O(N__13395),
            .I(N__13389));
    Odrv4 I__1187 (
            .O(N__13392),
            .I(tail_118));
    Odrv4 I__1186 (
            .O(N__13389),
            .I(tail_118));
    InMux I__1185 (
            .O(N__13384),
            .I(N__13381));
    LocalMux I__1184 (
            .O(N__13381),
            .I(N__13378));
    Span4Mux_v I__1183 (
            .O(N__13378),
            .I(N__13375));
    Span4Mux_v I__1182 (
            .O(N__13375),
            .I(N__13372));
    Odrv4 I__1181 (
            .O(N__13372),
            .I(\tok.table_wr_data_8 ));
    InMux I__1180 (
            .O(N__13369),
            .I(N__13365));
    InMux I__1179 (
            .O(N__13368),
            .I(N__13362));
    LocalMux I__1178 (
            .O(N__13365),
            .I(N__13359));
    LocalMux I__1177 (
            .O(N__13362),
            .I(\tok.A_stk.tail_89 ));
    Odrv4 I__1176 (
            .O(N__13359),
            .I(\tok.A_stk.tail_89 ));
    InMux I__1175 (
            .O(N__13354),
            .I(N__13350));
    InMux I__1174 (
            .O(N__13353),
            .I(N__13347));
    LocalMux I__1173 (
            .O(N__13350),
            .I(tail_122));
    LocalMux I__1172 (
            .O(N__13347),
            .I(tail_122));
    InMux I__1171 (
            .O(N__13342),
            .I(N__13336));
    InMux I__1170 (
            .O(N__13341),
            .I(N__13336));
    LocalMux I__1169 (
            .O(N__13336),
            .I(tail_80));
    InMux I__1168 (
            .O(N__13333),
            .I(N__13327));
    InMux I__1167 (
            .O(N__13332),
            .I(N__13327));
    LocalMux I__1166 (
            .O(N__13327),
            .I(\tok.A_stk.tail_64 ));
    InMux I__1165 (
            .O(N__13324),
            .I(N__13318));
    InMux I__1164 (
            .O(N__13323),
            .I(N__13318));
    LocalMux I__1163 (
            .O(N__13318),
            .I(tail_48));
    InMux I__1162 (
            .O(N__13315),
            .I(N__13309));
    InMux I__1161 (
            .O(N__13314),
            .I(N__13309));
    LocalMux I__1160 (
            .O(N__13309),
            .I(\tok.A_stk.tail_32 ));
    InMux I__1159 (
            .O(N__13306),
            .I(N__13300));
    InMux I__1158 (
            .O(N__13305),
            .I(N__13300));
    LocalMux I__1157 (
            .O(N__13300),
            .I(tail_16));
    InMux I__1156 (
            .O(N__13297),
            .I(N__13291));
    InMux I__1155 (
            .O(N__13296),
            .I(N__13291));
    LocalMux I__1154 (
            .O(N__13291),
            .I(\tok.A_stk.tail_9 ));
    InMux I__1153 (
            .O(N__13288),
            .I(N__13282));
    InMux I__1152 (
            .O(N__13287),
            .I(N__13282));
    LocalMux I__1151 (
            .O(N__13282),
            .I(\tok.A_stk.tail_25 ));
    InMux I__1150 (
            .O(N__13279),
            .I(N__13276));
    LocalMux I__1149 (
            .O(N__13276),
            .I(N__13273));
    Span4Mux_v I__1148 (
            .O(N__13273),
            .I(N__13269));
    InMux I__1147 (
            .O(N__13272),
            .I(N__13266));
    Odrv4 I__1146 (
            .O(N__13269),
            .I(\tok.A_stk.tail_57 ));
    LocalMux I__1145 (
            .O(N__13266),
            .I(\tok.A_stk.tail_57 ));
    InMux I__1144 (
            .O(N__13261),
            .I(N__13257));
    InMux I__1143 (
            .O(N__13260),
            .I(N__13254));
    LocalMux I__1142 (
            .O(N__13257),
            .I(N__13251));
    LocalMux I__1141 (
            .O(N__13254),
            .I(N__13248));
    Span4Mux_v I__1140 (
            .O(N__13251),
            .I(N__13245));
    Odrv4 I__1139 (
            .O(N__13248),
            .I(\tok.A_stk.tail_41 ));
    Odrv4 I__1138 (
            .O(N__13245),
            .I(\tok.A_stk.tail_41 ));
    InMux I__1137 (
            .O(N__13240),
            .I(N__13237));
    LocalMux I__1136 (
            .O(N__13237),
            .I(N__13234));
    Span4Mux_v I__1135 (
            .O(N__13234),
            .I(N__13231));
    Odrv4 I__1134 (
            .O(N__13231),
            .I(\tok.table_rd_10 ));
    CascadeMux I__1133 (
            .O(N__13228),
            .I(\tok.n203_adj_866_cascade_ ));
    CascadeMux I__1132 (
            .O(N__13225),
            .I(\tok.n212_adj_867_cascade_ ));
    CascadeMux I__1131 (
            .O(N__13222),
            .I(\tok.n6426_cascade_ ));
    InMux I__1130 (
            .O(N__13219),
            .I(N__13213));
    InMux I__1129 (
            .O(N__13218),
            .I(N__13213));
    LocalMux I__1128 (
            .O(N__13213),
            .I(\tok.A_stk.tail_85 ));
    InMux I__1127 (
            .O(N__13210),
            .I(N__13204));
    InMux I__1126 (
            .O(N__13209),
            .I(N__13204));
    LocalMux I__1125 (
            .O(N__13204),
            .I(\tok.A_stk.tail_69 ));
    InMux I__1124 (
            .O(N__13201),
            .I(N__13195));
    InMux I__1123 (
            .O(N__13200),
            .I(N__13195));
    LocalMux I__1122 (
            .O(N__13195),
            .I(\tok.A_stk.tail_53 ));
    InMux I__1121 (
            .O(N__13192),
            .I(N__13186));
    InMux I__1120 (
            .O(N__13191),
            .I(N__13186));
    LocalMux I__1119 (
            .O(N__13186),
            .I(\tok.A_stk.tail_37 ));
    InMux I__1118 (
            .O(N__13183),
            .I(N__13179));
    InMux I__1117 (
            .O(N__13182),
            .I(N__13176));
    LocalMux I__1116 (
            .O(N__13179),
            .I(\tok.A_stk.tail_21 ));
    LocalMux I__1115 (
            .O(N__13176),
            .I(\tok.A_stk.tail_21 ));
    CascadeMux I__1114 (
            .O(N__13171),
            .I(N__13168));
    InMux I__1113 (
            .O(N__13168),
            .I(N__13162));
    InMux I__1112 (
            .O(N__13167),
            .I(N__13162));
    LocalMux I__1111 (
            .O(N__13162),
            .I(\tok.A_stk.tail_5 ));
    InMux I__1110 (
            .O(N__13159),
            .I(N__13156));
    LocalMux I__1109 (
            .O(N__13156),
            .I(N__13152));
    InMux I__1108 (
            .O(N__13155),
            .I(N__13149));
    Odrv4 I__1107 (
            .O(N__13152),
            .I(\tok.A_stk.tail_11 ));
    LocalMux I__1106 (
            .O(N__13149),
            .I(\tok.A_stk.tail_11 ));
    InMux I__1105 (
            .O(N__13144),
            .I(N__13138));
    InMux I__1104 (
            .O(N__13143),
            .I(N__13138));
    LocalMux I__1103 (
            .O(N__13138),
            .I(\tok.A_stk.tail_29 ));
    CascadeMux I__1102 (
            .O(N__13135),
            .I(N__13132));
    InMux I__1101 (
            .O(N__13132),
            .I(N__13126));
    InMux I__1100 (
            .O(N__13131),
            .I(N__13126));
    LocalMux I__1099 (
            .O(N__13126),
            .I(\tok.A_stk.tail_13 ));
    InMux I__1098 (
            .O(N__13123),
            .I(N__13117));
    InMux I__1097 (
            .O(N__13122),
            .I(N__13117));
    LocalMux I__1096 (
            .O(N__13117),
            .I(\tok.A_stk.tail_75 ));
    InMux I__1095 (
            .O(N__13114),
            .I(N__13108));
    InMux I__1094 (
            .O(N__13113),
            .I(N__13108));
    LocalMux I__1093 (
            .O(N__13108),
            .I(\tok.A_stk.tail_59 ));
    InMux I__1092 (
            .O(N__13105),
            .I(N__13099));
    InMux I__1091 (
            .O(N__13104),
            .I(N__13099));
    LocalMux I__1090 (
            .O(N__13099),
            .I(\tok.A_stk.tail_43 ));
    InMux I__1089 (
            .O(N__13096),
            .I(N__13090));
    InMux I__1088 (
            .O(N__13095),
            .I(N__13090));
    LocalMux I__1087 (
            .O(N__13090),
            .I(\tok.A_stk.tail_27 ));
    InMux I__1086 (
            .O(N__13087),
            .I(N__13081));
    InMux I__1085 (
            .O(N__13086),
            .I(N__13081));
    LocalMux I__1084 (
            .O(N__13081),
            .I(\tok.A_stk.tail_73 ));
    InMux I__1083 (
            .O(N__13078),
            .I(N__13074));
    InMux I__1082 (
            .O(N__13077),
            .I(N__13071));
    LocalMux I__1081 (
            .O(N__13074),
            .I(\tok.A_stk.tail_93 ));
    LocalMux I__1080 (
            .O(N__13071),
            .I(\tok.A_stk.tail_93 ));
    InMux I__1079 (
            .O(N__13066),
            .I(N__13060));
    InMux I__1078 (
            .O(N__13065),
            .I(N__13060));
    LocalMux I__1077 (
            .O(N__13060),
            .I(\tok.A_stk.tail_77 ));
    InMux I__1076 (
            .O(N__13057),
            .I(N__13051));
    InMux I__1075 (
            .O(N__13056),
            .I(N__13051));
    LocalMux I__1074 (
            .O(N__13051),
            .I(\tok.A_stk.tail_61 ));
    InMux I__1073 (
            .O(N__13048),
            .I(N__13042));
    InMux I__1072 (
            .O(N__13047),
            .I(N__13042));
    LocalMux I__1071 (
            .O(N__13042),
            .I(\tok.A_stk.tail_45 ));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\tok.uart.n4837 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(\tok.n4788_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(\tok.n4796 ),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(\tok.n4781 ),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_6_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_2_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(\tok.n4803_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(\tok.n4810_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_4_11_0_));
    GND GND (
            .Y(GNDG0));
    defparam OSCInst0.CLKHF_DIV="0b01";
    SB_HFOSC OSCInst0 (
            .CLKHFPU(N__17536),
            .CLKHFEN(N__17535),
            .CLKHF(clk));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i57_LC_0_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i57_LC_0_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i57_LC_0_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i57_LC_0_4_1  (
            .in0(N__13261),
            .in1(N__13087),
            .in2(_gnd_net_),
            .in3(N__18201),
            .lcout(\tok.A_stk.tail_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38428),
            .ce(N__17919),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i89_LC_0_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i89_LC_0_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i89_LC_0_4_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i89_LC_0_4_3  (
            .in0(N__13464),
            .in1(N__13086),
            .in2(_gnd_net_),
            .in3(N__18203),
            .lcout(\tok.A_stk.tail_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38428),
            .ce(N__17919),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i73_LC_0_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i73_LC_0_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i73_LC_0_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i73_LC_0_4_6  (
            .in0(N__18202),
            .in1(N__13368),
            .in2(_gnd_net_),
            .in3(N__13272),
            .lcout(\tok.A_stk.tail_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38428),
            .ce(N__17919),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i109_LC_0_5_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i109_LC_0_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i109_LC_0_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i109_LC_0_5_0  (
            .in0(N__13494),
            .in1(N__13077),
            .in2(_gnd_net_),
            .in3(N__18181),
            .lcout(tail_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38431),
            .ce(N__17936),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i93_LC_0_5_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i93_LC_0_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i93_LC_0_5_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i93_LC_0_5_1  (
            .in0(N__18187),
            .in1(N__13506),
            .in2(_gnd_net_),
            .in3(N__13065),
            .lcout(\tok.A_stk.tail_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38431),
            .ce(N__17936),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i77_LC_0_5_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i77_LC_0_5_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i77_LC_0_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i77_LC_0_5_2  (
            .in0(N__13078),
            .in1(N__13056),
            .in2(_gnd_net_),
            .in3(N__18186),
            .lcout(\tok.A_stk.tail_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38431),
            .ce(N__17936),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i61_LC_0_5_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i61_LC_0_5_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i61_LC_0_5_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i61_LC_0_5_3  (
            .in0(N__18185),
            .in1(N__13047),
            .in2(_gnd_net_),
            .in3(N__13066),
            .lcout(\tok.A_stk.tail_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38431),
            .ce(N__17936),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i45_LC_0_5_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i45_LC_0_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i45_LC_0_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i45_LC_0_5_4  (
            .in0(N__13143),
            .in1(N__13057),
            .in2(_gnd_net_),
            .in3(N__18184),
            .lcout(\tok.A_stk.tail_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38431),
            .ce(N__17936),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i29_LC_0_5_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i29_LC_0_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i29_LC_0_5_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.A_stk.tail_i0_i29_LC_0_5_5  (
            .in0(N__18183),
            .in1(_gnd_net_),
            .in2(N__13135),
            .in3(N__13048),
            .lcout(\tok.A_stk.tail_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38431),
            .ce(N__17936),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i13_LC_0_5_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i13_LC_0_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i13_LC_0_5_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i13_LC_0_5_6  (
            .in0(N__13144),
            .in1(N__18182),
            .in2(_gnd_net_),
            .in3(N__17288),
            .lcout(\tok.A_stk.tail_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38431),
            .ce(N__17936),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i13_LC_0_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i13_LC_0_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i13_LC_0_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i13_LC_0_5_7  (
            .in0(N__13131),
            .in1(N__18569),
            .in2(_gnd_net_),
            .in3(N__32232),
            .lcout(\tok.S_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38431),
            .ce(N__17936),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i91_LC_0_6_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i91_LC_0_6_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i91_LC_0_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i91_LC_0_6_1  (
            .in0(N__18194),
            .in1(N__13641),
            .in2(_gnd_net_),
            .in3(N__13122),
            .lcout(\tok.A_stk.tail_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38435),
            .ce(N__17874),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i75_LC_0_6_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i75_LC_0_6_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i75_LC_0_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i75_LC_0_6_2  (
            .in0(N__13666),
            .in1(N__13113),
            .in2(_gnd_net_),
            .in3(N__18192),
            .lcout(\tok.A_stk.tail_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38435),
            .ce(N__17874),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i59_LC_0_6_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i59_LC_0_6_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i59_LC_0_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i59_LC_0_6_3  (
            .in0(N__18191),
            .in1(N__13104),
            .in2(_gnd_net_),
            .in3(N__13123),
            .lcout(\tok.A_stk.tail_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38435),
            .ce(N__17874),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i43_LC_0_6_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i43_LC_0_6_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i43_LC_0_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i43_LC_0_6_4  (
            .in0(N__13095),
            .in1(N__13114),
            .in2(_gnd_net_),
            .in3(N__18190),
            .lcout(\tok.A_stk.tail_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38435),
            .ce(N__17874),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i27_LC_0_6_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i27_LC_0_6_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i27_LC_0_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i27_LC_0_6_5  (
            .in0(N__18189),
            .in1(N__13155),
            .in2(_gnd_net_),
            .in3(N__13105),
            .lcout(\tok.A_stk.tail_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38435),
            .ce(N__17874),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i11_LC_0_6_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i11_LC_0_6_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i11_LC_0_6_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i11_LC_0_6_6  (
            .in0(N__13096),
            .in1(N__18188),
            .in2(_gnd_net_),
            .in3(N__19470),
            .lcout(\tok.A_stk.tail_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38435),
            .ce(N__17874),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i84_LC_0_6_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i84_LC_0_6_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i84_LC_0_6_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.A_stk.tail_i0_i84_LC_0_6_7  (
            .in0(N__18193),
            .in1(_gnd_net_),
            .in2(N__13609),
            .in3(N__13699),
            .lcout(\tok.A_stk.tail_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38435),
            .ce(N__17874),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i101_LC_0_7_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i101_LC_0_7_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i101_LC_0_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i101_LC_0_7_0  (
            .in0(N__13729),
            .in1(N__13218),
            .in2(_gnd_net_),
            .in3(N__18356),
            .lcout(tail_101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38440),
            .ce(N__17946),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i85_LC_0_7_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i85_LC_0_7_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i85_LC_0_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i85_LC_0_7_1  (
            .in0(N__18362),
            .in1(N__13740),
            .in2(_gnd_net_),
            .in3(N__13209),
            .lcout(\tok.A_stk.tail_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38440),
            .ce(N__17946),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i69_LC_0_7_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i69_LC_0_7_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i69_LC_0_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i69_LC_0_7_2  (
            .in0(N__13200),
            .in1(N__13219),
            .in2(_gnd_net_),
            .in3(N__18361),
            .lcout(\tok.A_stk.tail_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38440),
            .ce(N__17946),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i53_LC_0_7_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i53_LC_0_7_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i53_LC_0_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i53_LC_0_7_3  (
            .in0(N__18359),
            .in1(N__13210),
            .in2(_gnd_net_),
            .in3(N__13191),
            .lcout(\tok.A_stk.tail_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38440),
            .ce(N__17946),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i37_LC_0_7_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i37_LC_0_7_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i37_LC_0_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i37_LC_0_7_4  (
            .in0(N__13201),
            .in1(N__13182),
            .in2(_gnd_net_),
            .in3(N__18358),
            .lcout(\tok.A_stk.tail_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38440),
            .ce(N__17946),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i21_LC_0_7_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i21_LC_0_7_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i21_LC_0_7_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.A_stk.tail_i0_i21_LC_0_7_5  (
            .in0(N__18357),
            .in1(_gnd_net_),
            .in2(N__13171),
            .in3(N__13192),
            .lcout(\tok.A_stk.tail_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38440),
            .ce(N__17946),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i5_LC_0_7_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i5_LC_0_7_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i5_LC_0_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i5_LC_0_7_6  (
            .in0(N__13183),
            .in1(N__18360),
            .in2(_gnd_net_),
            .in3(N__21986),
            .lcout(\tok.A_stk.tail_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38440),
            .ce(N__17946),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i5_LC_0_7_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i5_LC_0_7_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i5_LC_0_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i5_LC_0_7_7  (
            .in0(N__13167),
            .in1(N__18586),
            .in2(_gnd_net_),
            .in3(N__30343),
            .lcout(\tok.S_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38440),
            .ce(N__17946),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i11_LC_0_8_0 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i11_LC_0_8_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i11_LC_0_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i11_LC_0_8_0  (
            .in0(N__13159),
            .in1(N__18587),
            .in2(_gnd_net_),
            .in3(N__24000),
            .lcout(\tok.S_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38445),
            .ce(N__17923),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i9_LC_0_8_2 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i9_LC_0_8_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i9_LC_0_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i9_LC_0_8_2  (
            .in0(N__13296),
            .in1(N__18588),
            .in2(_gnd_net_),
            .in3(N__26803),
            .lcout(\tok.S_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38445),
            .ce(N__17923),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i15_LC_0_8_3 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i15_LC_0_8_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i15_LC_0_8_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \tok.A_stk.head_i0_i15_LC_0_8_3  (
            .in0(_gnd_net_),
            .in1(N__24198),
            .in2(N__14167),
            .in3(N__18589),
            .lcout(\tok.S_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38445),
            .ce(N__17923),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i9_LC_0_8_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i9_LC_0_8_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i9_LC_0_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i9_LC_0_8_4  (
            .in0(N__18347),
            .in1(N__13288),
            .in2(_gnd_net_),
            .in3(N__21737),
            .lcout(\tok.A_stk.tail_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38445),
            .ce(N__17923),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i25_LC_0_8_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i25_LC_0_8_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i25_LC_0_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i25_LC_0_8_5  (
            .in0(N__13260),
            .in1(N__13297),
            .in2(_gnd_net_),
            .in3(N__18345),
            .lcout(\tok.A_stk.tail_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38445),
            .ce(N__17923),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i41_LC_0_8_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i41_LC_0_8_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i41_LC_0_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i41_LC_0_8_6  (
            .in0(N__18346),
            .in1(N__13287),
            .in2(_gnd_net_),
            .in3(N__13279),
            .lcout(\tok.A_stk.tail_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38445),
            .ce(N__17923),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i120_LC_0_9_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i120_LC_0_9_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i120_LC_0_9_3 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \tok.A_stk.tail_i0_i120_LC_0_9_3  (
            .in0(N__18348),
            .in1(N__13864),
            .in2(N__13879),
            .in3(N__17935),
            .lcout(tail_120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38449),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i312_4_lut_adj_301_LC_0_10_1 .C_ON=1'b0;
    defparam \tok.i312_4_lut_adj_301_LC_0_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i312_4_lut_adj_301_LC_0_10_1 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \tok.i312_4_lut_adj_301_LC_0_10_1  (
            .in0(N__13240),
            .in1(N__33097),
            .in2(N__31214),
            .in3(N__14013),
            .lcout(),
            .ltout(\tok.n203_adj_866_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_302_LC_0_10_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_302_LC_0_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_302_LC_0_10_2 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \tok.i1_4_lut_adj_302_LC_0_10_2  (
            .in0(N__14014),
            .in1(N__19246),
            .in2(N__13228),
            .in3(N__31940),
            .lcout(),
            .ltout(\tok.n212_adj_867_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6917_4_lut_LC_0_10_3 .C_ON=1'b0;
    defparam \tok.i6917_4_lut_LC_0_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6917_4_lut_LC_0_10_3 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i6917_4_lut_LC_0_10_3  (
            .in0(N__31941),
            .in1(N__33430),
            .in2(N__13225),
            .in3(N__13939),
            .lcout(),
            .ltout(\tok.n6426_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_309_LC_0_10_4 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_309_LC_0_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_309_LC_0_10_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \tok.i308_4_lut_adj_309_LC_0_10_4  (
            .in0(N__26182),
            .in1(N__36981),
            .in2(N__13222),
            .in3(N__30322),
            .lcout(\tok.n242_adj_874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i300_4_lut_4_lut_LC_0_10_6 .C_ON=1'b0;
    defparam \tok.i300_4_lut_4_lut_LC_0_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i300_4_lut_4_lut_LC_0_10_6 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \tok.i300_4_lut_4_lut_LC_0_10_6  (
            .in0(N__20689),
            .in1(N__35972),
            .in2(N__24197),
            .in3(N__14866),
            .lcout(\tok.n206_adj_691 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i96_LC_1_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i96_LC_1_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i96_LC_1_2_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i96_LC_1_2_0  (
            .in0(N__18372),
            .in1(_gnd_net_),
            .in2(N__13420),
            .in3(N__13341),
            .lcout(tail_96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38426),
            .ce(N__17900),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i80_LC_1_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i80_LC_1_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i80_LC_1_2_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i80_LC_1_2_1  (
            .in0(N__13431),
            .in1(N__13332),
            .in2(_gnd_net_),
            .in3(N__18371),
            .lcout(tail_80),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38426),
            .ce(N__17900),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i64_LC_1_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i64_LC_1_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i64_LC_1_2_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i64_LC_1_2_2  (
            .in0(N__18370),
            .in1(N__13342),
            .in2(_gnd_net_),
            .in3(N__13323),
            .lcout(\tok.A_stk.tail_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38426),
            .ce(N__17900),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i48_LC_1_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i48_LC_1_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i48_LC_1_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i48_LC_1_2_3  (
            .in0(N__13314),
            .in1(N__13333),
            .in2(_gnd_net_),
            .in3(N__18369),
            .lcout(tail_48),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38426),
            .ce(N__17900),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i32_LC_1_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i32_LC_1_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i32_LC_1_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i32_LC_1_2_4  (
            .in0(N__18368),
            .in1(N__13305),
            .in2(_gnd_net_),
            .in3(N__13324),
            .lcout(\tok.A_stk.tail_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38426),
            .ce(N__17900),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i16_LC_1_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i16_LC_1_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i16_LC_1_2_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i16_LC_1_2_5  (
            .in0(N__13315),
            .in1(N__13788),
            .in2(_gnd_net_),
            .in3(N__18367),
            .lcout(tail_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38426),
            .ce(N__17900),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i0_LC_1_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i0_LC_1_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i0_LC_1_2_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i0_LC_1_2_6  (
            .in0(N__18365),
            .in1(N__13306),
            .in2(_gnd_net_),
            .in3(N__18813),
            .lcout(\tok.A_stk.tail_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38426),
            .ce(N__17900),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i102_LC_1_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i102_LC_1_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i102_LC_1_2_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i102_LC_1_2_7  (
            .in0(N__13402),
            .in1(N__15016),
            .in2(_gnd_net_),
            .in3(N__18366),
            .lcout(tail_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38426),
            .ce(N__17900),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i112_LC_1_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i112_LC_1_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i112_LC_1_3_0 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i112_LC_1_3_0  (
            .in0(N__13432),
            .in1(N__17813),
            .in2(N__13419),
            .in3(N__18216),
            .lcout(tail_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38429),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i122_LC_1_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i122_LC_1_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i122_LC_1_3_1 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \tok.A_stk.tail_i0_i122_LC_1_3_1  (
            .in0(N__18218),
            .in1(N__13353),
            .in2(N__17885),
            .in3(N__13563),
            .lcout(tail_122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38429),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7005_4_lut_4_lut_LC_1_3_2 .C_ON=1'b0;
    defparam \tok.i7005_4_lut_4_lut_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i7005_4_lut_4_lut_LC_1_3_2 .LUT_INIT=16'b0101001100010011;
    LogicCell40 \tok.i7005_4_lut_4_lut_LC_1_3_2  (
            .in0(N__31939),
            .in1(N__33296),
            .in2(N__34840),
            .in3(N__31296),
            .lcout(\tok.n6274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i118_LC_1_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i118_LC_1_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i118_LC_1_3_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \tok.A_stk.tail_i0_i118_LC_1_3_3  (
            .in0(N__18217),
            .in1(N__13401),
            .in2(N__17884),
            .in3(N__15030),
            .lcout(tail_118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38429),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i126_LC_1_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i126_LC_1_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i126_LC_1_3_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \tok.A_stk.tail_i0_i126_LC_1_3_5  (
            .in0(N__18219),
            .in1(N__14320),
            .in2(N__17886),
            .in3(N__14331),
            .lcout(tail_126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38429),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2626_2_lut_LC_1_3_7 .C_ON=1'b0;
    defparam \tok.i2626_2_lut_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2626_2_lut_LC_1_3_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i2626_2_lut_LC_1_3_7  (
            .in0(_gnd_net_),
            .in1(N__28474),
            .in2(_gnd_net_),
            .in3(N__17249),
            .lcout(\tok.table_wr_data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i105_LC_1_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i105_LC_1_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i105_LC_1_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i105_LC_1_4_0  (
            .in0(N__13447),
            .in1(N__13369),
            .in2(_gnd_net_),
            .in3(N__18168),
            .lcout(tail_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__17932),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i26_LC_1_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i26_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i26_LC_1_4_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i26_LC_1_4_1  (
            .in0(N__18170),
            .in1(_gnd_net_),
            .in2(N__13519),
            .in3(N__15202),
            .lcout(\tok.A_stk.tail_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__17932),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i100_LC_1_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i100_LC_1_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i100_LC_1_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i100_LC_1_4_2  (
            .in0(N__13678),
            .in1(N__13630),
            .in2(_gnd_net_),
            .in3(N__18167),
            .lcout(tail_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__17932),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i106_LC_1_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i106_LC_1_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i106_LC_1_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i106_LC_1_4_3  (
            .in0(N__18169),
            .in1(N__13354),
            .in2(_gnd_net_),
            .in3(N__13548),
            .lcout(tail_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__17932),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i90_LC_1_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i90_LC_1_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i90_LC_1_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i90_LC_1_4_4  (
            .in0(N__13564),
            .in1(N__13539),
            .in2(_gnd_net_),
            .in3(N__18174),
            .lcout(\tok.A_stk.tail_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__17932),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i74_LC_1_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i74_LC_1_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i74_LC_1_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i74_LC_1_4_5  (
            .in0(N__18173),
            .in1(N__13549),
            .in2(_gnd_net_),
            .in3(N__13527),
            .lcout(\tok.A_stk.tail_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__17932),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i58_LC_1_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i58_LC_1_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i58_LC_1_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i58_LC_1_4_6  (
            .in0(N__13540),
            .in1(N__13515),
            .in2(_gnd_net_),
            .in3(N__18172),
            .lcout(\tok.A_stk.tail_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__17932),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i42_LC_1_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i42_LC_1_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i42_LC_1_4_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i42_LC_1_4_7  (
            .in0(N__18171),
            .in1(N__14346),
            .in2(_gnd_net_),
            .in3(N__13528),
            .lcout(\tok.A_stk.tail_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__17932),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i125_LC_1_5_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i125_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i125_LC_1_5_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \tok.A_stk.tail_i0_i125_LC_1_5_0  (
            .in0(N__18116),
            .in1(N__13507),
            .in2(N__17812),
            .in3(N__13495),
            .lcout(tail_125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38436),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i49_4_lut_LC_1_5_1 .C_ON=1'b0;
    defparam \tok.i49_4_lut_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i49_4_lut_LC_1_5_1 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \tok.i49_4_lut_LC_1_5_1  (
            .in0(N__15328),
            .in1(N__35480),
            .in2(N__13483),
            .in3(N__36227),
            .lcout(\tok.n34 ),
            .ltout(\tok.n34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2541_2_lut_4_lut_LC_1_5_2 .C_ON=1'b0;
    defparam \tok.i2541_2_lut_4_lut_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2541_2_lut_4_lut_LC_1_5_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \tok.i2541_2_lut_4_lut_LC_1_5_2  (
            .in0(N__21348),
            .in1(N__32433),
            .in2(N__13471),
            .in3(N__25254),
            .lcout(A_stk_delta_1),
            .ltout(A_stk_delta_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i123_LC_1_5_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i123_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i123_LC_1_5_3 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \tok.A_stk.tail_i0_i123_LC_1_5_3  (
            .in0(N__13653),
            .in1(N__13642),
            .in2(N__13468),
            .in3(N__17753),
            .lcout(tail_123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38436),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i121_LC_1_5_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i121_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i121_LC_1_5_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \tok.A_stk.tail_i0_i121_LC_1_5_4  (
            .in0(N__18115),
            .in1(N__13443),
            .in2(N__17811),
            .in3(N__13465),
            .lcout(tail_121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38436),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i117_LC_1_5_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i117_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i117_LC_1_5_5 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i117_LC_1_5_5  (
            .in0(N__13747),
            .in1(N__17749),
            .in2(N__13725),
            .in3(N__18114),
            .lcout(tail_117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38436),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i426_2_lut_4_lut_LC_1_5_6 .C_ON=1'b0;
    defparam \tok.i426_2_lut_4_lut_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i426_2_lut_4_lut_LC_1_5_6 .LUT_INIT=16'b0101010111010101;
    LogicCell40 \tok.i426_2_lut_4_lut_LC_1_5_6  (
            .in0(N__21349),
            .in1(N__32434),
            .in2(N__13708),
            .in3(N__25255),
            .lcout(rd_15__N_300),
            .ltout(rd_15__N_300_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i116_LC_1_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i116_LC_1_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i116_LC_1_5_7 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \tok.A_stk.tail_i0_i116_LC_1_5_7  (
            .in0(N__13695),
            .in1(N__13677),
            .in2(N__13681),
            .in3(N__18113),
            .lcout(tail_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38436),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i107_LC_1_6_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i107_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i107_LC_1_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i107_LC_1_6_0  (
            .in0(N__13665),
            .in1(N__13654),
            .in2(_gnd_net_),
            .in3(N__18175),
            .lcout(tail_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__17933),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i4_LC_1_6_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i4_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i4_LC_1_6_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i4_LC_1_6_1  (
            .in0(N__18178),
            .in1(_gnd_net_),
            .in2(N__13576),
            .in3(N__23800),
            .lcout(\tok.A_stk.tail_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__17933),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i68_LC_1_6_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i68_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i68_LC_1_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i68_LC_1_6_2  (
            .in0(N__13593),
            .in1(N__13629),
            .in2(_gnd_net_),
            .in3(N__18180),
            .lcout(\tok.A_stk.tail_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__17933),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i52_LC_1_6_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i52_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i52_LC_1_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i52_LC_1_6_3  (
            .in0(N__18179),
            .in1(N__13584),
            .in2(_gnd_net_),
            .in3(N__13608),
            .lcout(\tok.A_stk.tail_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__17933),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i36_LC_1_6_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i36_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i36_LC_1_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i36_LC_1_6_4  (
            .in0(N__13594),
            .in1(N__13572),
            .in2(_gnd_net_),
            .in3(N__18177),
            .lcout(\tok.A_stk.tail_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__17933),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i20_LC_1_6_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i20_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i20_LC_1_6_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i20_LC_1_6_5  (
            .in0(N__18176),
            .in1(N__13585),
            .in2(_gnd_net_),
            .in3(N__13777),
            .lcout(\tok.A_stk.tail_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__17933),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i0_LC_1_6_6 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i0_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i0_LC_1_6_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i0_LC_1_6_6  (
            .in0(N__13792),
            .in1(N__18581),
            .in2(_gnd_net_),
            .in3(N__30526),
            .lcout(S_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__17933),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i4_LC_1_6_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i4_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i4_LC_1_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.head_i0_i4_LC_1_6_7  (
            .in0(N__18582),
            .in1(N__13776),
            .in2(_gnd_net_),
            .in3(N__27390),
            .lcout(\tok.S_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__17933),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_2_lut_LC_1_7_0 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_2_lut_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_2_lut_LC_1_7_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_2_lut_LC_1_7_0  (
            .in0(N__14515),
            .in1(N__14514),
            .in2(N__15739),
            .in3(N__13768),
            .lcout(\tok.n33_adj_631 ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\tok.n4767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_3_lut_LC_1_7_1 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_3_lut_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_3_lut_LC_1_7_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_3_lut_LC_1_7_1  (
            .in0(N__15461),
            .in1(N__15460),
            .in2(N__15723),
            .in3(N__13765),
            .lcout(\tok.n33_adj_632 ),
            .ltout(),
            .carryin(\tok.n4767 ),
            .carryout(\tok.n4768 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_4_lut_LC_1_7_2 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_4_lut_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_4_lut_LC_1_7_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_4_lut_LC_1_7_2  (
            .in0(N__15632),
            .in1(N__15631),
            .in2(N__15740),
            .in3(N__13762),
            .lcout(\tok.n33_adj_633 ),
            .ltout(),
            .carryin(\tok.n4768 ),
            .carryout(\tok.n4769 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_5_lut_LC_1_7_3 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_5_lut_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_5_lut_LC_1_7_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_5_lut_LC_1_7_3  (
            .in0(N__15542),
            .in1(N__15532),
            .in2(N__15724),
            .in3(N__13759),
            .lcout(\tok.n33_adj_661 ),
            .ltout(),
            .carryin(\tok.n4769 ),
            .carryout(\tok.n4770 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_6_lut_LC_1_7_4 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_6_lut_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_6_lut_LC_1_7_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_6_lut_LC_1_7_4  (
            .in0(N__14683),
            .in1(N__14682),
            .in2(N__15741),
            .in3(N__13756),
            .lcout(\tok.n33_adj_634 ),
            .ltout(),
            .carryin(\tok.n4770 ),
            .carryout(\tok.n4771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_7_lut_LC_1_7_5 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_7_lut_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_7_lut_LC_1_7_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_7_lut_LC_1_7_5  (
            .in0(N__15397),
            .in1(N__15398),
            .in2(N__15725),
            .in3(N__13753),
            .lcout(\tok.n33 ),
            .ltout(),
            .carryin(\tok.n4771 ),
            .carryout(\tok.n4772 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_8_lut_LC_1_7_6 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_8_lut_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_8_lut_LC_1_7_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_8_lut_LC_1_7_6  (
            .in0(N__15845),
            .in1(N__15844),
            .in2(N__15742),
            .in3(N__13750),
            .lcout(\tok.n33_adj_663 ),
            .ltout(),
            .carryin(\tok.n4772 ),
            .carryout(\tok.n4773 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_9_lut_LC_1_7_7 .C_ON=1'b0;
    defparam \tok.idx_7__I_0_9_lut_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_9_lut_LC_1_7_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_9_lut_LC_1_7_7  (
            .in0(N__14451),
            .in1(N__14452),
            .in2(N__15726),
            .in3(N__13882),
            .lcout(\tok.n33_adj_662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i104_LC_1_8_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i104_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i104_LC_1_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i104_LC_1_8_0  (
            .in0(N__13878),
            .in1(N__13851),
            .in2(_gnd_net_),
            .in3(N__18349),
            .lcout(tail_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38450),
            .ce(N__17926),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i88_LC_1_8_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i88_LC_1_8_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i88_LC_1_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i88_LC_1_8_1  (
            .in0(N__18354),
            .in1(N__13863),
            .in2(_gnd_net_),
            .in3(N__13839),
            .lcout(\tok.A_stk.tail_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38450),
            .ce(N__17926),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i72_LC_1_8_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i72_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i72_LC_1_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i72_LC_1_8_2  (
            .in0(N__13852),
            .in1(N__13830),
            .in2(_gnd_net_),
            .in3(N__18353),
            .lcout(\tok.A_stk.tail_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38450),
            .ce(N__17926),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i56_LC_1_8_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i56_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i56_LC_1_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i56_LC_1_8_3  (
            .in0(N__18352),
            .in1(N__13840),
            .in2(_gnd_net_),
            .in3(N__13821),
            .lcout(\tok.A_stk.tail_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38450),
            .ce(N__17926),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i40_LC_1_8_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i40_LC_1_8_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i40_LC_1_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i40_LC_1_8_4  (
            .in0(N__13812),
            .in1(N__13831),
            .in2(_gnd_net_),
            .in3(N__18351),
            .lcout(\tok.A_stk.tail_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38450),
            .ce(N__17926),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i24_LC_1_8_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i24_LC_1_8_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i24_LC_1_8_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.A_stk.tail_i0_i24_LC_1_8_5  (
            .in0(N__18350),
            .in1(_gnd_net_),
            .in2(N__13804),
            .in3(N__13822),
            .lcout(\tok.A_stk.tail_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38450),
            .ce(N__17926),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i8_LC_1_8_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i8_LC_1_8_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i8_LC_1_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i8_LC_1_8_6  (
            .in0(N__13813),
            .in1(N__18355),
            .in2(_gnd_net_),
            .in3(N__17220),
            .lcout(\tok.A_stk.tail_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38450),
            .ce(N__17926),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i8_LC_1_8_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i8_LC_1_8_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i8_LC_1_8_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i8_LC_1_8_7  (
            .in0(N__13800),
            .in1(N__18583),
            .in2(_gnd_net_),
            .in3(N__22251),
            .lcout(\tok.S_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38450),
            .ce(N__17926),
            .sr(_gnd_net_));
    defparam \tok.or_100_i14_2_lut_LC_1_9_0 .C_ON=1'b0;
    defparam \tok.or_100_i14_2_lut_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.or_100_i14_2_lut_LC_1_9_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.or_100_i14_2_lut_LC_1_9_0  (
            .in0(N__26797),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20767),
            .lcout(\tok.n226 ),
            .ltout(\tok.n226_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i312_4_lut_adj_34_LC_1_9_1 .C_ON=1'b0;
    defparam \tok.i312_4_lut_adj_34_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i312_4_lut_adj_34_LC_1_9_1 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.i312_4_lut_adj_34_LC_1_9_1  (
            .in0(N__13933),
            .in1(N__33098),
            .in2(N__13924),
            .in3(N__30972),
            .lcout(),
            .ltout(\tok.n203_adj_643_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_37_LC_1_9_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_37_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_37_LC_1_9_2 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \tok.i1_4_lut_adj_37_LC_1_9_2  (
            .in0(N__31919),
            .in1(N__19247),
            .in2(N__13921),
            .in3(N__13918),
            .lcout(),
            .ltout(\tok.n212_adj_646_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6897_4_lut_LC_1_9_3 .C_ON=1'b0;
    defparam \tok.i6897_4_lut_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6897_4_lut_LC_1_9_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \tok.i6897_4_lut_LC_1_9_3  (
            .in0(N__33415),
            .in1(N__31920),
            .in2(N__13912),
            .in3(N__13900),
            .lcout(\tok.n6383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6700_3_lut_4_lut_LC_1_9_4 .C_ON=1'b0;
    defparam \tok.i6700_3_lut_4_lut_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6700_3_lut_4_lut_LC_1_9_4 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \tok.i6700_3_lut_4_lut_LC_1_9_4  (
            .in0(N__30970),
            .in1(N__34537),
            .in2(N__26802),
            .in3(N__20766),
            .lcout(\tok.n6388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6738_3_lut_4_lut_LC_1_9_5 .C_ON=1'b0;
    defparam \tok.i6738_3_lut_4_lut_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6738_3_lut_4_lut_LC_1_9_5 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \tok.i6738_3_lut_4_lut_LC_1_9_5  (
            .in0(N__20768),
            .in1(N__30344),
            .in2(N__34706),
            .in3(N__30971),
            .lcout(),
            .ltout(\tok.n6448_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i300_4_lut_adj_265_LC_1_9_6 .C_ON=1'b0;
    defparam \tok.i300_4_lut_adj_265_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i300_4_lut_adj_265_LC_1_9_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \tok.i300_4_lut_adj_265_LC_1_9_6  (
            .in0(N__36048),
            .in1(N__20679),
            .in2(N__13909),
            .in3(N__26798),
            .lcout(\tok.n206_adj_834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i300_4_lut_adj_39_LC_1_9_7 .C_ON=1'b0;
    defparam \tok.i300_4_lut_adj_39_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i300_4_lut_adj_39_LC_1_9_7 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \tok.i300_4_lut_adj_39_LC_1_9_7  (
            .in0(N__20678),
            .in1(N__16927),
            .in2(N__36228),
            .in3(N__13906),
            .lcout(\tok.n206_adj_649 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i312_4_lut_adj_259_LC_1_10_0 .C_ON=1'b0;
    defparam \tok.i312_4_lut_adj_259_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i312_4_lut_adj_259_LC_1_10_0 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \tok.i312_4_lut_adj_259_LC_1_10_0  (
            .in0(N__13894),
            .in1(N__33099),
            .in2(N__31215),
            .in3(N__13956),
            .lcout(),
            .ltout(\tok.n203_adj_833_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_326_LC_1_10_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_326_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_326_LC_1_10_1 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_326_LC_1_10_1  (
            .in0(N__13957),
            .in1(N__31931),
            .in2(N__13975),
            .in3(N__19244),
            .lcout(),
            .ltout(\tok.n212_adj_835_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6922_4_lut_LC_1_10_2 .C_ON=1'b0;
    defparam \tok.i6922_4_lut_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6922_4_lut_LC_1_10_2 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i6922_4_lut_LC_1_10_2  (
            .in0(N__31932),
            .in1(N__33372),
            .in2(N__13972),
            .in3(N__13969),
            .lcout(),
            .ltout(\tok.n6443_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_269_LC_1_10_3 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_269_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_269_LC_1_10_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \tok.i308_4_lut_adj_269_LC_1_10_3  (
            .in0(N__26181),
            .in1(N__27363),
            .in2(N__13963),
            .in3(N__36982),
            .lcout(),
            .ltout(\tok.n242_adj_839_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_270_LC_1_10_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_270_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_270_LC_1_10_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_270_LC_1_10_4  (
            .in0(N__36983),
            .in1(N__16072),
            .in2(N__13960),
            .in3(N__35446),
            .lcout(\tok.n200_adj_840 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_100_i10_2_lut_LC_1_10_5 .C_ON=1'b0;
    defparam \tok.or_100_i10_2_lut_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.or_100_i10_2_lut_LC_1_10_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.or_100_i10_2_lut_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__30321),
            .in2(_gnd_net_),
            .in3(N__20765),
            .lcout(\tok.n230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_310_LC_1_10_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_310_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_310_LC_1_10_7 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_310_LC_1_10_7  (
            .in0(N__35445),
            .in1(N__36984),
            .in2(N__19039),
            .in3(N__13948),
            .lcout(\tok.n200_adj_875 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6730_3_lut_4_lut_LC_1_11_1 .C_ON=1'b0;
    defparam \tok.i6730_3_lut_4_lut_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6730_3_lut_4_lut_LC_1_11_1 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \tok.i6730_3_lut_4_lut_LC_1_11_1  (
            .in0(N__34547),
            .in1(N__30973),
            .in2(N__20781),
            .in3(N__30084),
            .lcout(),
            .ltout(\tok.n6431_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i300_4_lut_adj_304_LC_1_11_2 .C_ON=1'b0;
    defparam \tok.i300_4_lut_adj_304_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i300_4_lut_adj_304_LC_1_11_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \tok.i300_4_lut_adj_304_LC_1_11_2  (
            .in0(N__20656),
            .in1(N__35778),
            .in2(N__13942),
            .in3(N__29627),
            .lcout(\tok.n206_adj_869 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_238_LC_1_11_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_238_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_238_LC_1_11_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i1_2_lut_adj_238_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__33798),
            .in2(_gnd_net_),
            .in3(N__36897),
            .lcout(\tok.n9_adj_677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_74_LC_1_11_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_74_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_74_LC_1_11_4 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \tok.i1_4_lut_adj_74_LC_1_11_4  (
            .in0(N__31917),
            .in1(N__14917),
            .in2(N__19251),
            .in3(N__14896),
            .lcout(),
            .ltout(\tok.n212_adj_689_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6880_4_lut_LC_1_11_5 .C_ON=1'b0;
    defparam \tok.i6880_4_lut_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6880_4_lut_LC_1_11_5 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i6880_4_lut_LC_1_11_5  (
            .in0(N__14023),
            .in1(N__33445),
            .in2(N__14017),
            .in3(N__31918),
            .lcout(\tok.n6347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_100_i11_2_lut_LC_1_11_7 .C_ON=1'b0;
    defparam \tok.or_100_i11_2_lut_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.or_100_i11_2_lut_LC_1_11_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.or_100_i11_2_lut_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__30083),
            .in2(_gnd_net_),
            .in3(N__20761),
            .lcout(\tok.n229_adj_863 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i6139_3_lut_LC_1_12_1 .C_ON=1'b0;
    defparam \tok.uart.i6139_3_lut_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i6139_3_lut_LC_1_12_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.uart.i6139_3_lut_LC_1_12_1  (
            .in0(N__14055),
            .in1(N__14070),
            .in2(_gnd_net_),
            .in3(N__14100),
            .lcout(),
            .ltout(\tok.uart.n6223_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i7019_4_lut_LC_1_12_2 .C_ON=1'b0;
    defparam \tok.uart.i7019_4_lut_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i7019_4_lut_LC_1_12_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \tok.uart.i7019_4_lut_LC_1_12_2  (
            .in0(N__14115),
            .in1(N__14130),
            .in2(N__14005),
            .in3(N__13999),
            .lcout(txtick),
            .ltout(txtick_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i7027_2_lut_LC_1_12_3 .C_ON=1'b0;
    defparam \tok.uart.i7027_2_lut_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i7027_2_lut_LC_1_12_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \tok.uart.i7027_2_lut_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14002),
            .in3(N__37556),
            .lcout(\tok.uart.n950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i2_LC_1_12_5 .C_ON=1'b0;
    defparam \tok.uart.sender_i2_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i2_LC_1_12_5 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \tok.uart.sender_i2_LC_1_12_5  (
            .in0(N__14964),
            .in1(N__37591),
            .in2(N__17398),
            .in3(N__37557),
            .lcout(sender_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38472),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i5_4_lut_LC_1_12_6 .C_ON=1'b0;
    defparam \tok.uart.i5_4_lut_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5_4_lut_LC_1_12_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.uart.i5_4_lut_LC_1_12_6  (
            .in0(N__14038),
            .in1(N__14145),
            .in2(N__13993),
            .in3(N__14085),
            .lcout(\tok.uart.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_70_LC_1_12_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_70_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_70_LC_1_12_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \tok.i1_2_lut_adj_70_LC_1_12_7  (
            .in0(N__35267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30785),
            .lcout(\tok.n4_adj_636 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.txclkcounter_141__i0_LC_1_13_0 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_141__i0_LC_1_13_0 .SEQ_MODE=4'b1001;
    defparam \tok.uart.txclkcounter_141__i0_LC_1_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_141__i0_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__13992),
            .in2(_gnd_net_),
            .in3(N__13978),
            .lcout(\tok.uart.txclkcounter_0 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\tok.uart.n4830 ),
            .clk(N__38477),
            .ce(),
            .sr(N__37607));
    defparam \tok.uart.txclkcounter_141__i1_LC_1_13_1 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_141__i1_LC_1_13_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_141__i1_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_141__i1_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__14146),
            .in2(_gnd_net_),
            .in3(N__14134),
            .lcout(\tok.uart.txclkcounter_1 ),
            .ltout(),
            .carryin(\tok.uart.n4830 ),
            .carryout(\tok.uart.n4831 ),
            .clk(N__38477),
            .ce(),
            .sr(N__37607));
    defparam \tok.uart.txclkcounter_141__i2_LC_1_13_2 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_141__i2_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_141__i2_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_141__i2_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__14131),
            .in2(_gnd_net_),
            .in3(N__14119),
            .lcout(\tok.uart.txclkcounter_2 ),
            .ltout(),
            .carryin(\tok.uart.n4831 ),
            .carryout(\tok.uart.n4832 ),
            .clk(N__38477),
            .ce(),
            .sr(N__37607));
    defparam \tok.uart.txclkcounter_141__i3_LC_1_13_3 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_141__i3_LC_1_13_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_141__i3_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_141__i3_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__14116),
            .in2(_gnd_net_),
            .in3(N__14104),
            .lcout(\tok.uart.txclkcounter_3 ),
            .ltout(),
            .carryin(\tok.uart.n4832 ),
            .carryout(\tok.uart.n4833 ),
            .clk(N__38477),
            .ce(),
            .sr(N__37607));
    defparam \tok.uart.txclkcounter_141__i4_LC_1_13_4 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_141__i4_LC_1_13_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_141__i4_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_141__i4_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__14101),
            .in2(_gnd_net_),
            .in3(N__14089),
            .lcout(\tok.uart.txclkcounter_4 ),
            .ltout(),
            .carryin(\tok.uart.n4833 ),
            .carryout(\tok.uart.n4834 ),
            .clk(N__38477),
            .ce(),
            .sr(N__37607));
    defparam \tok.uart.txclkcounter_141__i5_LC_1_13_5 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_141__i5_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_141__i5_LC_1_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_141__i5_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__14086),
            .in2(_gnd_net_),
            .in3(N__14074),
            .lcout(\tok.uart.txclkcounter_5 ),
            .ltout(),
            .carryin(\tok.uart.n4834 ),
            .carryout(\tok.uart.n4835 ),
            .clk(N__38477),
            .ce(),
            .sr(N__37607));
    defparam \tok.uart.txclkcounter_141__i6_LC_1_13_6 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_141__i6_LC_1_13_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_141__i6_LC_1_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_141__i6_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__14071),
            .in2(_gnd_net_),
            .in3(N__14059),
            .lcout(\tok.uart.txclkcounter_6 ),
            .ltout(),
            .carryin(\tok.uart.n4835 ),
            .carryout(\tok.uart.n4836 ),
            .clk(N__38477),
            .ce(),
            .sr(N__37607));
    defparam \tok.uart.txclkcounter_141__i7_LC_1_13_7 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_141__i7_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_141__i7_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_141__i7_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__14056),
            .in2(_gnd_net_),
            .in3(N__14044),
            .lcout(\tok.uart.txclkcounter_7 ),
            .ltout(),
            .carryin(\tok.uart.n4836 ),
            .carryout(\tok.uart.n4837 ),
            .clk(N__38477),
            .ce(),
            .sr(N__37607));
    defparam \tok.uart.txclkcounter_141__i8_LC_1_14_0 .C_ON=1'b0;
    defparam \tok.uart.txclkcounter_141__i8_LC_1_14_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_141__i8_LC_1_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_141__i8_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__14037),
            .in2(_gnd_net_),
            .in3(N__14041),
            .lcout(\tok.uart.txclkcounter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38482),
            .ce(),
            .sr(N__37601));
    defparam \tok.A_stk.tail_i0_i119_LC_2_1_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i119_LC_2_1_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i119_LC_2_1_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i119_LC_2_1_1  (
            .in0(N__16243),
            .in1(N__17887),
            .in2(N__16260),
            .in3(N__18363),
            .lcout(tail_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38427),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i127_LC_2_1_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i127_LC_2_1_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i127_LC_2_1_6 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \tok.A_stk.tail_i0_i127_LC_2_1_6  (
            .in0(N__18364),
            .in1(N__14224),
            .in2(N__17931),
            .in3(N__14235),
            .lcout(tail_127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38427),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i111_LC_2_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i111_LC_2_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i111_LC_2_2_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i111_LC_2_2_0  (
            .in0(N__18376),
            .in1(N__14236),
            .in2(_gnd_net_),
            .in3(N__14211),
            .lcout(tail_111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38430),
            .ce(N__17901),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i95_LC_2_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i95_LC_2_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i95_LC_2_2_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i95_LC_2_2_1  (
            .in0(N__14223),
            .in1(N__18382),
            .in2(_gnd_net_),
            .in3(N__14202),
            .lcout(\tok.A_stk.tail_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38430),
            .ce(N__17901),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i79_LC_2_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i79_LC_2_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i79_LC_2_2_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i79_LC_2_2_2  (
            .in0(N__18381),
            .in1(N__14212),
            .in2(_gnd_net_),
            .in3(N__14193),
            .lcout(\tok.A_stk.tail_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38430),
            .ce(N__17901),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i63_LC_2_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i63_LC_2_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i63_LC_2_2_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.tail_i0_i63_LC_2_2_3  (
            .in0(N__14184),
            .in1(N__18380),
            .in2(_gnd_net_),
            .in3(N__14203),
            .lcout(\tok.A_stk.tail_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38430),
            .ce(N__17901),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i47_LC_2_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i47_LC_2_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i47_LC_2_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i47_LC_2_2_4  (
            .in0(N__18379),
            .in1(N__14175),
            .in2(_gnd_net_),
            .in3(N__14194),
            .lcout(\tok.A_stk.tail_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38430),
            .ce(N__17901),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i31_LC_2_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i31_LC_2_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i31_LC_2_2_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i31_LC_2_2_5  (
            .in0(N__14185),
            .in1(N__18378),
            .in2(_gnd_net_),
            .in3(N__14157),
            .lcout(\tok.A_stk.tail_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38430),
            .ce(N__17901),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i15_LC_2_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i15_LC_2_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i15_LC_2_2_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i15_LC_2_2_6  (
            .in0(N__18377),
            .in1(N__14176),
            .in2(_gnd_net_),
            .in3(N__18962),
            .lcout(\tok.A_stk.tail_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38430),
            .ce(N__17901),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i10_LC_2_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i10_LC_2_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i10_LC_2_2_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i10_LC_2_2_7  (
            .in0(N__14350),
            .in1(N__18375),
            .in2(_gnd_net_),
            .in3(N__20178),
            .lcout(\tok.A_stk.tail_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38430),
            .ce(N__17901),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i110_LC_2_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i110_LC_2_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i110_LC_2_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i110_LC_2_3_0  (
            .in0(N__14335),
            .in1(N__14301),
            .in2(_gnd_net_),
            .in3(N__18316),
            .lcout(tail_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38433),
            .ce(N__17948),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i94_LC_2_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i94_LC_2_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i94_LC_2_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i94_LC_2_3_1  (
            .in0(N__18322),
            .in1(N__14313),
            .in2(_gnd_net_),
            .in3(N__14289),
            .lcout(\tok.A_stk.tail_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38433),
            .ce(N__17948),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i78_LC_2_3_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i78_LC_2_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i78_LC_2_3_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i78_LC_2_3_2  (
            .in0(N__14302),
            .in1(N__14277),
            .in2(_gnd_net_),
            .in3(N__18321),
            .lcout(\tok.A_stk.tail_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38433),
            .ce(N__17948),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i46_LC_2_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i46_LC_2_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i46_LC_2_3_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i46_LC_2_3_3  (
            .in0(N__18319),
            .in1(_gnd_net_),
            .in2(N__14281),
            .in3(N__14256),
            .lcout(\tok.A_stk.tail_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38433),
            .ce(N__17948),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i62_LC_2_3_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i62_LC_2_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i62_LC_2_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i62_LC_2_3_4  (
            .in0(N__14290),
            .in1(N__14265),
            .in2(_gnd_net_),
            .in3(N__18320),
            .lcout(\tok.A_stk.tail_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38433),
            .ce(N__17948),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i30_LC_2_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i30_LC_2_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i30_LC_2_3_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i30_LC_2_3_5  (
            .in0(N__18318),
            .in1(_gnd_net_),
            .in2(N__14269),
            .in3(N__14248),
            .lcout(\tok.A_stk.tail_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38433),
            .ce(N__17948),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i14_LC_2_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i14_LC_2_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i14_LC_2_3_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i14_LC_2_3_6  (
            .in0(N__14257),
            .in1(N__18317),
            .in2(_gnd_net_),
            .in3(N__19304),
            .lcout(\tok.A_stk.tail_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38433),
            .ce(N__17948),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i14_LC_2_3_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i14_LC_2_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i14_LC_2_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i14_LC_2_3_7  (
            .in0(N__14247),
            .in1(N__18584),
            .in2(_gnd_net_),
            .in3(N__32380),
            .lcout(\tok.S_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38433),
            .ce(N__17948),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i18_LC_2_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i18_LC_2_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i18_LC_2_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i18_LC_2_4_0  (
            .in0(N__14425),
            .in1(N__17974),
            .in2(_gnd_net_),
            .in3(N__18195),
            .lcout(\tok.A_stk.tail_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38437),
            .ce(N__17934),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i34_LC_2_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i34_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i34_LC_2_4_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i34_LC_2_4_1  (
            .in0(N__18196),
            .in1(N__18468),
            .in2(_gnd_net_),
            .in3(N__14416),
            .lcout(\tok.A_stk.tail_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38437),
            .ce(N__17934),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i50_LC_2_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i50_LC_2_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i50_LC_2_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i50_LC_2_4_2  (
            .in0(N__14424),
            .in1(N__14407),
            .in2(_gnd_net_),
            .in3(N__18197),
            .lcout(\tok.A_stk.tail_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38437),
            .ce(N__17934),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i66_LC_2_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i66_LC_2_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i66_LC_2_4_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i66_LC_2_4_3  (
            .in0(N__18198),
            .in1(N__14415),
            .in2(_gnd_net_),
            .in3(N__14398),
            .lcout(\tok.A_stk.tail_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38437),
            .ce(N__17934),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i82_LC_2_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i82_LC_2_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i82_LC_2_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i82_LC_2_4_4  (
            .in0(N__14376),
            .in1(N__14406),
            .in2(_gnd_net_),
            .in3(N__18199),
            .lcout(\tok.A_stk.tail_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38437),
            .ce(N__17934),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i98_LC_2_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i98_LC_2_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i98_LC_2_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i98_LC_2_4_5  (
            .in0(N__18200),
            .in1(N__14364),
            .in2(_gnd_net_),
            .in3(N__14397),
            .lcout(tail_98),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38437),
            .ce(N__17934),
            .sr(_gnd_net_));
    defparam \tok.i6975_2_lut_3_lut_LC_2_4_7 .C_ON=1'b0;
    defparam \tok.i6975_2_lut_3_lut_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6975_2_lut_3_lut_LC_2_4_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \tok.i6975_2_lut_3_lut_LC_2_4_7  (
            .in0(N__36220),
            .in1(N__33161),
            .in2(_gnd_net_),
            .in3(N__31285),
            .lcout(\tok.n6644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1412_3_lut_LC_2_5_0.C_ON=1'b0;
    defparam i1412_3_lut_LC_2_5_0.SEQ_MODE=4'b0000;
    defparam i1412_3_lut_LC_2_5_0.LUT_INIT=16'b1010111110100000;
    LogicCell40 i1412_3_lut_LC_2_5_0 (
            .in0(N__18812),
            .in1(_gnd_net_),
            .in2(N__28473),
            .in3(N__21172),
            .lcout(table_wr_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i114_LC_2_5_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i114_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i114_LC_2_5_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i114_LC_2_5_1  (
            .in0(N__14377),
            .in1(N__17757),
            .in2(N__14365),
            .in3(N__18117),
            .lcout(tail_114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38442),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_86_LC_2_5_2 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_86_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_86_LC_2_5_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_adj_86_LC_2_5_2  (
            .in0(N__32967),
            .in1(N__31828),
            .in2(N__34560),
            .in3(N__31092),
            .lcout(\tok.n4_adj_642 ),
            .ltout(\tok.n4_adj_642_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6118_3_lut_LC_2_5_3 .C_ON=1'b0;
    defparam \tok.i6118_3_lut_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6118_3_lut_LC_2_5_3 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \tok.i6118_3_lut_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(N__16568),
            .in2(N__14593),
            .in3(N__30145),
            .lcout(\tok.n2532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_adj_262_LC_2_5_4 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_adj_262_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_adj_262_LC_2_5_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i1_3_lut_4_lut_adj_262_LC_2_5_4  (
            .in0(N__32966),
            .in1(N__31827),
            .in2(N__34559),
            .in3(N__31091),
            .lcout(\tok.n4_adj_641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2619_2_lut_LC_2_5_5 .C_ON=1'b0;
    defparam \tok.i2619_2_lut_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2619_2_lut_LC_2_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i2619_2_lut_LC_2_5_5  (
            .in0(_gnd_net_),
            .in1(N__28450),
            .in2(_gnd_net_),
            .in3(N__17298),
            .lcout(\tok.table_wr_data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2622_2_lut_LC_2_5_6 .C_ON=1'b0;
    defparam \tok.i2622_2_lut_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2622_2_lut_LC_2_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i2622_2_lut_LC_2_5_6  (
            .in0(N__28451),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20177),
            .lcout(\tok.table_wr_data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2617_2_lut_LC_2_5_7 .C_ON=1'b0;
    defparam \tok.i2617_2_lut_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2617_2_lut_LC_2_5_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i2617_2_lut_LC_2_5_7  (
            .in0(N__18951),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28449),
            .lcout(\tok.table_wr_data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_LC_2_6_1 .C_ON=1'b0;
    defparam \tok.i50_4_lut_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_LC_2_6_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \tok.i50_4_lut_LC_2_6_1  (
            .in0(N__25360),
            .in1(N__14551),
            .in2(N__30535),
            .in3(N__15801),
            .lcout(),
            .ltout(\tok.n27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i0_LC_2_6_2 .C_ON=1'b0;
    defparam \tok.idx_i0_LC_2_6_2 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i0_LC_2_6_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.idx_i0_LC_2_6_2  (
            .in0(N__14516),
            .in1(N__16779),
            .in2(N__14545),
            .in3(N__16677),
            .lcout(\tok.n41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38446),
            .ce(),
            .sr(N__29254));
    defparam \tok.i50_4_lut_adj_100_LC_2_6_3 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_100_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_100_LC_2_6_3 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \tok.i50_4_lut_adj_100_LC_2_6_3  (
            .in0(N__14488),
            .in1(N__15797),
            .in2(N__25375),
            .in3(N__37467),
            .lcout(),
            .ltout(\tok.n27_adj_709_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i7_LC_2_6_4 .C_ON=1'b0;
    defparam \tok.idx_i7_LC_2_6_4 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i7_LC_2_6_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.idx_i7_LC_2_6_4  (
            .in0(N__14453),
            .in1(N__16780),
            .in2(N__14482),
            .in3(N__16678),
            .lcout(\tok.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38446),
            .ce(),
            .sr(N__29254));
    defparam \tok.i50_4_lut_adj_94_LC_2_6_6 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_94_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_94_LC_2_6_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \tok.i50_4_lut_adj_94_LC_2_6_6  (
            .in0(N__25353),
            .in1(N__14719),
            .in2(N__15802),
            .in3(N__27389),
            .lcout(),
            .ltout(\tok.n27_adj_706_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i4_LC_2_6_7 .C_ON=1'b0;
    defparam \tok.idx_i4_LC_2_6_7 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i4_LC_2_6_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.idx_i4_LC_2_6_7  (
            .in0(N__16671),
            .in1(N__14684),
            .in2(N__14713),
            .in3(N__16781),
            .lcout(\tok.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38446),
            .ce(),
            .sr(N__29254));
    defparam \tok.i10_4_lut_LC_2_7_0 .C_ON=1'b0;
    defparam \tok.i10_4_lut_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_LC_2_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i10_4_lut_LC_2_7_0  (
            .in0(N__16608),
            .in1(N__16629),
            .in2(N__16884),
            .in3(N__16854),
            .lcout(\tok.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6974_4_lut_LC_2_7_1 .C_ON=1'b0;
    defparam \tok.i6974_4_lut_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6974_4_lut_LC_2_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i6974_4_lut_LC_2_7_1  (
            .in0(N__16864),
            .in1(N__15676),
            .in2(N__14602),
            .in3(N__15916),
            .lcout(),
            .ltout(\tok.n6667_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_41_LC_2_7_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_41_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_41_LC_2_7_2 .LUT_INIT=16'b0000100000101010;
    LogicCell40 \tok.i1_4_lut_adj_41_LC_2_7_2  (
            .in0(N__25367),
            .in1(N__14767),
            .in2(N__14656),
            .in3(N__14653),
            .lcout(\tok.found_slot ),
            .ltout(\tok.found_slot_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_4_lut_adj_291_LC_2_7_3 .C_ON=1'b0;
    defparam \tok.i2_2_lut_4_lut_adj_291_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_4_lut_adj_291_LC_2_7_3 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \tok.i2_2_lut_4_lut_adj_291_LC_2_7_3  (
            .in0(N__14644),
            .in1(N__16576),
            .in2(N__14635),
            .in3(N__30134),
            .lcout(\tok.write_slot ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6632_3_lut_LC_2_7_7 .C_ON=1'b0;
    defparam \tok.i6632_3_lut_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6632_3_lut_LC_2_7_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \tok.i6632_3_lut_LC_2_7_7  (
            .in0(N__35260),
            .in1(N__14761),
            .in2(_gnd_net_),
            .in3(N__31826),
            .lcout(\tok.n6326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_LC_2_8_0 .C_ON=1'b0;
    defparam \tok.i5_4_lut_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_LC_2_8_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \tok.i5_4_lut_LC_2_8_0  (
            .in0(N__29595),
            .in1(N__14799),
            .in2(N__14790),
            .in3(N__27039),
            .lcout(),
            .ltout(\tok.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i14_4_lut_LC_2_8_1 .C_ON=1'b0;
    defparam \tok.i14_4_lut_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i14_4_lut_LC_2_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i14_4_lut_LC_2_8_1  (
            .in0(N__14725),
            .in1(N__18673),
            .in2(N__14605),
            .in3(N__18715),
            .lcout(\tok.n30_adj_647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_100_i13_2_lut_LC_2_8_2 .C_ON=1'b0;
    defparam \tok.or_100_i13_2_lut_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.or_100_i13_2_lut_LC_2_8_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.or_100_i13_2_lut_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__22241),
            .in2(_gnd_net_),
            .in3(N__20769),
            .lcout(\tok.n227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i11_4_lut_LC_2_8_4 .C_ON=1'b0;
    defparam \tok.i11_4_lut_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i11_4_lut_LC_2_8_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i11_4_lut_LC_2_8_4  (
            .in0(N__14752),
            .in1(N__14800),
            .in2(N__14791),
            .in3(N__14739),
            .lcout(),
            .ltout(\tok.n27_adj_639_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i15_4_lut_LC_2_8_5 .C_ON=1'b0;
    defparam \tok.i15_4_lut_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i15_4_lut_LC_2_8_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i15_4_lut_LC_2_8_5  (
            .in0(N__15946),
            .in1(N__14776),
            .in2(N__14770),
            .in3(N__18766),
            .lcout(\tok.found_slot_N_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6657_4_lut_LC_2_8_6 .C_ON=1'b0;
    defparam \tok.i6657_4_lut_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6657_4_lut_LC_2_8_6 .LUT_INIT=16'b0000101100111011;
    LogicCell40 \tok.i6657_4_lut_LC_2_8_6  (
            .in0(N__36049),
            .in1(N__34710),
            .in2(N__33163),
            .in3(N__22242),
            .lcout(\tok.n6322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i13_1_lut_LC_2_9_0 .C_ON=1'b0;
    defparam \tok.inv_105_i13_1_lut_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i13_1_lut_LC_2_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i13_1_lut_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27018),
            .lcout(\tok.n313 ),
            .ltout(\tok.n313_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i300_4_lut_LC_2_9_1 .C_ON=1'b0;
    defparam \tok.i300_4_lut_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i300_4_lut_LC_2_9_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \tok.i300_4_lut_LC_2_9_1  (
            .in0(N__20677),
            .in1(N__36044),
            .in2(N__14755),
            .in3(N__14854),
            .lcout(\tok.n206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_LC_2_9_2 .C_ON=1'b0;
    defparam \tok.i6_4_lut_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_LC_2_9_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i6_4_lut_LC_2_9_2  (
            .in0(N__14751),
            .in1(N__37401),
            .in2(N__14740),
            .in3(N__33625),
            .lcout(\tok.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i11_1_lut_LC_2_9_3 .C_ON=1'b0;
    defparam \tok.inv_105_i11_1_lut_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i11_1_lut_LC_2_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i11_1_lut_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29620),
            .lcout(\tok.n315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i8_1_lut_LC_2_9_4 .C_ON=1'b0;
    defparam \tok.inv_105_i8_1_lut_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i8_1_lut_LC_2_9_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \tok.inv_105_i8_1_lut_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__37402),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i312_4_lut_LC_2_9_5 .C_ON=1'b0;
    defparam \tok.i312_4_lut_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i312_4_lut_LC_2_9_5 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \tok.i312_4_lut_LC_2_9_5  (
            .in0(N__14845),
            .in1(N__32851),
            .in2(N__31111),
            .in3(N__14835),
            .lcout(),
            .ltout(\tok.n203_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_LC_2_9_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_LC_2_9_6 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \tok.i1_4_lut_LC_2_9_6  (
            .in0(N__14836),
            .in1(N__19240),
            .in2(N__14827),
            .in3(N__31921),
            .lcout(),
            .ltout(\tok.n212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6903_4_lut_LC_2_9_7 .C_ON=1'b0;
    defparam \tok.i6903_4_lut_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6903_4_lut_LC_2_9_7 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i6903_4_lut_LC_2_9_7  (
            .in0(N__31922),
            .in1(N__33414),
            .in2(N__14824),
            .in3(N__14821),
            .lcout(\tok.n6397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_224_LC_2_10_0 .C_ON=1'b1;
    defparam \tok.i1_2_lut_adj_224_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_224_LC_2_10_0 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \tok.i1_2_lut_adj_224_LC_2_10_0  (
            .in0(N__36698),
            .in1(_gnd_net_),
            .in2(N__30857),
            .in3(_gnd_net_),
            .lcout(\tok.n5_adj_713 ),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\tok.n4774 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_99_add_2_3_lut_LC_2_10_1 .C_ON=1'b1;
    defparam \tok.sub_99_add_2_3_lut_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_99_add_2_3_lut_LC_2_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_99_add_2_3_lut_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__32827),
            .in2(_gnd_net_),
            .in3(N__14815),
            .lcout(\tok.n238 ),
            .ltout(),
            .carryin(\tok.n4774 ),
            .carryout(\tok.n4775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_99_add_2_4_lut_LC_2_10_2 .C_ON=1'b1;
    defparam \tok.sub_99_add_2_4_lut_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.sub_99_add_2_4_lut_LC_2_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_99_add_2_4_lut_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__31572),
            .in2(_gnd_net_),
            .in3(N__14812),
            .lcout(\tok.n237 ),
            .ltout(),
            .carryin(\tok.n4775 ),
            .carryout(\tok.n4776 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_99_add_2_5_lut_LC_2_10_3 .C_ON=1'b1;
    defparam \tok.sub_99_add_2_5_lut_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.sub_99_add_2_5_lut_LC_2_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_99_add_2_5_lut_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__17515),
            .in2(N__34428),
            .in3(N__14809),
            .lcout(\tok.n236 ),
            .ltout(),
            .carryin(\tok.n4776 ),
            .carryout(\tok.n4777 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_99_add_2_6_lut_LC_2_10_4 .C_ON=1'b1;
    defparam \tok.sub_99_add_2_6_lut_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.sub_99_add_2_6_lut_LC_2_10_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_99_add_2_6_lut_LC_2_10_4  (
            .in0(N__30503),
            .in1(N__35612),
            .in2(_gnd_net_),
            .in3(N__14806),
            .lcout(\tok.n235 ),
            .ltout(),
            .carryin(\tok.n4777 ),
            .carryout(\tok.n4778 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_99_add_2_7_lut_LC_2_10_5 .C_ON=1'b1;
    defparam \tok.sub_99_add_2_7_lut_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_99_add_2_7_lut_LC_2_10_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_99_add_2_7_lut_LC_2_10_5  (
            .in0(N__27560),
            .in1(N__36697),
            .in2(_gnd_net_),
            .in3(N__14803),
            .lcout(\tok.n234 ),
            .ltout(),
            .carryin(\tok.n4778 ),
            .carryout(\tok.n4779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_99_add_2_8_lut_LC_2_10_6 .C_ON=1'b1;
    defparam \tok.sub_99_add_2_8_lut_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_99_add_2_8_lut_LC_2_10_6 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_99_add_2_8_lut_LC_2_10_6  (
            .in0(N__33633),
            .in1(N__17508),
            .in2(N__35057),
            .in3(N__14878),
            .lcout(\tok.n233 ),
            .ltout(),
            .carryin(\tok.n4779 ),
            .carryout(\tok.n4780 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_99_add_2_9_lut_LC_2_10_7 .C_ON=1'b1;
    defparam \tok.sub_99_add_2_9_lut_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.sub_99_add_2_9_lut_LC_2_10_7 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_99_add_2_9_lut_LC_2_10_7  (
            .in0(N__36528),
            .in1(N__17516),
            .in2(N__33797),
            .in3(N__14875),
            .lcout(\tok.n232 ),
            .ltout(),
            .carryin(\tok.n4780 ),
            .carryout(\tok.n4781 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_99_add_2_10_lut_LC_2_11_0 .C_ON=1'b0;
    defparam \tok.sub_99_add_2_10_lut_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_99_add_2_10_lut_LC_2_11_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \tok.sub_99_add_2_10_lut_LC_2_11_0  (
            .in0(N__17507),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14872),
            .lcout(\tok.n214 ),
            .ltout(\tok.n214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6679_3_lut_4_lut_LC_2_11_1 .C_ON=1'b0;
    defparam \tok.i6679_3_lut_4_lut_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6679_3_lut_4_lut_LC_2_11_1 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \tok.i6679_3_lut_4_lut_LC_2_11_1  (
            .in0(N__30716),
            .in1(N__34269),
            .in2(N__14869),
            .in3(N__23994),
            .lcout(\tok.n6358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_258_LC_2_11_2 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_258_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_258_LC_2_11_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_258_LC_2_11_2  (
            .in0(N__34268),
            .in1(N__32781),
            .in2(_gnd_net_),
            .in3(N__30715),
            .lcout(\tok.n786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_49_LC_2_11_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_49_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_49_LC_2_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_49_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__35611),
            .in2(_gnd_net_),
            .in3(N__34267),
            .lcout(\tok.n289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_117_LC_2_11_4 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_117_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_117_LC_2_11_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_adj_117_LC_2_11_4  (
            .in0(N__35610),
            .in1(N__34917),
            .in2(N__36727),
            .in3(N__33711),
            .lcout(\tok.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6710_3_lut_4_lut_LC_2_11_6 .C_ON=1'b0;
    defparam \tok.i6710_3_lut_4_lut_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6710_3_lut_4_lut_LC_2_11_6 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \tok.i6710_3_lut_4_lut_LC_2_11_6  (
            .in0(N__34270),
            .in1(N__30717),
            .in2(N__22250),
            .in3(N__20740),
            .lcout(\tok.n6402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i14_1_lut_LC_2_11_7 .C_ON=1'b0;
    defparam \tok.inv_105_i14_1_lut_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i14_1_lut_LC_2_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i14_1_lut_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32210),
            .lcout(\tok.n312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_100_i15_2_lut_LC_2_12_0 .C_ON=1'b0;
    defparam \tok.or_100_i15_2_lut_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.or_100_i15_2_lut_LC_2_12_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.or_100_i15_2_lut_LC_2_12_0  (
            .in0(N__29621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20758),
            .lcout(\tok.n225 ),
            .ltout(\tok.n225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i312_4_lut_adj_50_LC_2_12_1 .C_ON=1'b0;
    defparam \tok.i312_4_lut_adj_50_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i312_4_lut_adj_50_LC_2_12_1 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.i312_4_lut_adj_50_LC_2_12_1  (
            .in0(N__14941),
            .in1(N__32785),
            .in2(N__14929),
            .in3(N__30721),
            .lcout(),
            .ltout(\tok.n203_adj_664_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_51_LC_2_12_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_51_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_51_LC_2_12_2 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \tok.i1_4_lut_adj_51_LC_2_12_2  (
            .in0(N__31538),
            .in1(N__19218),
            .in2(N__14926),
            .in3(N__14923),
            .lcout(\tok.n212_adj_665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_100_i16_2_lut_LC_2_12_3 .C_ON=1'b0;
    defparam \tok.or_100_i16_2_lut_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.or_100_i16_2_lut_LC_2_12_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.or_100_i16_2_lut_LC_2_12_3  (
            .in0(N__20759),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23995),
            .lcout(\tok.n224 ),
            .ltout(\tok.n224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i312_4_lut_adj_73_LC_2_12_4 .C_ON=1'b0;
    defparam \tok.i312_4_lut_adj_73_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i312_4_lut_adj_73_LC_2_12_4 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \tok.i312_4_lut_adj_73_LC_2_12_4  (
            .in0(N__30720),
            .in1(N__14911),
            .in2(N__14899),
            .in3(N__32786),
            .lcout(\tok.n203_adj_688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6689_3_lut_4_lut_LC_2_12_5 .C_ON=1'b0;
    defparam \tok.i6689_3_lut_4_lut_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6689_3_lut_4_lut_LC_2_12_5 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \tok.i6689_3_lut_4_lut_LC_2_12_5  (
            .in0(N__20760),
            .in1(N__34397),
            .in2(N__30974),
            .in3(N__29622),
            .lcout(),
            .ltout(\tok.n6373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i300_4_lut_adj_52_LC_2_12_6 .C_ON=1'b0;
    defparam \tok.i300_4_lut_adj_52_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i300_4_lut_adj_52_LC_2_12_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \tok.i300_4_lut_adj_52_LC_2_12_6  (
            .in0(N__20670),
            .in1(N__32281),
            .in2(N__14890),
            .in3(N__35722),
            .lcout(),
            .ltout(\tok.n206_adj_666_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6890_4_lut_LC_2_12_7 .C_ON=1'b0;
    defparam \tok.i6890_4_lut_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6890_4_lut_LC_2_12_7 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \tok.i6890_4_lut_LC_2_12_7  (
            .in0(N__31547),
            .in1(N__33371),
            .in2(N__14887),
            .in3(N__14884),
            .lcout(\tok.n6368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_294_LC_2_13_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_294_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_294_LC_2_13_0 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \tok.i1_4_lut_adj_294_LC_2_13_0  (
            .in0(N__36946),
            .in1(N__14974),
            .in2(N__17548),
            .in3(N__34004),
            .lcout(),
            .ltout(\tok.n281_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_300_LC_2_13_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_300_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_300_LC_2_13_1 .LUT_INIT=16'b1010000010101000;
    LogicCell40 \tok.i1_4_lut_adj_300_LC_2_13_1  (
            .in0(N__35272),
            .in1(N__14980),
            .in2(N__15001),
            .in3(N__30510),
            .lcout(),
            .ltout(\tok.n236_adj_864_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_306_LC_2_13_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_306_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_306_LC_2_13_2 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \tok.i1_4_lut_adj_306_LC_2_13_2  (
            .in0(N__30729),
            .in1(N__14992),
            .in2(N__14998),
            .in3(N__31546),
            .lcout(\tok.n5_adj_871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2624_4_lut_LC_2_13_3 .C_ON=1'b0;
    defparam \tok.i2624_4_lut_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2624_4_lut_LC_2_13_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i2624_4_lut_LC_2_13_3  (
            .in0(N__36051),
            .in1(N__30509),
            .in2(N__35444),
            .in3(N__34275),
            .lcout(),
            .ltout(\tok.n2648_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i360_4_lut_LC_2_13_4 .C_ON=1'b0;
    defparam \tok.i360_4_lut_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i360_4_lut_LC_2_13_4 .LUT_INIT=16'b0000111100100010;
    LogicCell40 \tok.i360_4_lut_LC_2_13_4  (
            .in0(N__14986),
            .in1(N__34003),
            .in2(N__14995),
            .in3(N__32789),
            .lcout(\tok.n226_adj_865 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6994_3_lut_LC_2_13_5 .C_ON=1'b0;
    defparam \tok.i6994_3_lut_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6994_3_lut_LC_2_13_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.i6994_3_lut_LC_2_13_5  (
            .in0(N__35268),
            .in1(N__36945),
            .in2(_gnd_net_),
            .in3(N__30727),
            .lcout(\tok.n6334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_LC_2_13_6 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_LC_2_13_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \tok.i1_3_lut_4_lut_LC_2_13_6  (
            .in0(N__34274),
            .in1(N__31545),
            .in2(N__33135),
            .in3(N__36052),
            .lcout(\tok.n4_adj_762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6661_4_lut_LC_2_13_7 .C_ON=1'b0;
    defparam \tok.i6661_4_lut_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6661_4_lut_LC_2_13_7 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \tok.i6661_4_lut_LC_2_13_7  (
            .in0(N__36050),
            .in1(N__34273),
            .in2(_gnd_net_),
            .in3(N__30728),
            .lcout(\tok.n6316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i1_LC_2_14_0 .C_ON=1'b0;
    defparam \tok.uart.sender_i1_LC_2_14_0 .SEQ_MODE=4'b1001;
    defparam \tok.uart.sender_i1_LC_2_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tok.uart.sender_i1_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14968),
            .lcout(tx_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38485),
            .ce(N__27163),
            .sr(N__37566));
    defparam \tok.A_stk.tail_i0_i65_LC_4_1_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i65_LC_4_1_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i65_LC_4_1_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i65_LC_4_1_0  (
            .in0(N__18448),
            .in1(N__15078),
            .in2(_gnd_net_),
            .in3(N__15070),
            .lcout(\tok.A_stk.tail_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38434),
            .ce(N__17955),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i49_LC_4_1_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i49_LC_4_1_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i49_LC_4_1_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i49_LC_4_1_1  (
            .in0(N__15088),
            .in1(N__15060),
            .in2(_gnd_net_),
            .in3(N__18447),
            .lcout(tail_49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38434),
            .ce(N__17955),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i81_LC_4_1_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i81_LC_4_1_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i81_LC_4_1_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i81_LC_4_1_2  (
            .in0(N__18449),
            .in1(N__16389),
            .in2(_gnd_net_),
            .in3(N__15087),
            .lcout(tail_81),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38434),
            .ce(N__17955),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i33_LC_4_1_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i33_LC_4_1_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i33_LC_4_1_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i33_LC_4_1_3  (
            .in0(N__15079),
            .in1(N__15048),
            .in2(_gnd_net_),
            .in3(N__18446),
            .lcout(\tok.A_stk.tail_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38434),
            .ce(N__17955),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i97_LC_4_1_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i97_LC_4_1_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i97_LC_4_1_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i97_LC_4_1_4  (
            .in0(N__18450),
            .in1(N__16378),
            .in2(_gnd_net_),
            .in3(N__15069),
            .lcout(tail_97),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38434),
            .ce(N__17955),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i17_LC_4_1_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i17_LC_4_1_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i17_LC_4_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i17_LC_4_1_5  (
            .in0(N__15040),
            .in1(N__15061),
            .in2(_gnd_net_),
            .in3(N__18444),
            .lcout(tail_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38434),
            .ce(N__17955),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i1_LC_4_1_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i1_LC_4_1_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i1_LC_4_1_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_stk.tail_i0_i1_LC_4_1_6  (
            .in0(N__18445),
            .in1(_gnd_net_),
            .in2(N__15052),
            .in3(N__23496),
            .lcout(\tok.A_stk.tail_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38434),
            .ce(N__17955),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i1_LC_4_1_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i1_LC_4_1_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i1_LC_4_1_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i1_LC_4_1_7  (
            .in0(N__15039),
            .in1(N__18585),
            .in2(_gnd_net_),
            .in3(N__27562),
            .lcout(S_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38434),
            .ce(N__17955),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i108_LC_4_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i108_LC_4_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i108_LC_4_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i108_LC_4_2_0  (
            .in0(N__16350),
            .in1(N__15258),
            .in2(_gnd_net_),
            .in3(N__18383),
            .lcout(tail_108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38438),
            .ce(N__17925),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i86_LC_4_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i86_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i86_LC_4_2_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i86_LC_4_2_1  (
            .in0(N__18389),
            .in1(N__15031),
            .in2(_gnd_net_),
            .in3(N__15144),
            .lcout(\tok.A_stk.tail_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38438),
            .ce(N__17925),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i70_LC_4_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i70_LC_4_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i70_LC_4_2_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i70_LC_4_2_2  (
            .in0(N__15135),
            .in1(N__15015),
            .in2(_gnd_net_),
            .in3(N__18388),
            .lcout(\tok.A_stk.tail_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38438),
            .ce(N__17925),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i54_LC_4_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i54_LC_4_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i54_LC_4_2_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i54_LC_4_2_3  (
            .in0(N__18386),
            .in1(N__15145),
            .in2(_gnd_net_),
            .in3(N__15126),
            .lcout(\tok.A_stk.tail_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38438),
            .ce(N__17925),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i38_LC_4_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i38_LC_4_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i38_LC_4_2_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i38_LC_4_2_4  (
            .in0(N__15136),
            .in1(N__15117),
            .in2(_gnd_net_),
            .in3(N__18385),
            .lcout(\tok.A_stk.tail_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38438),
            .ce(N__17925),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i22_LC_4_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i22_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i22_LC_4_2_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i22_LC_4_2_5  (
            .in0(N__18384),
            .in1(N__15127),
            .in2(_gnd_net_),
            .in3(N__15225),
            .lcout(\tok.A_stk.tail_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38438),
            .ce(N__17925),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i6_LC_4_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i6_LC_4_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i6_LC_4_2_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i6_LC_4_2_6  (
            .in0(N__15118),
            .in1(N__18387),
            .in2(_gnd_net_),
            .in3(N__25937),
            .lcout(\tok.A_stk.tail_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38438),
            .ce(N__17925),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i92_LC_4_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i92_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i92_LC_4_2_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i92_LC_4_2_7  (
            .in0(N__18390),
            .in1(N__16365),
            .in2(_gnd_net_),
            .in3(N__15237),
            .lcout(\tok.A_stk.tail_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38438),
            .ce(N__17925),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i12_LC_4_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i12_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i12_LC_4_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i12_LC_4_3_0  (
            .in0(N__18439),
            .in1(N__15106),
            .in2(_gnd_net_),
            .in3(N__20226),
            .lcout(\tok.A_stk.tail_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38443),
            .ce(N__17927),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i28_LC_4_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i28_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i28_LC_4_3_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i28_LC_4_3_1  (
            .in0(N__15214),
            .in1(N__15097),
            .in2(_gnd_net_),
            .in3(N__18440),
            .lcout(\tok.A_stk.tail_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38443),
            .ce(N__17927),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i44_LC_4_3_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i44_LC_4_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i44_LC_4_3_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i44_LC_4_3_2  (
            .in0(N__18441),
            .in1(N__15105),
            .in2(_gnd_net_),
            .in3(N__15247),
            .lcout(\tok.A_stk.tail_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38443),
            .ce(N__17927),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i60_LC_4_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i60_LC_4_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i60_LC_4_3_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i60_LC_4_3_3  (
            .in0(N__15238),
            .in1(N__15096),
            .in2(_gnd_net_),
            .in3(N__18442),
            .lcout(\tok.A_stk.tail_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38443),
            .ce(N__17927),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i76_LC_4_3_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i76_LC_4_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i76_LC_4_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i76_LC_4_3_4  (
            .in0(N__18443),
            .in1(N__15259),
            .in2(_gnd_net_),
            .in3(N__15246),
            .lcout(\tok.A_stk.tail_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38443),
            .ce(N__17927),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i6_LC_4_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i6_LC_4_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i6_LC_4_3_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.head_i0_i6_LC_4_3_5  (
            .in0(N__18565),
            .in1(N__15226),
            .in2(_gnd_net_),
            .in3(N__30073),
            .lcout(\tok.S_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38443),
            .ce(N__17927),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i12_LC_4_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i12_LC_4_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i12_LC_4_3_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i12_LC_4_3_6  (
            .in0(N__15213),
            .in1(N__18564),
            .in2(_gnd_net_),
            .in3(N__27038),
            .lcout(\tok.S_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38443),
            .ce(N__17927),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i10_LC_4_3_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i10_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i10_LC_4_3_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.head_i0_i10_LC_4_3_7  (
            .in0(N__18563),
            .in1(N__15201),
            .in2(_gnd_net_),
            .in3(N__29628),
            .lcout(\tok.S_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38443),
            .ce(N__17927),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i99_LC_4_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i99_LC_4_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i99_LC_4_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i99_LC_4_4_0  (
            .in0(N__18397),
            .in1(N__15273),
            .in2(_gnd_net_),
            .in3(N__15180),
            .lcout(tail_99),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38447),
            .ce(N__17924),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i83_LC_4_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i83_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i83_LC_4_4_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i83_LC_4_4_1  (
            .in0(N__15285),
            .in1(N__15171),
            .in2(_gnd_net_),
            .in3(N__18396),
            .lcout(\tok.A_stk.tail_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38447),
            .ce(N__17924),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i67_LC_4_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i67_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i67_LC_4_4_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i67_LC_4_4_2  (
            .in0(N__18395),
            .in1(N__15162),
            .in2(_gnd_net_),
            .in3(N__15181),
            .lcout(\tok.A_stk.tail_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38447),
            .ce(N__17924),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i51_LC_4_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i51_LC_4_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i51_LC_4_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i51_LC_4_4_3  (
            .in0(N__15153),
            .in1(N__15172),
            .in2(_gnd_net_),
            .in3(N__18394),
            .lcout(\tok.A_stk.tail_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38447),
            .ce(N__17924),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i35_LC_4_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i35_LC_4_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i35_LC_4_4_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i35_LC_4_4_4  (
            .in0(N__18392),
            .in1(N__15351),
            .in2(_gnd_net_),
            .in3(N__15163),
            .lcout(\tok.A_stk.tail_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38447),
            .ce(N__17924),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i19_LC_4_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i19_LC_4_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i19_LC_4_4_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \tok.A_stk.tail_i0_i19_LC_4_4_5  (
            .in0(N__15154),
            .in1(_gnd_net_),
            .in2(N__15343),
            .in3(N__18391),
            .lcout(\tok.A_stk.tail_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38447),
            .ce(N__17924),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i3_LC_4_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i3_LC_4_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i3_LC_4_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i3_LC_4_4_6  (
            .in0(N__18393),
            .in1(N__15352),
            .in2(_gnd_net_),
            .in3(N__23178),
            .lcout(\tok.A_stk.tail_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38447),
            .ce(N__17924),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i3_LC_4_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i3_LC_4_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i3_LC_4_4_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i3_LC_4_4_7  (
            .in0(N__15339),
            .in1(N__18550),
            .in2(_gnd_net_),
            .in3(N__36513),
            .lcout(\tok.S_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38447),
            .ce(N__17924),
            .sr(_gnd_net_));
    defparam \tok.i6631_4_lut_LC_4_5_1 .C_ON=1'b0;
    defparam \tok.i6631_4_lut_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6631_4_lut_LC_4_5_1 .LUT_INIT=16'b0001000000100000;
    LogicCell40 \tok.i6631_4_lut_LC_4_5_1  (
            .in0(N__34661),
            .in1(N__26512),
            .in2(N__18610),
            .in3(N__31095),
            .lcout(\tok.n6252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_4_lut_adj_299_LC_4_5_2 .C_ON=1'b0;
    defparam \tok.i1_2_lut_4_lut_adj_299_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_4_lut_adj_299_LC_4_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \tok.i1_2_lut_4_lut_adj_299_LC_4_5_2  (
            .in0(N__33240),
            .in1(N__34660),
            .in2(N__36231),
            .in3(N__32111),
            .lcout(\tok.n4 ),
            .ltout(\tok.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6594_2_lut_LC_4_5_3 .C_ON=1'b0;
    defparam \tok.i6594_2_lut_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6594_2_lut_LC_4_5_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \tok.i6594_2_lut_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15331),
            .in3(N__31094),
            .lcout(\tok.n6273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2623_2_lut_LC_4_5_4 .C_ON=1'b0;
    defparam \tok.i2623_2_lut_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2623_2_lut_LC_4_5_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i2623_2_lut_LC_4_5_4  (
            .in0(N__28425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21768),
            .lcout(\tok.table_wr_data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6993_4_lut_LC_4_5_5 .C_ON=1'b0;
    defparam \tok.i6993_4_lut_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6993_4_lut_LC_4_5_5 .LUT_INIT=16'b0000000011010001;
    LogicCell40 \tok.i6993_4_lut_LC_4_5_5  (
            .in0(N__21514),
            .in1(N__37042),
            .in2(N__15307),
            .in3(N__31096),
            .lcout(),
            .ltout(\tok.n6253_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6119_4_lut_LC_4_5_6 .C_ON=1'b0;
    defparam \tok.i6119_4_lut_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6119_4_lut_LC_4_5_6 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \tok.i6119_4_lut_LC_4_5_6  (
            .in0(N__15298),
            .in1(N__16552),
            .in2(N__15289),
            .in3(N__35199),
            .lcout(\tok.n6203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i115_LC_4_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i115_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i115_LC_4_5_7 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \tok.A_stk.tail_i0_i115_LC_4_5_7  (
            .in0(N__15286),
            .in1(N__17904),
            .in2(N__15274),
            .in3(N__18253),
            .lcout(tail_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38451),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_90_LC_4_6_0 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_90_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_90_LC_4_6_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \tok.i50_4_lut_adj_90_LC_4_6_0  (
            .in0(N__25338),
            .in1(N__15661),
            .in2(N__33646),
            .in3(N__15787),
            .lcout(),
            .ltout(\tok.n27_adj_704_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i2_LC_4_6_1 .C_ON=1'b0;
    defparam \tok.idx_i2_LC_4_6_1 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i2_LC_4_6_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.idx_i2_LC_4_6_1  (
            .in0(N__15602),
            .in1(N__16770),
            .in2(N__15649),
            .in3(N__16668),
            .lcout(\tok.n38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38457),
            .ce(),
            .sr(N__29216));
    defparam \tok.i314_4_lut_adj_266_LC_4_6_2 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_266_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_266_LC_4_6_2 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \tok.i314_4_lut_adj_266_LC_4_6_2  (
            .in0(N__27553),
            .in1(N__34461),
            .in2(N__15985),
            .in3(N__31907),
            .lcout(\tok.n161_adj_836 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_88_LC_4_6_3 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_88_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_88_LC_4_6_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \tok.i50_4_lut_adj_88_LC_4_6_3  (
            .in0(N__25343),
            .in1(N__15580),
            .in2(N__15796),
            .in3(N__27554),
            .lcout(\tok.n27_adj_703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_92_LC_4_6_4 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_92_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_92_LC_4_6_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \tok.i50_4_lut_adj_92_LC_4_6_4  (
            .in0(N__25339),
            .in1(N__36479),
            .in2(N__15568),
            .in3(N__15788),
            .lcout(),
            .ltout(\tok.n27_adj_705_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i3_LC_4_6_5 .C_ON=1'b0;
    defparam \tok.idx_i3_LC_4_6_5 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i3_LC_4_6_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.idx_i3_LC_4_6_5  (
            .in0(N__15513),
            .in1(N__16771),
            .in2(N__15553),
            .in3(N__16669),
            .lcout(\tok.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38457),
            .ce(),
            .sr(N__29216));
    defparam \tok.idx_i1_LC_4_6_6 .C_ON=1'b0;
    defparam \tok.idx_i1_LC_4_6_6 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i1_LC_4_6_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.idx_i1_LC_4_6_6  (
            .in0(N__16666),
            .in1(N__15441),
            .in2(N__16782),
            .in3(N__15484),
            .lcout(\tok.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38457),
            .ce(),
            .sr(N__29216));
    defparam \tok.idx_i5_LC_4_6_7 .C_ON=1'b0;
    defparam \tok.idx_i5_LC_4_6_7 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i5_LC_4_6_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.idx_i5_LC_4_6_7  (
            .in0(N__15378),
            .in1(N__16667),
            .in2(N__16786),
            .in3(N__15880),
            .lcout(\tok.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38457),
            .ce(),
            .sr(N__29216));
    defparam \tok.i314_4_lut_adj_40_LC_4_7_0 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_40_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_40_LC_4_7_0 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \tok.i314_4_lut_adj_40_LC_4_7_0  (
            .in0(N__30328),
            .in1(N__34481),
            .in2(N__16036),
            .in3(N__31908),
            .lcout(\tok.n161_adj_650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i6_1_lut_LC_4_7_1 .C_ON=1'b0;
    defparam \tok.inv_105_i6_1_lut_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i6_1_lut_LC_4_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i6_1_lut_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30327),
            .lcout(\tok.n320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_96_LC_4_7_2 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_96_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_96_LC_4_7_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \tok.i50_4_lut_adj_96_LC_4_7_2  (
            .in0(N__30329),
            .in1(N__25329),
            .in2(N__15783),
            .in3(N__15889),
            .lcout(\tok.n27_adj_707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_98_LC_4_7_3 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_98_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_98_LC_4_7_3 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \tok.i50_4_lut_adj_98_LC_4_7_3  (
            .in0(N__30054),
            .in1(N__15771),
            .in2(N__25359),
            .in3(N__15874),
            .lcout(),
            .ltout(\tok.n27_adj_708_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i6_LC_4_7_4 .C_ON=1'b0;
    defparam \tok.idx_i6_LC_4_7_4 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i6_LC_4_7_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.idx_i6_LC_4_7_4  (
            .in0(N__15840),
            .in1(N__16775),
            .in2(N__15865),
            .in3(N__16670),
            .lcout(\tok.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38462),
            .ce(),
            .sr(N__29259));
    defparam \tok.search_clk_I_0_1_lut_LC_4_7_5 .C_ON=1'b0;
    defparam \tok.search_clk_I_0_1_lut_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.search_clk_I_0_1_lut_LC_4_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.search_clk_I_0_1_lut_LC_4_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15767),
            .lcout(\tok.search_clk_N_137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.search_clk_359_LC_4_7_6 .C_ON=1'b0;
    defparam \tok.search_clk_359_LC_4_7_6 .SEQ_MODE=4'b1010;
    defparam \tok.search_clk_359_LC_4_7_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \tok.search_clk_359_LC_4_7_6  (
            .in0(N__15772),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.search_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38462),
            .ce(),
            .sr(N__29259));
    defparam \tok.i1_2_lut_LC_4_7_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_LC_4_7_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.i1_2_lut_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(N__15766),
            .in2(_gnd_net_),
            .in3(N__15713),
            .lcout(\tok.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_375_i13_2_lut_LC_4_8_0 .C_ON=1'b0;
    defparam \tok.T_7__I_0_375_i13_2_lut_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_375_i13_2_lut_LC_4_8_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \tok.T_7__I_0_375_i13_2_lut_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(N__33802),
            .in2(_gnd_net_),
            .in3(N__35237),
            .lcout(\tok.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7002_4_lut_LC_4_8_1 .C_ON=1'b0;
    defparam \tok.i7002_4_lut_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i7002_4_lut_LC_4_8_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i7002_4_lut_LC_4_8_1  (
            .in0(N__15955),
            .in1(N__30010),
            .in2(N__15967),
            .in3(N__30478),
            .lcout(\tok.n6670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_LC_4_8_2 .C_ON=1'b0;
    defparam \tok.i9_4_lut_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_LC_4_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_LC_4_8_2  (
            .in0(N__15924),
            .in1(N__15963),
            .in2(N__15937),
            .in3(N__15954),
            .lcout(\tok.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_31_LC_4_8_3 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_31_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_31_LC_4_8_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i2_4_lut_adj_31_LC_4_8_3  (
            .in0(N__27524),
            .in1(N__15933),
            .in2(N__27387),
            .in3(N__15925),
            .lcout(\tok.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_281_LC_4_8_4 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_281_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_281_LC_4_8_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i2_4_lut_adj_281_LC_4_8_4  (
            .in0(N__23548),
            .in1(N__27353),
            .in2(N__23843),
            .in3(N__27523),
            .lcout(\tok.n18_adj_850 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i317_4_lut_LC_4_8_5 .C_ON=1'b0;
    defparam \tok.i317_4_lut_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i317_4_lut_LC_4_8_5 .LUT_INIT=16'b0001000111000000;
    LogicCell40 \tok.i317_4_lut_LC_4_8_5  (
            .in0(N__27357),
            .in1(N__36841),
            .in2(N__23844),
            .in3(N__31041),
            .lcout(\tok.n177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6817_4_lut_LC_4_8_6 .C_ON=1'b0;
    defparam \tok.i6817_4_lut_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6817_4_lut_LC_4_8_6 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \tok.i6817_4_lut_LC_4_8_6  (
            .in0(N__16006),
            .in1(N__23616),
            .in2(N__32075),
            .in3(N__16813),
            .lcout(),
            .ltout(\tok.n6575_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i303_4_lut_adj_169_LC_4_8_7 .C_ON=1'b0;
    defparam \tok.i303_4_lut_adj_169_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i303_4_lut_adj_169_LC_4_8_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \tok.i303_4_lut_adj_169_LC_4_8_7  (
            .in0(N__35238),
            .in1(N__25892),
            .in2(N__15904),
            .in3(N__15901),
            .lcout(\tok.n252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_2_lut_LC_4_9_0 .C_ON=1'b1;
    defparam \tok.add_103_2_lut_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_2_lut_LC_4_9_0 .LUT_INIT=16'b1111111110010110;
    LogicCell40 \tok.add_103_2_lut_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(N__18828),
            .in2(N__30508),
            .in3(N__31671),
            .lcout(\tok.n2579 ),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\tok.n4797 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_3_lut_LC_4_9_1 .C_ON=1'b1;
    defparam \tok.add_103_3_lut_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_3_lut_LC_4_9_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.add_103_3_lut_LC_4_9_1  (
            .in0(N__31672),
            .in1(N__27552),
            .in2(N__23546),
            .in3(N__15895),
            .lcout(\tok.n2635 ),
            .ltout(),
            .carryin(\tok.n4797 ),
            .carryout(\tok.n4798 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_4_lut_LC_4_9_2 .C_ON=1'b1;
    defparam \tok.add_103_4_lut_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_4_lut_LC_4_9_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_4_lut_LC_4_9_2  (
            .in0(N__34460),
            .in1(N__33597),
            .in2(N__20095),
            .in3(N__15892),
            .lcout(\tok.n6615 ),
            .ltout(),
            .carryin(\tok.n4798 ),
            .carryout(\tok.n4799 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_5_lut_LC_4_9_3 .C_ON=1'b1;
    defparam \tok.add_103_5_lut_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_5_lut_LC_4_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.add_103_5_lut_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__23210),
            .in2(N__36541),
            .in3(N__16009),
            .lcout(\tok.n288 ),
            .ltout(),
            .carryin(\tok.n4799 ),
            .carryout(\tok.n4800 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_6_lut_LC_4_9_4 .C_ON=1'b1;
    defparam \tok.add_103_6_lut_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_6_lut_LC_4_9_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_6_lut_LC_4_9_4  (
            .in0(N__32853),
            .in1(N__27386),
            .in2(N__23839),
            .in3(N__16000),
            .lcout(\tok.n6556 ),
            .ltout(),
            .carryin(\tok.n4800 ),
            .carryout(\tok.n4801 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_7_lut_LC_4_9_5 .C_ON=1'b1;
    defparam \tok.add_103_7_lut_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_7_lut_LC_4_9_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_7_lut_LC_4_9_5  (
            .in0(N__32877),
            .in1(N__30319),
            .in2(N__22027),
            .in3(N__15997),
            .lcout(\tok.n6514 ),
            .ltout(),
            .carryin(\tok.n4801 ),
            .carryout(\tok.n4802 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_8_lut_LC_4_9_6 .C_ON=1'b1;
    defparam \tok.add_103_8_lut_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_8_lut_LC_4_9_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_8_lut_LC_4_9_6  (
            .in0(N__32852),
            .in1(N__30042),
            .in2(N__25971),
            .in3(N__15994),
            .lcout(\tok.n6490 ),
            .ltout(),
            .carryin(\tok.n4802 ),
            .carryout(\tok.n4803 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_8_THRU_CRY_0_LC_4_9_7 .C_ON=1'b1;
    defparam \tok.add_103_8_THRU_CRY_0_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_8_THRU_CRY_0_LC_4_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \tok.add_103_8_THRU_CRY_0_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(N__17517),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\tok.n4803 ),
            .carryout(\tok.n4803_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_9_lut_LC_4_10_0 .C_ON=1'b1;
    defparam \tok.add_103_9_lut_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_9_lut_LC_4_10_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_9_lut_LC_4_10_0  (
            .in0(N__33093),
            .in1(N__37443),
            .in2(N__28330),
            .in3(N__15991),
            .lcout(\tok.n6466 ),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\tok.n4804 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_10_lut_LC_4_10_1 .C_ON=1'b1;
    defparam \tok.add_103_10_lut_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_10_lut_LC_4_10_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_10_lut_LC_4_10_1  (
            .in0(N__16116),
            .in1(N__22233),
            .in2(N__17261),
            .in3(N__15988),
            .lcout(\tok.n6452 ),
            .ltout(),
            .carryin(\tok.n4804 ),
            .carryout(\tok.n4805 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_11_lut_LC_4_10_2 .C_ON=1'b1;
    defparam \tok.add_103_11_lut_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_11_lut_LC_4_10_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_11_lut_LC_4_10_2  (
            .in0(N__16113),
            .in1(N__26775),
            .in2(N__21772),
            .in3(N__15973),
            .lcout(\tok.n6437 ),
            .ltout(),
            .carryin(\tok.n4805 ),
            .carryout(\tok.n4806 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_12_lut_LC_4_10_3 .C_ON=1'b1;
    defparam \tok.add_103_12_lut_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_12_lut_LC_4_10_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_12_lut_LC_4_10_3  (
            .in0(N__16117),
            .in1(N__29577),
            .in2(N__20173),
            .in3(N__15970),
            .lcout(\tok.n6421 ),
            .ltout(),
            .carryin(\tok.n4806 ),
            .carryout(\tok.n4807 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_13_lut_LC_4_10_4 .C_ON=1'b1;
    defparam \tok.add_103_13_lut_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_13_lut_LC_4_10_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_13_lut_LC_4_10_4  (
            .in0(N__16115),
            .in1(N__23992),
            .in2(N__19503),
            .in3(N__16042),
            .lcout(\tok.n6406 ),
            .ltout(),
            .carryin(\tok.n4807 ),
            .carryout(\tok.n4808 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_14_lut_LC_4_10_5 .C_ON=1'b1;
    defparam \tok.add_103_14_lut_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_14_lut_LC_4_10_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_14_lut_LC_4_10_5  (
            .in0(N__16118),
            .in1(N__27036),
            .in2(N__20258),
            .in3(N__16039),
            .lcout(\tok.n6392 ),
            .ltout(),
            .carryin(\tok.n4808 ),
            .carryout(\tok.n4809 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_15_lut_LC_4_10_6 .C_ON=1'b1;
    defparam \tok.add_103_15_lut_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_15_lut_LC_4_10_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_15_lut_LC_4_10_6  (
            .in0(N__16114),
            .in1(N__32200),
            .in2(N__17320),
            .in3(N__16024),
            .lcout(\tok.n6377 ),
            .ltout(),
            .carryin(\tok.n4809 ),
            .carryout(\tok.n4810 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_15_THRU_CRY_0_LC_4_10_7 .C_ON=1'b1;
    defparam \tok.add_103_15_THRU_CRY_0_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_15_THRU_CRY_0_LC_4_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \tok.add_103_15_THRU_CRY_0_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(N__17485),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\tok.n4810 ),
            .carryout(\tok.n4810_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_16_lut_LC_4_11_0 .C_ON=1'b1;
    defparam \tok.add_103_16_lut_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_16_lut_LC_4_11_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_103_16_lut_LC_4_11_0  (
            .in0(N__16119),
            .in1(N__32368),
            .in2(N__19336),
            .in3(N__16021),
            .lcout(\tok.n6362 ),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\tok.n4811 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_103_17_lut_LC_4_11_1 .C_ON=1'b0;
    defparam \tok.add_103_17_lut_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_103_17_lut_LC_4_11_1 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \tok.add_103_17_lut_LC_4_11_1  (
            .in0(N__18963),
            .in1(N__16120),
            .in2(N__24199),
            .in3(N__16018),
            .lcout(\tok.n6339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_adj_53_LC_4_11_2 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_53_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_53_LC_4_11_2 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \tok.i314_4_lut_adj_53_LC_4_11_2  (
            .in0(N__31470),
            .in1(N__16015),
            .in2(N__30066),
            .in3(N__34266),
            .lcout(\tok.n161_adj_667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_4_lut_LC_4_11_3 .C_ON=1'b0;
    defparam \tok.i2_3_lut_4_lut_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_4_lut_LC_4_11_3 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \tok.i2_3_lut_4_lut_LC_4_11_3  (
            .in0(N__34265),
            .in1(N__35715),
            .in2(N__36980),
            .in3(N__32695),
            .lcout(\tok.n260_adj_717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_284_LC_4_11_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_284_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_284_LC_4_11_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i1_4_lut_adj_284_LC_4_11_4  (
            .in0(N__30043),
            .in1(N__18835),
            .in2(N__25984),
            .in3(N__30531),
            .lcout(\tok.n17_adj_853 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_1_lut_LC_4_11_5 .C_ON=1'b0;
    defparam \tok.i7_1_lut_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i7_1_lut_LC_4_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.i7_1_lut_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32694),
            .lcout(\tok.n21_adj_660 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_LC_4_11_6 .C_ON=1'b0;
    defparam \tok.i2_2_lut_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_LC_4_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i2_2_lut_LC_4_11_6  (
            .in0(N__31469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34264),
            .lcout(\tok.n4_adj_635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i402_1_lut_LC_4_11_7 .C_ON=1'b0;
    defparam \tok.i402_1_lut_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i402_1_lut_LC_4_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.i402_1_lut_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31468),
            .lcout(\tok.n83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_248_LC_4_12_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_248_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_248_LC_4_12_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_248_LC_4_12_0  (
            .in0(N__20341),
            .in1(N__24288),
            .in2(N__17266),
            .in3(N__17155),
            .lcout(\tok.n248_adj_827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i299_4_lut_adj_267_LC_4_12_1 .C_ON=1'b0;
    defparam \tok.i299_4_lut_adj_267_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i299_4_lut_adj_267_LC_4_12_1 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \tok.i299_4_lut_adj_267_LC_4_12_1  (
            .in0(N__35716),
            .in1(N__16087),
            .in2(N__17119),
            .in3(N__32779),
            .lcout(),
            .ltout(\tok.n197_adj_837_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_268_LC_4_12_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_268_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_268_LC_4_12_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_268_LC_4_12_2  (
            .in0(N__20342),
            .in1(N__24289),
            .in2(N__16075),
            .in3(N__21761),
            .lcout(\tok.n248_adj_838 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6699_4_lut_LC_4_12_3 .C_ON=1'b0;
    defparam \tok.i6699_4_lut_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6699_4_lut_LC_4_12_3 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \tok.i6699_4_lut_LC_4_12_3  (
            .in0(N__23731),
            .in1(N__20396),
            .in2(N__35874),
            .in3(N__16900),
            .lcout(),
            .ltout(\tok.n6386_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i299_4_lut_adj_42_LC_4_12_4 .C_ON=1'b0;
    defparam \tok.i299_4_lut_adj_42_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i299_4_lut_adj_42_LC_4_12_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \tok.i299_4_lut_adj_42_LC_4_12_4  (
            .in0(N__32780),
            .in1(N__16060),
            .in2(N__16048),
            .in3(N__35721),
            .lcout(),
            .ltout(\tok.n197_adj_652_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_43_LC_4_12_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_43_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_43_LC_4_12_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_43_LC_4_12_5  (
            .in0(N__24290),
            .in1(N__20343),
            .in2(N__16045),
            .in3(N__17319),
            .lcout(\tok.n248_adj_653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6706_4_lut_LC_4_12_6 .C_ON=1'b0;
    defparam \tok.i6706_4_lut_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6706_4_lut_LC_4_12_6 .LUT_INIT=16'b0010000011100000;
    LogicCell40 \tok.i6706_4_lut_LC_4_12_6  (
            .in0(N__17068),
            .in1(N__35717),
            .in2(N__20412),
            .in3(N__23730),
            .lcout(\tok.n6356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i335_rep_143_2_lut_LC_4_12_7 .C_ON=1'b0;
    defparam \tok.i335_rep_143_2_lut_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i335_rep_143_2_lut_LC_4_12_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.i335_rep_143_2_lut_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(N__32778),
            .in2(_gnd_net_),
            .in3(N__30714),
            .lcout(\tok.n7269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_100_i12_2_lut_LC_4_13_0 .C_ON=1'b0;
    defparam \tok.or_100_i12_2_lut_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.or_100_i12_2_lut_LC_4_13_0 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \tok.or_100_i12_2_lut_LC_4_13_0  (
            .in0(N__20785),
            .in1(N__37445),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n228 ),
            .ltout(\tok.n228_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i312_4_lut_adj_320_LC_4_13_1 .C_ON=1'b0;
    defparam \tok.i312_4_lut_adj_320_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i312_4_lut_adj_320_LC_4_13_1 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \tok.i312_4_lut_adj_320_LC_4_13_1  (
            .in0(N__30719),
            .in1(N__16180),
            .in2(N__16168),
            .in3(N__32787),
            .lcout(),
            .ltout(\tok.n203_adj_879_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_321_LC_4_13_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_321_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_321_LC_4_13_2 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \tok.i1_4_lut_adj_321_LC_4_13_2  (
            .in0(N__31743),
            .in1(N__19214),
            .in2(N__16165),
            .in3(N__16162),
            .lcout(),
            .ltout(\tok.n212_adj_880_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6911_4_lut_LC_4_13_3 .C_ON=1'b0;
    defparam \tok.i6911_4_lut_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6911_4_lut_LC_4_13_3 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i6911_4_lut_LC_4_13_3  (
            .in0(N__31548),
            .in1(N__33490),
            .in2(N__16156),
            .in3(N__16126),
            .lcout(\tok.n6412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6719_3_lut_4_lut_LC_4_13_4 .C_ON=1'b0;
    defparam \tok.i6719_3_lut_4_lut_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6719_3_lut_4_lut_LC_4_13_4 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \tok.i6719_3_lut_4_lut_LC_4_13_4  (
            .in0(N__34271),
            .in1(N__30718),
            .in2(N__20792),
            .in3(N__37444),
            .lcout(\tok.n6417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_adj_76_LC_4_13_5 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_76_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_76_LC_4_13_5 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \tok.i314_4_lut_adj_76_LC_4_13_5  (
            .in0(N__31549),
            .in1(N__16153),
            .in2(N__37469),
            .in3(N__34272),
            .lcout(),
            .ltout(\tok.n161_adj_692_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i299_4_lut_adj_77_LC_4_13_6 .C_ON=1'b0;
    defparam \tok.i299_4_lut_adj_77_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.i299_4_lut_adj_77_LC_4_13_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \tok.i299_4_lut_adj_77_LC_4_13_6  (
            .in0(N__32788),
            .in1(N__36142),
            .in2(N__16144),
            .in3(N__16141),
            .lcout(\tok.n197_adj_693 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i300_4_lut_adj_322_LC_4_13_7 .C_ON=1'b0;
    defparam \tok.i300_4_lut_adj_322_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.i300_4_lut_adj_322_LC_4_13_7 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \tok.i300_4_lut_adj_322_LC_4_13_7  (
            .in0(N__20690),
            .in1(N__20610),
            .in2(N__36283),
            .in3(N__16132),
            .lcout(\tok.n206_adj_881 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2579_2_lut_LC_4_14_3 .C_ON=1'b0;
    defparam \tok.i2579_2_lut_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2579_2_lut_LC_4_14_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i2579_2_lut_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__33936),
            .in2(_gnd_net_),
            .in3(N__36548),
            .lcout(\tok.n2602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_327_LC_4_14_7 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_327_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_327_LC_4_14_7 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \tok.i308_4_lut_adj_327_LC_4_14_7  (
            .in0(N__30072),
            .in1(N__36852),
            .in2(N__26226),
            .in3(N__16267),
            .lcout(\tok.n242_adj_885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i103_LC_5_1_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i103_LC_5_1_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i103_LC_5_1_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i103_LC_5_1_0  (
            .in0(N__16261),
            .in1(N__16227),
            .in2(_gnd_net_),
            .in3(N__18451),
            .lcout(tail_103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38439),
            .ce(N__17947),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i87_LC_5_1_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i87_LC_5_1_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i87_LC_5_1_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i87_LC_5_1_1  (
            .in0(N__18457),
            .in1(N__16239),
            .in2(_gnd_net_),
            .in3(N__16218),
            .lcout(\tok.A_stk.tail_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38439),
            .ce(N__17947),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i71_LC_5_1_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i71_LC_5_1_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i71_LC_5_1_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.A_stk.tail_i0_i71_LC_5_1_2  (
            .in0(N__16209),
            .in1(N__16228),
            .in2(_gnd_net_),
            .in3(N__18455),
            .lcout(\tok.A_stk.tail_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38439),
            .ce(N__17947),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i55_LC_5_1_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i55_LC_5_1_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i55_LC_5_1_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.A_stk.tail_i0_i55_LC_5_1_3  (
            .in0(N__18454),
            .in1(N__16219),
            .in2(_gnd_net_),
            .in3(N__16200),
            .lcout(\tok.A_stk.tail_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38439),
            .ce(N__17947),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i39_LC_5_1_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i39_LC_5_1_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i39_LC_5_1_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.tail_i0_i39_LC_5_1_4  (
            .in0(N__16210),
            .in1(N__16191),
            .in2(_gnd_net_),
            .in3(N__18453),
            .lcout(\tok.A_stk.tail_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38439),
            .ce(N__17947),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i23_LC_5_1_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i23_LC_5_1_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i23_LC_5_1_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.A_stk.tail_i0_i23_LC_5_1_5  (
            .in0(N__18452),
            .in1(_gnd_net_),
            .in2(N__16408),
            .in3(N__16201),
            .lcout(\tok.A_stk.tail_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38439),
            .ce(N__17947),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i7_LC_5_1_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i7_LC_5_1_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i7_LC_5_1_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i7_LC_5_1_6  (
            .in0(N__16192),
            .in1(N__18456),
            .in2(_gnd_net_),
            .in3(N__28297),
            .lcout(\tok.A_stk.tail_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38439),
            .ce(N__17947),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i7_LC_5_1_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i7_LC_5_1_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i7_LC_5_1_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i7_LC_5_1_7  (
            .in0(N__16404),
            .in1(N__18562),
            .in2(_gnd_net_),
            .in3(N__37477),
            .lcout(\tok.S_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38439),
            .ce(N__17947),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i113_LC_5_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i113_LC_5_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i113_LC_5_2_0 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \tok.A_stk.tail_i0_i113_LC_5_2_0  (
            .in0(N__18373),
            .in1(N__16377),
            .in2(N__16396),
            .in3(N__17902),
            .lcout(tail_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38444),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i124_LC_5_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i124_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i124_LC_5_2_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \tok.A_stk.tail_i0_i124_LC_5_2_1  (
            .in0(N__17903),
            .in1(N__16366),
            .in2(N__16354),
            .in3(N__18374),
            .lcout(tail_124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38444),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.S_15__I_0_i4_3_lut_LC_5_2_2 .C_ON=1'b0;
    defparam \tok.S_15__I_0_i4_3_lut_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \tok.S_15__I_0_i4_3_lut_LC_5_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.S_15__I_0_i4_3_lut_LC_5_2_2  (
            .in0(N__23218),
            .in1(N__22646),
            .in2(_gnd_net_),
            .in3(N__28476),
            .lcout(\tok.table_wr_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1379_3_lut_LC_5_2_3.C_ON=1'b0;
    defparam i1379_3_lut_LC_5_2_3.SEQ_MODE=4'b0000;
    defparam i1379_3_lut_LC_5_2_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 i1379_3_lut_LC_5_2_3 (
            .in0(N__28475),
            .in1(N__24986),
            .in2(_gnd_net_),
            .in3(N__23495),
            .lcout(table_wr_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1464_3_lut_LC_5_2_4 .C_ON=1'b0;
    defparam \tok.ram.i1464_3_lut_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1464_3_lut_LC_5_2_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.ram.i1464_3_lut_LC_5_2_4  (
            .in0(N__27738),
            .in1(N__28477),
            .in2(_gnd_net_),
            .in3(N__25936),
            .lcout(\tok.table_wr_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1536_3_lut_LC_5_2_6 .C_ON=1'b0;
    defparam \tok.ram.i1536_3_lut_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1536_3_lut_LC_5_2_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.ram.i1536_3_lut_LC_5_2_6  (
            .in0(N__23851),
            .in1(N__21057),
            .in2(_gnd_net_),
            .in3(N__28478),
            .lcout(\tok.table_wr_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1572_3_lut_LC_5_2_7 .C_ON=1'b0;
    defparam \tok.ram.i1572_3_lut_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1572_3_lut_LC_5_2_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.ram.i1572_3_lut_LC_5_2_7  (
            .in0(N__28479),
            .in1(N__22487),
            .in2(_gnd_net_),
            .in3(N__20094),
            .lcout(\tok.table_wr_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6634_4_lut_LC_5_3_0 .C_ON=1'b0;
    defparam \tok.ram.i6634_4_lut_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6634_4_lut_LC_5_3_0 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \tok.ram.i6634_4_lut_LC_5_3_0  (
            .in0(N__22939),
            .in1(N__22875),
            .in2(N__27685),
            .in3(N__27736),
            .lcout(),
            .ltout(\tok.ram.n6266_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1456_4_lut_LC_5_3_1 .C_ON=1'b0;
    defparam \tok.ram.i1456_4_lut_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1456_4_lut_LC_5_3_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.ram.i1456_4_lut_LC_5_3_1  (
            .in0(N__22807),
            .in1(N__27684),
            .in2(N__16459),
            .in3(N__31934),
            .lcout(),
            .ltout(\tok.n1495_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_167_LC_5_3_2 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_167_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_167_LC_5_3_2 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i27_4_lut_adj_167_LC_5_3_2  (
            .in0(N__16417),
            .in1(N__35522),
            .in2(N__16456),
            .in3(N__31331),
            .lcout(\tok.n13_adj_766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i6_LC_5_3_3 .C_ON=1'b0;
    defparam \tok.tc_i6_LC_5_3_3 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i6_LC_5_3_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.tc_i6_LC_5_3_3  (
            .in0(N__16447),
            .in1(N__27707),
            .in2(_gnd_net_),
            .in3(N__19738),
            .lcout(tc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38448),
            .ce(),
            .sr(N__29220));
    defparam \tok.i1_4_lut_adj_168_LC_5_3_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_168_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_168_LC_5_3_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_168_LC_5_3_4  (
            .in0(N__25809),
            .in1(N__16453),
            .in2(N__29725),
            .in3(N__27737),
            .lcout(n10_adj_907),
            .ltout(n10_adj_907_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_200_LC_5_3_5 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_200_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_200_LC_5_3_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \tok.i26_3_lut_adj_200_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(N__27706),
            .in2(N__16441),
            .in3(N__19737),
            .lcout(\tok.tc_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_164_LC_5_3_6 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_164_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_164_LC_5_3_6 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_164_LC_5_3_6  (
            .in0(N__27680),
            .in1(N__33295),
            .in2(N__24060),
            .in3(N__31330),
            .lcout(),
            .ltout(\tok.n83_adj_765_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6725_2_lut_3_lut_LC_5_3_7 .C_ON=1'b0;
    defparam \tok.i6725_2_lut_3_lut_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6725_2_lut_3_lut_LC_5_3_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \tok.i6725_2_lut_3_lut_LC_5_3_7  (
            .in0(N__36306),
            .in1(_gnd_net_),
            .in2(N__16420),
            .in3(N__31933),
            .lcout(\tok.n6435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6614_4_lut_LC_5_4_0 .C_ON=1'b0;
    defparam \tok.i6614_4_lut_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6614_4_lut_LC_5_4_0 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \tok.i6614_4_lut_LC_5_4_0  (
            .in0(N__22945),
            .in1(N__21102),
            .in2(N__21167),
            .in3(N__22864),
            .lcout(),
            .ltout(\tok.n6283_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i124_4_lut_LC_5_4_1 .C_ON=1'b0;
    defparam \tok.i124_4_lut_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.i124_4_lut_LC_5_4_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.i124_4_lut_LC_5_4_1  (
            .in0(N__22806),
            .in1(N__21101),
            .in2(N__16411),
            .in3(N__32022),
            .lcout(),
            .ltout(\tok.n80_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i126_4_lut_LC_5_4_2 .C_ON=1'b0;
    defparam \tok.i126_4_lut_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i126_4_lut_LC_5_4_2 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i126_4_lut_LC_5_4_2  (
            .in0(N__16534),
            .in1(N__35504),
            .in2(N__16543),
            .in3(N__31252),
            .lcout(),
            .ltout(\tok.n89_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_131_LC_5_4_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_131_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_131_LC_5_4_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_131_LC_5_4_3  (
            .in0(N__29718),
            .in1(N__25805),
            .in2(N__16540),
            .in3(N__21160),
            .lcout(n92_adj_897),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_LC_5_4_4 .C_ON=1'b0;
    defparam \tok.i125_4_lut_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_LC_5_4_4 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \tok.i125_4_lut_LC_5_4_4  (
            .in0(N__16527),
            .in1(N__33137),
            .in2(N__21103),
            .in3(N__31251),
            .lcout(),
            .ltout(\tok.n83_adj_734_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6637_2_lut_3_lut_LC_5_4_5 .C_ON=1'b0;
    defparam \tok.i6637_2_lut_3_lut_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6637_2_lut_3_lut_LC_5_4_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i6637_2_lut_3_lut_LC_5_4_5  (
            .in0(_gnd_net_),
            .in1(N__36183),
            .in2(N__16537),
            .in3(N__32021),
            .lcout(\tok.n6279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i358_4_lut_LC_5_4_6 .C_ON=1'b0;
    defparam \tok.i358_4_lut_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i358_4_lut_LC_5_4_6 .LUT_INIT=16'b1010101011111100;
    LogicCell40 \tok.i358_4_lut_LC_5_4_6  (
            .in0(N__17421),
            .in1(N__33136),
            .in2(N__16528),
            .in3(N__31250),
            .lcout(\tok.n2696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2618_2_lut_LC_5_4_7 .C_ON=1'b0;
    defparam \tok.i2618_2_lut_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2618_2_lut_LC_5_4_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i2618_2_lut_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(N__28424),
            .in2(_gnd_net_),
            .in3(N__19333),
            .lcout(\tok.table_wr_data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2583_2_lut_LC_5_5_0 .C_ON=1'b0;
    defparam \tok.i2583_2_lut_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2583_2_lut_LC_5_5_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \tok.i2583_2_lut_LC_5_5_0  (
            .in0(N__28448),
            .in1(N__19514),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.table_wr_data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2542_2_lut_LC_5_5_1 .C_ON=1'b0;
    defparam \tok.i2542_2_lut_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2542_2_lut_LC_5_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i2542_2_lut_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__28447),
            .in2(_gnd_net_),
            .in3(N__20238),
            .lcout(\tok.table_wr_data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_292_LC_5_5_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_292_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_292_LC_5_5_2 .LUT_INIT=16'b0101000001110011;
    LogicCell40 \tok.i1_4_lut_adj_292_LC_5_5_2  (
            .in0(N__17422),
            .in1(N__16465),
            .in2(N__19252),
            .in3(N__32109),
            .lcout(\tok.n268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.stall_I_0_369_i11_2_lut_LC_5_5_3 .C_ON=1'b0;
    defparam \tok.stall_I_0_369_i11_2_lut_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.stall_I_0_369_i11_2_lut_LC_5_5_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.stall_I_0_369_i11_2_lut_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__31093),
            .in2(_gnd_net_),
            .in3(N__33236),
            .lcout(\tok.n9_adj_651 ),
            .ltout(\tok.n9_adj_651_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_4_lut_adj_293_LC_5_5_4 .C_ON=1'b0;
    defparam \tok.i2_2_lut_4_lut_adj_293_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_4_lut_adj_293_LC_5_5_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.i2_2_lut_4_lut_adj_293_LC_5_5_4  (
            .in0(N__30142),
            .in1(N__34643),
            .in2(N__16594),
            .in3(N__32110),
            .lcout(n15),
            .ltout(n15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_69_LC_5_5_5 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_69_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_69_LC_5_5_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \tok.i2_4_lut_adj_69_LC_5_5_5  (
            .in0(N__16591),
            .in1(N__21363),
            .in2(N__16582),
            .in3(N__19609),
            .lcout(),
            .ltout(\tok.n6_adj_687_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_71_LC_5_5_6 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_71_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_71_LC_5_5_6 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \tok.i3_4_lut_adj_71_LC_5_5_6  (
            .in0(N__30144),
            .in1(N__27923),
            .in2(N__16579),
            .in3(N__16575),
            .lcout(\tok.n2702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_4_lut_adj_275_LC_5_5_7 .C_ON=1'b0;
    defparam \tok.i2_3_lut_4_lut_adj_275_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_4_lut_adj_275_LC_5_5_7 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \tok.i2_3_lut_4_lut_adj_275_LC_5_5_7  (
            .in0(N__32108),
            .in1(N__26129),
            .in2(N__34780),
            .in3(N__30143),
            .lcout(\tok.n891 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_255_LC_5_6_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_255_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_255_LC_5_6_0 .LUT_INIT=16'b1010101010101111;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_255_LC_5_6_0  (
            .in0(N__29448),
            .in1(_gnd_net_),
            .in2(N__37241),
            .in3(N__37203),
            .lcout(\tok.uart_stall ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_257_LC_5_6_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_257_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_257_LC_5_6_1 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_257_LC_5_6_1  (
            .in0(N__37202),
            .in1(N__37230),
            .in2(_gnd_net_),
            .in3(N__29447),
            .lcout(\tok.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_33_LC_5_6_2 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_33_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_33_LC_5_6_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i1_2_lut_adj_33_LC_5_6_2  (
            .in0(N__16728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16714),
            .lcout(\tok.n6170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_4_lut_adj_312_LC_5_6_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_4_lut_adj_312_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_4_lut_adj_312_LC_5_6_3 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \tok.i1_2_lut_4_lut_adj_312_LC_5_6_3  (
            .in0(N__37234),
            .in1(N__29449),
            .in2(N__37207),
            .in3(N__16727),
            .lcout(\tok.n796 ),
            .ltout(\tok.n796_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_28_LC_5_6_4 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_28_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_28_LC_5_6_4 .LUT_INIT=16'b1111110011011100;
    LogicCell40 \tok.i2_4_lut_adj_28_LC_5_6_4  (
            .in0(N__25354),
            .in1(N__16715),
            .in2(N__16546),
            .in3(N__16794),
            .lcout(stall_),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.stall_361_LC_5_6_5 .C_ON=1'b0;
    defparam \tok.stall_361_LC_5_6_5 .SEQ_MODE=4'b1010;
    defparam \tok.stall_361_LC_5_6_5 .LUT_INIT=16'b1111111110001100;
    LogicCell40 \tok.stall_361_LC_5_6_5  (
            .in0(N__16795),
            .in1(N__16769),
            .in2(N__25358),
            .in3(N__16717),
            .lcout(\tok.stall ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38463),
            .ce(),
            .sr(N__29242));
    defparam \tok.i36_4_lut_4_lut_LC_5_6_6 .C_ON=1'b0;
    defparam \tok.i36_4_lut_4_lut_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i36_4_lut_4_lut_LC_5_6_6 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \tok.i36_4_lut_4_lut_LC_5_6_6  (
            .in0(N__16729),
            .in1(N__16716),
            .in2(N__25374),
            .in3(N__16699),
            .lcout(),
            .ltout(\tok.n31_adj_637_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_29_LC_5_6_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_29_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_29_LC_5_6_7 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \tok.i1_4_lut_adj_29_LC_5_6_7  (
            .in0(N__25325),
            .in1(N__16693),
            .in2(N__16687),
            .in3(N__16684),
            .lcout(\tok.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_276_LC_5_7_0 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_276_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_276_LC_5_7_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \tok.i4_4_lut_adj_276_LC_5_7_0  (
            .in0(N__21987),
            .in1(N__30324),
            .in2(N__23215),
            .in3(N__36454),
            .lcout(\tok.n20_adj_845 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_154_LC_5_7_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_154_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_154_LC_5_7_1 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \tok.i1_4_lut_adj_154_LC_5_7_1  (
            .in0(N__36457),
            .in1(N__25153),
            .in2(N__19870),
            .in3(N__28993),
            .lcout(),
            .ltout(\tok.n221_adj_753_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i4_LC_5_7_2 .C_ON=1'b0;
    defparam \tok.A_i4_LC_5_7_2 .SEQ_MODE=4'b1010;
    defparam \tok.A_i4_LC_5_7_2 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \tok.A_i4_LC_5_7_2  (
            .in0(N__25499),
            .in1(N__18658),
            .in2(N__16636),
            .in3(N__23209),
            .lcout(\tok.A_low_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38469),
            .ce(N__25640),
            .sr(N__29260));
    defparam \tok.i189_1_lut_LC_5_7_3 .C_ON=1'b0;
    defparam \tok.i189_1_lut_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i189_1_lut_LC_5_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.i189_1_lut_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36453),
            .lcout(\tok.n127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_LC_5_7_4 .C_ON=1'b0;
    defparam \tok.i4_4_lut_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_LC_5_7_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i4_4_lut_LC_5_7_4  (
            .in0(N__16633),
            .in1(N__30325),
            .in2(N__16615),
            .in3(N__36455),
            .lcout(),
            .ltout(\tok.n20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_35_LC_5_7_5 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_35_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_35_LC_5_7_5 .LUT_INIT=16'b1111110111111110;
    LogicCell40 \tok.i10_4_lut_adj_35_LC_5_7_5  (
            .in0(N__16885),
            .in1(N__16840),
            .in2(N__16867),
            .in3(N__22232),
            .lcout(\tok.n26_adj_645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_185_LC_5_7_6 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_185_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_185_LC_5_7_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i10_4_lut_adj_185_LC_5_7_6  (
            .in0(N__32190),
            .in1(N__30326),
            .in2(N__22249),
            .in3(N__36456),
            .lcout(\tok.n26_adj_781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.key_rd_15__I_0_401_i14_2_lut_LC_5_7_7 .C_ON=1'b0;
    defparam \tok.key_rd_15__I_0_401_i14_2_lut_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.key_rd_15__I_0_401_i14_2_lut_LC_5_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.key_rd_15__I_0_401_i14_2_lut_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(N__16855),
            .in2(_gnd_net_),
            .in3(N__32189),
            .lcout(\tok.n14_adj_644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_2_lut_LC_5_8_0 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_2_lut_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_2_lut_LC_5_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_104_add_2_2_lut_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__18865),
            .in2(N__18832),
            .in3(N__16834),
            .lcout(\tok.n308 ),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\tok.n4782 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_3_lut_LC_5_8_1 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_3_lut_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_3_lut_LC_5_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_104_add_2_3_lut_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__23374),
            .in2(N__23547),
            .in3(N__16831),
            .lcout(\tok.n307 ),
            .ltout(),
            .carryin(\tok.n4782 ),
            .carryout(\tok.n4783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_4_lut_LC_5_8_2 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_4_lut_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_4_lut_LC_5_8_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_104_add_2_4_lut_LC_5_8_2  (
            .in0(N__31898),
            .in1(N__20087),
            .in2(N__18874),
            .in3(N__16828),
            .lcout(\tok.n6616 ),
            .ltout(),
            .carryin(\tok.n4783 ),
            .carryout(\tok.n4784 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_5_lut_LC_5_8_3 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_5_lut_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_5_lut_LC_5_8_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_104_add_2_5_lut_LC_5_8_3  (
            .in0(N__33022),
            .in1(N__23211),
            .in2(N__16825),
            .in3(N__16816),
            .lcout(\tok.n2613 ),
            .ltout(),
            .carryin(\tok.n4784 ),
            .carryout(\tok.n4785 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_6_lut_LC_5_8_4 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_6_lut_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_6_lut_LC_5_8_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_104_add_2_6_lut_LC_5_8_4  (
            .in0(N__17012),
            .in1(N__20587),
            .in2(N__23852),
            .in3(N__16807),
            .lcout(\tok.n6557 ),
            .ltout(),
            .carryin(\tok.n4785 ),
            .carryout(\tok.n4786 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_7_lut_LC_5_8_5 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_7_lut_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_7_lut_LC_5_8_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_104_add_2_7_lut_LC_5_8_5  (
            .in0(N__17014),
            .in1(N__16804),
            .in2(N__22030),
            .in3(N__16798),
            .lcout(\tok.n6515 ),
            .ltout(),
            .carryin(\tok.n4786 ),
            .carryout(\tok.n4787 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_8_lut_LC_5_8_6 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_8_lut_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_8_lut_LC_5_8_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_104_add_2_8_lut_LC_5_8_6  (
            .in0(N__17011),
            .in1(N__18637),
            .in2(N__25988),
            .in3(N__17017),
            .lcout(\tok.n6491 ),
            .ltout(),
            .carryin(\tok.n4787 ),
            .carryout(\tok.n4788 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_8_THRU_CRY_0_LC_5_8_7 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_8_THRU_CRY_0_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_8_THRU_CRY_0_LC_5_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \tok.sub_104_add_2_8_THRU_CRY_0_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__17509),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\tok.n4788 ),
            .carryout(\tok.n4788_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_9_lut_LC_5_9_0 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_9_lut_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_9_lut_LC_5_9_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_104_add_2_9_lut_LC_5_9_0  (
            .in0(N__17013),
            .in1(N__28328),
            .in2(N__16981),
            .in3(N__16969),
            .lcout(\tok.n6467 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\tok.n4789 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_10_lut_LC_5_9_1 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_10_lut_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_10_lut_LC_5_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_104_add_2_10_lut_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__20500),
            .in2(N__17265),
            .in3(N__16966),
            .lcout(\tok.n300 ),
            .ltout(),
            .carryin(\tok.n4789 ),
            .carryout(\tok.n4790 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_11_lut_LC_5_9_2 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_11_lut_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_11_lut_LC_5_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_104_add_2_11_lut_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__21773),
            .in2(N__24019),
            .in3(N__16963),
            .lcout(\tok.n299 ),
            .ltout(),
            .carryin(\tok.n4790 ),
            .carryout(\tok.n4791 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_12_lut_LC_5_9_3 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_12_lut_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_12_lut_LC_5_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_104_add_2_12_lut_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__20180),
            .in2(N__16960),
            .in3(N__16948),
            .lcout(\tok.n298 ),
            .ltout(),
            .carryin(\tok.n4791 ),
            .carryout(\tok.n4792 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_13_lut_LC_5_9_4 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_13_lut_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_13_lut_LC_5_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_104_add_2_13_lut_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__19504),
            .in2(N__20614),
            .in3(N__16945),
            .lcout(\tok.n297 ),
            .ltout(),
            .carryin(\tok.n4792 ),
            .carryout(\tok.n4793 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_14_lut_LC_5_9_5 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_14_lut_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_14_lut_LC_5_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_104_add_2_14_lut_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(N__20248),
            .in2(N__16942),
            .in3(N__16930),
            .lcout(\tok.n296 ),
            .ltout(),
            .carryin(\tok.n4793 ),
            .carryout(\tok.n4794 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_15_lut_LC_5_9_6 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_15_lut_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_15_lut_LC_5_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_104_add_2_15_lut_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__17318),
            .in2(N__16926),
            .in3(N__16888),
            .lcout(\tok.n295 ),
            .ltout(),
            .carryin(\tok.n4794 ),
            .carryout(\tok.n4795 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_16_lut_LC_5_9_7 .C_ON=1'b1;
    defparam \tok.sub_104_add_2_16_lut_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_16_lut_LC_5_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_104_add_2_16_lut_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__19321),
            .in2(N__32274),
            .in3(N__17074),
            .lcout(\tok.n294 ),
            .ltout(),
            .carryin(\tok.n4795 ),
            .carryout(\tok.n4796 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_104_add_2_17_lut_LC_5_10_0 .C_ON=1'b0;
    defparam \tok.sub_104_add_2_17_lut_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_104_add_2_17_lut_LC_5_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \tok.sub_104_add_2_17_lut_LC_5_10_0  (
            .in0(N__18955),
            .in1(N__17053),
            .in2(_gnd_net_),
            .in3(N__17071),
            .lcout(\tok.n293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6717_4_lut_LC_5_10_1 .C_ON=1'b0;
    defparam \tok.i6717_4_lut_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6717_4_lut_LC_5_10_1 .LUT_INIT=16'b0010000011100000;
    LogicCell40 \tok.i6717_4_lut_LC_5_10_1  (
            .in0(N__17059),
            .in1(N__36010),
            .in2(N__20406),
            .in3(N__23720),
            .lcout(\tok.n6415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i16_1_lut_LC_5_10_2 .C_ON=1'b0;
    defparam \tok.inv_105_i16_1_lut_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i16_1_lut_LC_5_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i16_1_lut_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24143),
            .lcout(\tok.n310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_adj_246_LC_5_10_3 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_246_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_246_LC_5_10_3 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \tok.i314_4_lut_adj_246_LC_5_10_3  (
            .in0(N__31912),
            .in1(N__17047),
            .in2(N__34711),
            .in3(N__30487),
            .lcout(\tok.n161_adj_825 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i356_4_lut_LC_5_10_4 .C_ON=1'b0;
    defparam \tok.i356_4_lut_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i356_4_lut_LC_5_10_4 .LUT_INIT=16'b0100011101000100;
    LogicCell40 \tok.i356_4_lut_LC_5_10_4  (
            .in0(N__17041),
            .in1(N__34551),
            .in2(N__37747),
            .in3(N__31913),
            .lcout(\tok.n208_adj_857 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_LC_5_10_5 .C_ON=1'b0;
    defparam \tok.i314_4_lut_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_LC_5_10_5 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \tok.i314_4_lut_LC_5_10_5  (
            .in0(N__31915),
            .in1(N__17035),
            .in2(N__34712),
            .in3(N__27370),
            .lcout(\tok.n161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_adj_305_LC_5_10_6 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_305_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_305_LC_5_10_6 .LUT_INIT=16'b1010110010100000;
    LogicCell40 \tok.i314_4_lut_adj_305_LC_5_10_6  (
            .in0(N__17029),
            .in1(N__33582),
            .in2(N__34713),
            .in3(N__31914),
            .lcout(\tok.n161_adj_870 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6746_4_lut_LC_5_10_7 .C_ON=1'b0;
    defparam \tok.i6746_4_lut_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6746_4_lut_LC_5_10_7 .LUT_INIT=16'b0010000011100000;
    LogicCell40 \tok.i6746_4_lut_LC_5_10_7  (
            .in0(N__17023),
            .in1(N__36009),
            .in2(N__20405),
            .in3(N__23719),
            .lcout(\tok.n6460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i299_4_lut_adj_247_LC_5_11_0 .C_ON=1'b0;
    defparam \tok.i299_4_lut_adj_247_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i299_4_lut_adj_247_LC_5_11_0 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \tok.i299_4_lut_adj_247_LC_5_11_0  (
            .in0(N__17170),
            .in1(N__35831),
            .in2(N__17164),
            .in3(N__33234),
            .lcout(\tok.n197_adj_826 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_103_LC_5_11_1 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_103_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_103_LC_5_11_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.i1_3_lut_adj_103_LC_5_11_1  (
            .in0(N__36780),
            .in1(N__31765),
            .in2(_gnd_net_),
            .in3(N__34528),
            .lcout(\tok.n4_adj_711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i15_4_lut_adj_285_LC_5_11_2 .C_ON=1'b0;
    defparam \tok.i15_4_lut_adj_285_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i15_4_lut_adj_285_LC_5_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i15_4_lut_adj_285_LC_5_11_2  (
            .in0(N__17149),
            .in1(N__17137),
            .in2(N__18886),
            .in3(N__17179),
            .lcout(\tok.n31 ),
            .ltout(\tok.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6736_4_lut_LC_5_11_3 .C_ON=1'b0;
    defparam \tok.i6736_4_lut_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6736_4_lut_LC_5_11_3 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \tok.i6736_4_lut_LC_5_11_3  (
            .in0(N__35829),
            .in1(N__20400),
            .in2(N__17131),
            .in3(N__17128),
            .lcout(\tok.n6446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6667_4_lut_LC_5_11_4 .C_ON=1'b0;
    defparam \tok.i6667_4_lut_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6667_4_lut_LC_5_11_4 .LUT_INIT=16'b1101000000010000;
    LogicCell40 \tok.i6667_4_lut_LC_5_11_4  (
            .in0(N__17110),
            .in1(N__35830),
            .in2(N__20416),
            .in3(N__23726),
            .lcout(\tok.n6328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6688_4_lut_LC_5_11_5 .C_ON=1'b0;
    defparam \tok.i6688_4_lut_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6688_4_lut_LC_5_11_5 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \tok.i6688_4_lut_LC_5_11_5  (
            .in0(N__23727),
            .in1(N__20404),
            .in2(N__36031),
            .in3(N__17101),
            .lcout(),
            .ltout(\tok.n6371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i299_4_lut_adj_54_LC_5_11_6 .C_ON=1'b0;
    defparam \tok.i299_4_lut_adj_54_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i299_4_lut_adj_54_LC_5_11_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.i299_4_lut_adj_54_LC_5_11_6  (
            .in0(N__17092),
            .in1(N__35835),
            .in2(N__17086),
            .in3(N__33235),
            .lcout(\tok.n197_adj_668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_172_LC_5_11_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_172_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_172_LC_5_11_7 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_172_LC_5_11_7  (
            .in0(N__35828),
            .in1(_gnd_net_),
            .in2(N__36935),
            .in3(N__34527),
            .lcout(\tok.n4_adj_680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_45_LC_5_12_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_45_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_45_LC_5_12_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_45_LC_5_12_0  (
            .in0(N__37083),
            .in1(N__35206),
            .in2(N__17083),
            .in3(N__17326),
            .lcout(),
            .ltout(\tok.n200_adj_655_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_48_LC_5_12_1 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_48_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_48_LC_5_12_1 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \tok.i2_4_lut_adj_48_LC_5_12_1  (
            .in0(N__26611),
            .in1(N__32188),
            .in2(N__17350),
            .in3(N__33935),
            .lcout(),
            .ltout(\tok.n6_adj_658_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i14_LC_5_12_2 .C_ON=1'b0;
    defparam \tok.A_i14_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \tok.A_i14_LC_5_12_2 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \tok.A_i14_LC_5_12_2  (
            .in0(N__25517),
            .in1(N__24484),
            .in2(N__17347),
            .in3(N__17314),
            .lcout(\tok.n44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38489),
            .ce(N__25650),
            .sr(N__29269));
    defparam \tok.i2_4_lut_adj_254_LC_5_12_3 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_254_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_254_LC_5_12_3 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \tok.i2_4_lut_adj_254_LC_5_12_3  (
            .in0(N__22189),
            .in1(N__33934),
            .in2(N__26617),
            .in3(N__19396),
            .lcout(),
            .ltout(\tok.n6_adj_832_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i9_LC_5_12_4 .C_ON=1'b0;
    defparam \tok.A_i9_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \tok.A_i9_LC_5_12_4 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \tok.A_i9_LC_5_12_4  (
            .in0(N__25518),
            .in1(N__20824),
            .in2(N__17344),
            .in3(N__17251),
            .lcout(\tok.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38489),
            .ce(N__25650),
            .sr(N__29269));
    defparam \tok.i308_4_lut_adj_44_LC_5_12_5 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_44_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_44_LC_5_12_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \tok.i308_4_lut_adj_44_LC_5_12_5  (
            .in0(N__22188),
            .in1(N__37082),
            .in2(N__26222),
            .in3(N__17341),
            .lcout(\tok.n242_adj_654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_106_i14_2_lut_LC_5_12_6 .C_ON=1'b0;
    defparam \tok.equal_106_i14_2_lut_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.equal_106_i14_2_lut_LC_5_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.equal_106_i14_2_lut_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__32169),
            .in2(_gnd_net_),
            .in3(N__17313),
            .lcout(),
            .ltout(\tok.n14_adj_844_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_282_LC_5_12_7 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_282_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_282_LC_5_12_7 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \tok.i10_4_lut_adj_282_LC_5_12_7  (
            .in0(N__17250),
            .in1(N__22167),
            .in2(N__17191),
            .in3(N__17188),
            .lcout(\tok.n26_adj_851 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6663_3_lut_4_lut_LC_5_13_1 .C_ON=1'b0;
    defparam \tok.i6663_3_lut_4_lut_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6663_3_lut_4_lut_LC_5_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \tok.i6663_3_lut_4_lut_LC_5_13_1  (
            .in0(N__34558),
            .in1(N__36030),
            .in2(N__30534),
            .in3(N__33100),
            .lcout(),
            .ltout(\tok.n6324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i366_4_lut_LC_5_13_2 .C_ON=1'b0;
    defparam \tok.i366_4_lut_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i366_4_lut_LC_5_13_2 .LUT_INIT=16'b1010000010110001;
    LogicCell40 \tok.i366_4_lut_LC_5_13_2  (
            .in0(N__30859),
            .in1(N__33431),
            .in2(N__17173),
            .in3(N__17414),
            .lcout(),
            .ltout(\tok.n262_adj_858_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6669_4_lut_LC_5_13_3 .C_ON=1'b0;
    defparam \tok.i6669_4_lut_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6669_4_lut_LC_5_13_3 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \tok.i6669_4_lut_LC_5_13_3  (
            .in0(N__31916),
            .in1(N__33432),
            .in2(N__17563),
            .in3(N__17560),
            .lcout(\tok.n6315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_13_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_13_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_13_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(CONSTANT_ONE_NET_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_99_add_2_2_lut_LC_5_13_5 .C_ON=1'b0;
    defparam \tok.sub_99_add_2_2_lut_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_99_add_2_2_lut_LC_5_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_99_add_2_2_lut_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17425),
            .in3(N__30858),
            .lcout(\tok.n239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i3_LC_5_13_7 .C_ON=1'b0;
    defparam \tok.uart.sender_i3_LC_5_13_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i3_LC_5_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.uart.sender_i3_LC_5_13_7  (
            .in0(N__30524),
            .in1(N__20863),
            .in2(_gnd_net_),
            .in3(N__37540),
            .lcout(sender_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38494),
            .ce(N__27171),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_80_LC_5_14_0 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_80_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_80_LC_5_14_0 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \tok.i308_4_lut_adj_80_LC_5_14_0  (
            .in0(N__29618),
            .in1(N__37077),
            .in2(N__26227),
            .in3(N__17380),
            .lcout(\tok.n242_adj_695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_79_LC_5_14_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_79_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_79_LC_5_14_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_79_LC_5_14_1  (
            .in0(N__24328),
            .in1(N__20344),
            .in2(N__18973),
            .in3(N__17368),
            .lcout(),
            .ltout(\tok.n248_adj_694_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_81_LC_5_14_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_81_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_81_LC_5_14_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_81_LC_5_14_2  (
            .in0(N__35266),
            .in1(N__37078),
            .in2(N__17362),
            .in3(N__17359),
            .lcout(),
            .ltout(\tok.n200_adj_696_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_84_LC_5_14_3 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_84_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_84_LC_5_14_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \tok.i2_4_lut_adj_84_LC_5_14_3  (
            .in0(N__33994),
            .in1(N__26609),
            .in2(N__17353),
            .in3(N__24133),
            .lcout(),
            .ltout(\tok.n6_adj_699_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i16_LC_5_14_4 .C_ON=1'b0;
    defparam \tok.A_i16_LC_5_14_4 .SEQ_MODE=4'b1010;
    defparam \tok.A_i16_LC_5_14_4 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \tok.A_i16_LC_5_14_4  (
            .in0(N__25519),
            .in1(N__18972),
            .in2(N__17584),
            .in3(N__20908),
            .lcout(\tok.n42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38499),
            .ce(N__25642),
            .sr(N__29272));
    defparam \tok.i6872_2_lut_3_lut_4_lut_LC_5_14_5 .C_ON=1'b0;
    defparam \tok.i6872_2_lut_3_lut_4_lut_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6872_2_lut_3_lut_4_lut_LC_5_14_5 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \tok.i6872_2_lut_3_lut_4_lut_LC_5_14_5  (
            .in0(N__37076),
            .in1(N__24426),
            .in2(N__34080),
            .in3(N__29617),
            .lcout(\tok.n6367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6865_2_lut_3_lut_4_lut_LC_5_14_6 .C_ON=1'b0;
    defparam \tok.i6865_2_lut_3_lut_4_lut_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6865_2_lut_3_lut_4_lut_LC_5_14_6 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \tok.i6865_2_lut_3_lut_4_lut_LC_5_14_6  (
            .in0(N__27362),
            .in1(N__33987),
            .in2(N__24453),
            .in3(N__37075),
            .lcout(\tok.n6456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6869_2_lut_3_lut_4_lut_LC_5_14_7 .C_ON=1'b0;
    defparam \tok.i6869_2_lut_3_lut_4_lut_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6869_2_lut_3_lut_4_lut_LC_5_14_7 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \tok.i6869_2_lut_3_lut_4_lut_LC_5_14_7  (
            .in0(N__37074),
            .in1(N__24425),
            .in2(N__34079),
            .in3(N__37470),
            .lcout(\tok.n6411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_404_2_lut_LC_6_2_0 .C_ON=1'b1;
    defparam \tok.add_404_2_lut_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_404_2_lut_LC_6_2_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.add_404_2_lut_LC_6_2_0  (
            .in0(_gnd_net_),
            .in1(N__21124),
            .in2(_gnd_net_),
            .in3(N__17581),
            .lcout(tc_plus_1_0),
            .ltout(),
            .carryin(bfn_6_2_0_),
            .carryout(\tok.n4812 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_404_3_lut_LC_6_2_1 .C_ON=1'b1;
    defparam \tok.add_404_3_lut_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_404_3_lut_LC_6_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.add_404_3_lut_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(N__24955),
            .in2(_gnd_net_),
            .in3(N__17578),
            .lcout(tc_plus_1_1),
            .ltout(),
            .carryin(\tok.n4812 ),
            .carryout(\tok.n4813 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_404_4_lut_LC_6_2_2 .C_ON=1'b1;
    defparam \tok.add_404_4_lut_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_404_4_lut_LC_6_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.add_404_4_lut_LC_6_2_2  (
            .in0(_gnd_net_),
            .in1(N__22456),
            .in2(_gnd_net_),
            .in3(N__17575),
            .lcout(\tok.tc_plus_1_2 ),
            .ltout(),
            .carryin(\tok.n4813 ),
            .carryout(\tok.n4814 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_404_5_lut_LC_6_2_3 .C_ON=1'b1;
    defparam \tok.add_404_5_lut_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_404_5_lut_LC_6_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.add_404_5_lut_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(N__22606),
            .in2(_gnd_net_),
            .in3(N__17572),
            .lcout(\tok.tc_plus_1_3 ),
            .ltout(),
            .carryin(\tok.n4814 ),
            .carryout(\tok.n4815 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_404_6_lut_LC_6_2_4 .C_ON=1'b1;
    defparam \tok.add_404_6_lut_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_404_6_lut_LC_6_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.add_404_6_lut_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(N__21028),
            .in2(_gnd_net_),
            .in3(N__17569),
            .lcout(\tok.tc_plus_1_4 ),
            .ltout(),
            .carryin(\tok.n4815 ),
            .carryout(\tok.n4816 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_404_7_lut_LC_6_2_5 .C_ON=1'b1;
    defparam \tok.add_404_7_lut_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_404_7_lut_LC_6_2_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.add_404_7_lut_LC_6_2_5  (
            .in0(_gnd_net_),
            .in1(N__22306),
            .in2(_gnd_net_),
            .in3(N__17566),
            .lcout(\tok.tc_plus_1_5 ),
            .ltout(),
            .carryin(\tok.n4816 ),
            .carryout(\tok.n4817 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_404_8_lut_LC_6_2_6 .C_ON=1'b1;
    defparam \tok.add_404_8_lut_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_404_8_lut_LC_6_2_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.add_404_8_lut_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27711),
            .in3(N__17635),
            .lcout(\tok.tc_plus_1_6 ),
            .ltout(),
            .carryin(\tok.n4817 ),
            .carryout(\tok.n4818 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_404_9_lut_LC_6_2_7 .C_ON=1'b0;
    defparam \tok.add_404_9_lut_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_404_9_lut_LC_6_2_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.add_404_9_lut_LC_6_2_7  (
            .in0(_gnd_net_),
            .in1(N__27977),
            .in2(_gnd_net_),
            .in3(N__17632),
            .lcout(\tok.tc_plus_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_162_LC_6_3_0 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_162_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_162_LC_6_3_0 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \tok.i27_4_lut_adj_162_LC_6_3_0  (
            .in0(N__31333),
            .in1(N__17602),
            .in2(N__17593),
            .in3(N__35502),
            .lcout(),
            .ltout(\tok.n13_adj_760_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_163_LC_6_3_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_163_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_163_LC_6_3_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_163_LC_6_3_1  (
            .in0(N__29711),
            .in1(N__25813),
            .in2(N__17629),
            .in3(N__22334),
            .lcout(n10_adj_905),
            .ltout(n10_adj_905_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_201_LC_6_3_2 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_201_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_201_LC_6_3_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.i26_3_lut_adj_201_LC_6_3_2  (
            .in0(N__19730),
            .in1(_gnd_net_),
            .in2(N__17626),
            .in3(N__22307),
            .lcout(\tok.tc_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6619_4_lut_LC_6_3_3 .C_ON=1'b0;
    defparam \tok.ram.i6619_4_lut_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6619_4_lut_LC_6_3_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \tok.ram.i6619_4_lut_LC_6_3_3  (
            .in0(N__22931),
            .in1(N__22333),
            .in2(N__22876),
            .in3(N__22287),
            .lcout(),
            .ltout(\tok.ram.n6263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1492_4_lut_LC_6_3_4 .C_ON=1'b0;
    defparam \tok.ram.i1492_4_lut_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1492_4_lut_LC_6_3_4 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.ram.i1492_4_lut_LC_6_3_4  (
            .in0(N__22288),
            .in1(N__22801),
            .in2(N__17605),
            .in3(N__31938),
            .lcout(\tok.n1530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_160_LC_6_3_5 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_160_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_160_LC_6_3_5 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \tok.i125_4_lut_adj_160_LC_6_3_5  (
            .in0(N__33101),
            .in1(N__22286),
            .in2(N__19906),
            .in3(N__31332),
            .lcout(),
            .ltout(\tok.n83_adj_759_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6973_2_lut_3_lut_LC_6_3_6 .C_ON=1'b0;
    defparam \tok.i6973_2_lut_3_lut_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6973_2_lut_3_lut_LC_6_3_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i6973_2_lut_3_lut_LC_6_3_6  (
            .in0(_gnd_net_),
            .in1(N__36324),
            .in2(N__17596),
            .in3(N__31937),
            .lcout(\tok.n6660 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i5_LC_6_3_7 .C_ON=1'b0;
    defparam \tok.tc_i5_LC_6_3_7 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i5_LC_6_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.tc_i5_LC_6_3_7  (
            .in0(N__22308),
            .in1(N__17695),
            .in2(_gnd_net_),
            .in3(N__19731),
            .lcout(tc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38452),
            .ce(),
            .sr(N__29230));
    defparam \tok.i125_4_lut_adj_195_LC_6_4_0 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_195_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_195_LC_6_4_0 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_195_LC_6_4_0  (
            .in0(N__27854),
            .in1(N__33162),
            .in2(N__21681),
            .in3(N__31324),
            .lcout(),
            .ltout(\tok.n83_adj_764_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6978_2_lut_3_lut_LC_6_4_1 .C_ON=1'b0;
    defparam \tok.i6978_2_lut_3_lut_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6978_2_lut_3_lut_LC_6_4_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i6978_2_lut_3_lut_LC_6_4_1  (
            .in0(_gnd_net_),
            .in1(N__36184),
            .in2(N__17689),
            .in3(N__32023),
            .lcout(\tok.n6662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6596_4_lut_LC_6_4_2 .C_ON=1'b0;
    defparam \tok.ram.i6596_4_lut_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6596_4_lut_LC_6_4_2 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \tok.ram.i6596_4_lut_LC_6_4_2  (
            .in0(N__28363),
            .in1(N__22944),
            .in2(N__27859),
            .in3(N__22863),
            .lcout(),
            .ltout(\tok.ram.n6277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1600_4_lut_LC_6_4_3 .C_ON=1'b0;
    defparam \tok.ram.i1600_4_lut_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1600_4_lut_LC_6_4_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.ram.i1600_4_lut_LC_6_4_3  (
            .in0(N__22802),
            .in1(N__27858),
            .in2(N__17686),
            .in3(N__32024),
            .lcout(\tok.n1635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_197_LC_6_4_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_197_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_197_LC_6_4_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_197_LC_6_4_4  (
            .in0(N__17647),
            .in1(N__29719),
            .in2(N__28373),
            .in3(N__25806),
            .lcout(n10),
            .ltout(n10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_LC_6_4_5 .C_ON=1'b0;
    defparam \tok.i26_3_lut_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_LC_6_4_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \tok.i26_3_lut_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(N__27970),
            .in2(N__17683),
            .in3(N__19728),
            .lcout(\tok.tc_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_196_LC_6_4_6 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_196_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_196_LC_6_4_6 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \tok.i27_4_lut_adj_196_LC_6_4_6  (
            .in0(N__17662),
            .in1(N__35443),
            .in2(N__17656),
            .in3(N__31325),
            .lcout(\tok.n13_adj_790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i7_LC_6_4_7 .C_ON=1'b0;
    defparam \tok.tc_i7_LC_6_4_7 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i7_LC_6_4_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.tc_i7_LC_6_4_7  (
            .in0(N__27979),
            .in1(N__17641),
            .in2(_gnd_net_),
            .in3(N__19729),
            .lcout(tc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38458),
            .ce(),
            .sr(N__29180));
    defparam \tok.i1_2_lut_adj_236_LC_6_5_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_236_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_236_LC_6_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i1_2_lut_adj_236_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__35394),
            .in2(_gnd_net_),
            .in3(N__37003),
            .lcout(\tok.n5_adj_715 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_78_LC_6_5_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_78_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_78_LC_6_5_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \tok.i1_2_lut_adj_78_LC_6_5_1  (
            .in0(N__37002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36179),
            .lcout(\tok.n5_adj_675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6962_4_lut_LC_6_5_2 .C_ON=1'b0;
    defparam \tok.i6962_4_lut_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6962_4_lut_LC_6_5_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \tok.i6962_4_lut_LC_6_5_2  (
            .in0(N__33609),
            .in1(N__35395),
            .in2(N__36294),
            .in3(N__34704),
            .lcout(\tok.n6632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_98_i7_3_lut_4_lut_LC_6_5_3 .C_ON=1'b0;
    defparam \tok.or_98_i7_3_lut_4_lut_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.or_98_i7_3_lut_4_lut_LC_6_5_3 .LUT_INIT=16'b1111111110000111;
    LogicCell40 \tok.or_98_i7_3_lut_4_lut_LC_6_5_3  (
            .in0(N__37001),
            .in1(N__36178),
            .in2(N__35495),
            .in3(N__33608),
            .lcout(\tok.n206_adj_794 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6121_2_lut_LC_6_5_4 .C_ON=1'b0;
    defparam \tok.i6121_2_lut_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6121_2_lut_LC_6_5_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i6121_2_lut_LC_6_5_4  (
            .in0(N__29413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31110),
            .lcout(),
            .ltout(\tok.n6205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_127_LC_6_5_5 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_127_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_127_LC_6_5_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \tok.i4_4_lut_adj_127_LC_6_5_5  (
            .in0(N__27133),
            .in1(N__18606),
            .in2(N__18592),
            .in3(N__26260),
            .lcout(\tok.n270 ),
            .ltout(\tok.n270_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i2_LC_6_5_6 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i2_LC_6_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i2_LC_6_5_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \tok.A_stk.head_i0_i2_LC_6_5_6  (
            .in0(N__33610),
            .in1(_gnd_net_),
            .in2(N__18481),
            .in3(N__17967),
            .lcout(\tok.S_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38464),
            .ce(N__17956),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i2_LC_6_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i2_LC_6_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i2_LC_6_5_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.tail_i0_i2_LC_6_5_7  (
            .in0(N__18478),
            .in1(N__18254),
            .in2(_gnd_net_),
            .in3(N__20076),
            .lcout(\tok.A_stk.tail_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38464),
            .ce(N__17956),
            .sr(_gnd_net_));
    defparam \tok.i339_4_lut_LC_6_6_0 .C_ON=1'b0;
    defparam \tok.i339_4_lut_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i339_4_lut_LC_6_6_0 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \tok.i339_4_lut_LC_6_6_0  (
            .in0(N__22984),
            .in1(N__21310),
            .in2(N__23458),
            .in3(N__36950),
            .lcout(),
            .ltout(\tok.n283_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i347_4_lut_LC_6_6_1 .C_ON=1'b0;
    defparam \tok.i347_4_lut_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i347_4_lut_LC_6_6_1 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \tok.i347_4_lut_LC_6_6_1  (
            .in0(N__21394),
            .in1(N__26317),
            .in2(N__18664),
            .in3(N__35479),
            .lcout(),
            .ltout(\tok.n223_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_153_LC_6_6_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_153_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_153_LC_6_6_2 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \tok.i1_4_lut_adj_153_LC_6_6_2  (
            .in0(N__34083),
            .in1(N__36951),
            .in2(N__18661),
            .in3(N__18649),
            .lcout(\tok.n4_adj_752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6826_4_lut_LC_6_6_3 .C_ON=1'b0;
    defparam \tok.i6826_4_lut_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6826_4_lut_LC_6_6_3 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \tok.i6826_4_lut_LC_6_6_3  (
            .in0(N__20695),
            .in1(N__34082),
            .in2(N__36534),
            .in3(N__19951),
            .lcout(),
            .ltout(\tok.n6586_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i340_4_lut_LC_6_6_4 .C_ON=1'b0;
    defparam \tok.i340_4_lut_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i340_4_lut_LC_6_6_4 .LUT_INIT=16'b1111000011011101;
    LogicCell40 \tok.i340_4_lut_LC_6_6_4  (
            .in0(N__23035),
            .in1(N__18643),
            .in2(N__18652),
            .in3(N__36185),
            .lcout(\tok.n226_adj_744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_146_LC_6_6_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_146_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_146_LC_6_6_5 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \tok.i1_4_lut_adj_146_LC_6_6_5  (
            .in0(N__21415),
            .in1(N__34081),
            .in2(N__19975),
            .in3(N__35478),
            .lcout(\tok.n254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i7_1_lut_LC_6_6_7 .C_ON=1'b0;
    defparam \tok.inv_105_i7_1_lut_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i7_1_lut_LC_6_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i7_1_lut_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29931),
            .lcout(\tok.n319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6811_2_lut_3_lut_LC_6_7_0 .C_ON=1'b0;
    defparam \tok.i6811_2_lut_3_lut_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6811_2_lut_3_lut_LC_6_7_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \tok.i6811_2_lut_3_lut_LC_6_7_0  (
            .in0(N__36948),
            .in1(N__30393),
            .in2(_gnd_net_),
            .in3(N__33945),
            .lcout(\tok.n6567 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i364_4_lut_LC_6_7_1 .C_ON=1'b0;
    defparam \tok.i364_4_lut_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i364_4_lut_LC_6_7_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \tok.i364_4_lut_LC_6_7_1  (
            .in0(N__35474),
            .in1(N__18628),
            .in2(N__19141),
            .in3(N__31222),
            .lcout(),
            .ltout(\tok.n387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_296_LC_6_7_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_296_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_296_LC_6_7_2 .LUT_INIT=16'b0000000011110010;
    LogicCell40 \tok.i1_4_lut_adj_296_LC_6_7_2  (
            .in0(N__23020),
            .in1(N__18833),
            .in2(N__18616),
            .in3(N__33946),
            .lcout(),
            .ltout(\tok.n254_adj_860_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_297_LC_6_7_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_297_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_297_LC_6_7_3 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \tok.i1_4_lut_adj_297_LC_6_7_3  (
            .in0(N__21916),
            .in1(N__34705),
            .in2(N__18613),
            .in3(N__31223),
            .lcout(\tok.n256_adj_862 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i178_1_lut_LC_6_7_4 .C_ON=1'b0;
    defparam \tok.i178_1_lut_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i178_1_lut_LC_6_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.i178_1_lut_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30391),
            .lcout(\tok.n163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_303_LC_6_7_5 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_303_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_303_LC_6_7_5 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \tok.i2_4_lut_adj_303_LC_6_7_5  (
            .in0(N__30394),
            .in1(N__36949),
            .in2(N__19846),
            .in3(N__18859),
            .lcout(),
            .ltout(\tok.n6_adj_868_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i1_LC_6_7_6 .C_ON=1'b0;
    defparam \tok.A_i1_LC_6_7_6 .SEQ_MODE=4'b1010;
    defparam \tok.A_i1_LC_6_7_6 .LUT_INIT=16'b0011011100000100;
    LogicCell40 \tok.A_i1_LC_6_7_6  (
            .in0(N__18853),
            .in1(N__25482),
            .in2(N__18838),
            .in3(N__18834),
            .lcout(\tok.A_low_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38473),
            .ce(N__25639),
            .sr(N__29237));
    defparam \tok.i6804_2_lut_3_lut_LC_6_7_7 .C_ON=1'b0;
    defparam \tok.i6804_2_lut_3_lut_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6804_2_lut_3_lut_LC_6_7_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \tok.i6804_2_lut_3_lut_LC_6_7_7  (
            .in0(N__30392),
            .in1(N__36947),
            .in2(_gnd_net_),
            .in3(N__31221),
            .lcout(\tok.n6532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i12_4_lut_LC_6_8_0 .C_ON=1'b0;
    defparam \tok.i12_4_lut_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i12_4_lut_LC_6_8_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i12_4_lut_LC_6_8_0  (
            .in0(N__18705),
            .in1(N__18688),
            .in2(N__18733),
            .in3(N__18753),
            .lcout(\tok.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_LC_6_8_1 .C_ON=1'b0;
    defparam \tok.i7_4_lut_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_LC_6_8_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i7_4_lut_LC_6_8_1  (
            .in0(N__23966),
            .in1(N__32356),
            .in2(N__18754),
            .in3(N__18729),
            .lcout(\tok.n23_adj_638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_4_lut_LC_6_8_2 .C_ON=1'b0;
    defparam \tok.i8_4_lut_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i8_4_lut_LC_6_8_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i8_4_lut_LC_6_8_2  (
            .in0(N__26773),
            .in1(N__24185),
            .in2(N__18706),
            .in3(N__18687),
            .lcout(\tok.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i12_4_lut_adj_182_LC_6_8_3 .C_ON=1'b0;
    defparam \tok.i12_4_lut_adj_182_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i12_4_lut_adj_182_LC_6_8_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i12_4_lut_adj_182_LC_6_8_3  (
            .in0(N__23967),
            .in1(N__24186),
            .in2(N__32373),
            .in3(N__26774),
            .lcout(),
            .ltout(\tok.n28_adj_778_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i15_4_lut_adj_192_LC_6_8_4 .C_ON=1'b0;
    defparam \tok.i15_4_lut_adj_192_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i15_4_lut_adj_192_LC_6_8_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i15_4_lut_adj_192_LC_6_8_4  (
            .in0(N__18988),
            .in1(N__19063),
            .in2(N__18982),
            .in3(N__18979),
            .lcout(\tok.tc__7__N_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_191_LC_6_8_5 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_191_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_191_LC_6_8_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_191_LC_6_8_5  (
            .in0(N__27358),
            .in1(N__27510),
            .in2(N__30053),
            .in3(N__30410),
            .lcout(\tok.n25_adj_788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_279_LC_6_8_6 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_279_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_279_LC_6_8_6 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \tok.i7_4_lut_adj_279_LC_6_8_6  (
            .in0(N__32355),
            .in1(N__19320),
            .in2(N__19487),
            .in3(N__23965),
            .lcout(\tok.n23_adj_848 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_4_lut_adj_277_LC_6_8_7 .C_ON=1'b0;
    defparam \tok.i8_4_lut_adj_277_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i8_4_lut_adj_277_LC_6_8_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i8_4_lut_adj_277_LC_6_8_7  (
            .in0(N__24184),
            .in1(N__26772),
            .in2(N__21777),
            .in3(N__18950),
            .lcout(\tok.n24_adj_846 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i3_LC_6_9_0 .C_ON=1'b0;
    defparam \tok.A_i3_LC_6_9_0 .SEQ_MODE=4'b1010;
    defparam \tok.A_i3_LC_6_9_0 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \tok.A_i3_LC_6_9_0  (
            .in0(N__25500),
            .in1(N__18907),
            .in2(N__20090),
            .in3(N__23413),
            .lcout(\tok.A_low_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38483),
            .ce(N__25641),
            .sr(N__29117));
    defparam \tok.i6983_4_lut_LC_6_9_1 .C_ON=1'b0;
    defparam \tok.i6983_4_lut_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6983_4_lut_LC_6_9_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i6983_4_lut_LC_6_9_1  (
            .in0(N__33564),
            .in1(N__36375),
            .in2(N__19627),
            .in3(N__19591),
            .lcout(\tok.n6634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_280_LC_6_9_2 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_280_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_280_LC_6_9_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i5_4_lut_adj_280_LC_6_9_2  (
            .in0(N__20249),
            .in1(N__20179),
            .in2(N__29562),
            .in3(N__26987),
            .lcout(),
            .ltout(\tok.n21_adj_849_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i14_4_lut_adj_283_LC_6_9_3 .C_ON=1'b0;
    defparam \tok.i14_4_lut_adj_283_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i14_4_lut_adj_283_LC_6_9_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i14_4_lut_adj_283_LC_6_9_3  (
            .in0(N__18901),
            .in1(N__19069),
            .in2(N__18895),
            .in3(N__18892),
            .lcout(\tok.n30_adj_852 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i3_1_lut_LC_6_9_5 .C_ON=1'b0;
    defparam \tok.inv_105_i3_1_lut_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i3_1_lut_LC_6_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \tok.inv_105_i3_1_lut_LC_6_9_5  (
            .in0(N__33561),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_278_LC_6_9_6 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_278_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_278_LC_6_9_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i6_4_lut_adj_278_LC_6_9_6  (
            .in0(N__28298),
            .in1(N__20077),
            .in2(N__37400),
            .in3(N__33562),
            .lcout(\tok.n22_adj_847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i11_4_lut_adj_186_LC_6_9_7 .C_ON=1'b0;
    defparam \tok.i11_4_lut_adj_186_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i11_4_lut_adj_186_LC_6_9_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i11_4_lut_adj_186_LC_6_9_7  (
            .in0(N__33563),
            .in1(N__37359),
            .in2(N__27012),
            .in3(N__29529),
            .lcout(\tok.n27_adj_782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6728_4_lut_LC_6_10_0 .C_ON=1'b0;
    defparam \tok.i6728_4_lut_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6728_4_lut_LC_6_10_0 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \tok.i6728_4_lut_LC_6_10_0  (
            .in0(N__23728),
            .in1(N__20426),
            .in2(N__36213),
            .in3(N__19057),
            .lcout(),
            .ltout(\tok.n6429_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i299_4_lut_adj_307_LC_6_10_1 .C_ON=1'b0;
    defparam \tok.i299_4_lut_adj_307_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i299_4_lut_adj_307_LC_6_10_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.i299_4_lut_adj_307_LC_6_10_1  (
            .in0(N__19051),
            .in1(N__36015),
            .in2(N__19045),
            .in3(N__32960),
            .lcout(),
            .ltout(\tok.n197_adj_872_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_308_LC_6_10_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_308_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_308_LC_6_10_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_308_LC_6_10_2  (
            .in0(N__20322),
            .in1(N__24333),
            .in2(N__19042),
            .in3(N__20190),
            .lcout(\tok.n248_adj_873 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6708_4_lut_LC_6_10_3 .C_ON=1'b0;
    defparam \tok.i6708_4_lut_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6708_4_lut_LC_6_10_3 .LUT_INIT=16'b0010000011100000;
    LogicCell40 \tok.i6708_4_lut_LC_6_10_3  (
            .in0(N__19024),
            .in1(N__36014),
            .in2(N__20433),
            .in3(N__23729),
            .lcout(),
            .ltout(\tok.n6400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i299_4_lut_LC_6_10_4 .C_ON=1'b0;
    defparam \tok.i299_4_lut_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i299_4_lut_LC_6_10_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \tok.i299_4_lut_LC_6_10_4  (
            .in0(N__36016),
            .in1(N__32958),
            .in2(N__19018),
            .in3(N__19015),
            .lcout(\tok.n197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_adj_323_LC_6_10_5 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_323_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_323_LC_6_10_5 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \tok.i314_4_lut_adj_323_LC_6_10_5  (
            .in0(N__34535),
            .in1(N__36509),
            .in2(N__19009),
            .in3(N__32020),
            .lcout(),
            .ltout(\tok.n161_adj_882_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i299_4_lut_adj_324_LC_6_10_6 .C_ON=1'b0;
    defparam \tok.i299_4_lut_adj_324_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i299_4_lut_adj_324_LC_6_10_6 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \tok.i299_4_lut_adj_324_LC_6_10_6  (
            .in0(N__36018),
            .in1(N__18997),
            .in2(N__18991),
            .in3(N__32959),
            .lcout(\tok.n197_adj_883 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i363_4_lut_LC_6_10_7 .C_ON=1'b0;
    defparam \tok.i363_4_lut_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i363_4_lut_LC_6_10_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.i363_4_lut_LC_6_10_7  (
            .in0(N__19159),
            .in1(N__36017),
            .in2(N__19150),
            .in3(N__32961),
            .lcout(\tok.n250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_237_LC_6_11_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_237_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_237_LC_6_11_0 .LUT_INIT=16'b0101101001001000;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_adj_237_LC_6_11_0  (
            .in0(N__36747),
            .in1(N__32018),
            .in2(N__30499),
            .in3(N__31049),
            .lcout(\tok.n190_adj_774 ),
            .ltout(\tok.n190_adj_774_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_adj_176_LC_6_11_1 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_176_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_176_LC_6_11_1 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \tok.i314_4_lut_adj_176_LC_6_11_1  (
            .in0(N__26383),
            .in1(N__19935),
            .in2(N__19129),
            .in3(N__36748),
            .lcout(\tok.n255_adj_775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_206_LC_6_11_2 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_206_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_206_LC_6_11_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_206_LC_6_11_2  (
            .in0(N__36746),
            .in1(N__35723),
            .in2(_gnd_net_),
            .in3(N__31048),
            .lcout(\tok.n833 ),
            .ltout(\tok.n833_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6800_4_lut_LC_6_11_3 .C_ON=1'b0;
    defparam \tok.i6800_4_lut_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6800_4_lut_LC_6_11_3 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \tok.i6800_4_lut_LC_6_11_3  (
            .in0(N__32019),
            .in1(N__19126),
            .in2(N__19114),
            .in3(N__19111),
            .lcout(),
            .ltout(\tok.n6534_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i303_4_lut_adj_187_LC_6_11_4 .C_ON=1'b0;
    defparam \tok.i303_4_lut_adj_187_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i303_4_lut_adj_187_LC_6_11_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \tok.i303_4_lut_adj_187_LC_6_11_4  (
            .in0(N__25893),
            .in1(N__19075),
            .in2(N__19102),
            .in3(N__35300),
            .lcout(),
            .ltout(\tok.n252_adj_783_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_189_LC_6_11_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_189_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_189_LC_6_11_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_189_LC_6_11_5  (
            .in0(N__35301),
            .in1(N__19081),
            .in2(N__19099),
            .in3(N__34536),
            .lcout(\tok.n4_adj_786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_184_LC_6_11_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_184_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_184_LC_6_11_6 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \tok.i1_4_lut_adj_184_LC_6_11_6  (
            .in0(N__26316),
            .in1(N__19096),
            .in2(N__19090),
            .in3(N__35724),
            .lcout(\tok.n258_adj_780 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i317_4_lut_adj_183_LC_6_11_7 .C_ON=1'b0;
    defparam \tok.i317_4_lut_adj_183_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i317_4_lut_adj_183_LC_6_11_7 .LUT_INIT=16'b0100010000001010;
    LogicCell40 \tok.i317_4_lut_adj_183_LC_6_11_7  (
            .in0(N__31050),
            .in1(N__22014),
            .in2(N__30312),
            .in3(N__36749),
            .lcout(\tok.n177_adj_779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_56_LC_6_12_0 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_56_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_56_LC_6_12_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \tok.i308_4_lut_adj_56_LC_6_12_0  (
            .in0(N__36978),
            .in1(N__26780),
            .in2(N__26217),
            .in3(N__19363),
            .lcout(\tok.n242_adj_670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_55_LC_6_12_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_55_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_55_LC_6_12_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_55_LC_6_12_1  (
            .in0(N__19354),
            .in1(N__20340),
            .in2(N__24317),
            .in3(N__19334),
            .lcout(),
            .ltout(\tok.n248_adj_669_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_57_LC_6_12_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_57_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_57_LC_6_12_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_57_LC_6_12_2  (
            .in0(N__36979),
            .in1(N__35198),
            .in2(N__19348),
            .in3(N__19345),
            .lcout(),
            .ltout(\tok.n200_adj_671_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_60_LC_6_12_3 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_60_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_60_LC_6_12_3 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i2_4_lut_adj_60_LC_6_12_3  (
            .in0(N__26587),
            .in1(N__33995),
            .in2(N__19339),
            .in3(N__32330),
            .lcout(),
            .ltout(\tok.n6_adj_674_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i15_LC_6_12_4 .C_ON=1'b0;
    defparam \tok.A_i15_LC_6_12_4 .SEQ_MODE=4'b1010;
    defparam \tok.A_i15_LC_6_12_4 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \tok.A_i15_LC_6_12_4  (
            .in0(N__19335),
            .in1(N__25515),
            .in2(N__19270),
            .in3(N__20896),
            .lcout(\tok.n43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38495),
            .ce(N__25644),
            .sr(N__29262));
    defparam \tok.i312_4_lut_adj_244_LC_6_13_0 .C_ON=1'b0;
    defparam \tok.i312_4_lut_adj_244_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.i312_4_lut_adj_244_LC_6_13_0 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \tok.i312_4_lut_adj_244_LC_6_13_0  (
            .in0(N__32965),
            .in1(N__30907),
            .in2(N__19267),
            .in3(N__19389),
            .lcout(),
            .ltout(\tok.n203_adj_822_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_319_LC_6_13_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_319_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_319_LC_6_13_1 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_319_LC_6_13_1  (
            .in0(N__19390),
            .in1(N__19245),
            .in2(N__19168),
            .in3(N__32064),
            .lcout(),
            .ltout(\tok.n212_adj_824_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6928_4_lut_LC_6_13_2 .C_ON=1'b0;
    defparam \tok.i6928_4_lut_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6928_4_lut_LC_6_13_2 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i6928_4_lut_LC_6_13_2  (
            .in0(N__32065),
            .in1(N__33471),
            .in2(N__19165),
            .in3(N__20620),
            .lcout(),
            .ltout(\tok.n6457_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_249_LC_6_13_3 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_249_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_249_LC_6_13_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \tok.i308_4_lut_adj_249_LC_6_13_3  (
            .in0(N__26207),
            .in1(N__36957),
            .in2(N__19162),
            .in3(N__36535),
            .lcout(),
            .ltout(\tok.n242_adj_828_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_250_LC_6_13_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_250_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_250_LC_6_13_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_250_LC_6_13_4  (
            .in0(N__36958),
            .in1(N__19411),
            .in2(N__19399),
            .in3(N__35329),
            .lcout(\tok.n200_adj_829 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_32_LC_6_13_5 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_32_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_32_LC_6_13_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_32_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(N__35264),
            .in2(_gnd_net_),
            .in3(N__36029),
            .lcout(\tok.n4_adj_640 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_100_i9_2_lut_LC_6_13_6 .C_ON=1'b0;
    defparam \tok.or_100_i9_2_lut_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.or_100_i9_2_lut_LC_6_13_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.or_100_i9_2_lut_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__27374),
            .in2(_gnd_net_),
            .in3(N__20793),
            .lcout(\tok.n231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_2_lut_3_lut_LC_6_13_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_2_lut_3_lut_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_2_lut_3_lut_LC_6_13_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \tok.i1_2_lut_2_lut_3_lut_LC_6_13_7  (
            .in0(N__30906),
            .in1(N__36956),
            .in2(_gnd_net_),
            .in3(N__32063),
            .lcout(\tok.n838 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_328_LC_6_14_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_328_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_328_LC_6_14_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_328_LC_6_14_0  (
            .in0(N__35465),
            .in1(N__36955),
            .in2(N__19423),
            .in3(N__19381),
            .lcout(),
            .ltout(\tok.n200_adj_886_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_331_LC_6_14_1 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_331_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_331_LC_6_14_1 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i2_4_lut_adj_331_LC_6_14_1  (
            .in0(N__26610),
            .in1(N__33952),
            .in2(N__19372),
            .in3(N__23953),
            .lcout(),
            .ltout(\tok.n6_adj_889_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i12_LC_6_14_2 .C_ON=1'b0;
    defparam \tok.A_i12_LC_6_14_2 .SEQ_MODE=4'b1010;
    defparam \tok.A_i12_LC_6_14_2 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \tok.A_i12_LC_6_14_2  (
            .in0(N__25516),
            .in1(N__22390),
            .in2(N__19369),
            .in3(N__19522),
            .lcout(\tok.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38502),
            .ce(N__25643),
            .sr(N__29271));
    defparam \tok.i289_2_lut_3_lut_4_lut_LC_6_14_4 .C_ON=1'b0;
    defparam \tok.i289_2_lut_3_lut_4_lut_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \tok.i289_2_lut_3_lut_4_lut_LC_6_14_4 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \tok.i289_2_lut_3_lut_4_lut_LC_6_14_4  (
            .in0(N__36032),
            .in1(N__35265),
            .in2(N__34060),
            .in3(N__36952),
            .lcout(\tok.n8 ),
            .ltout(\tok.n8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6868_2_lut_3_lut_4_lut_LC_6_14_5 .C_ON=1'b0;
    defparam \tok.i6868_2_lut_3_lut_4_lut_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6868_2_lut_3_lut_4_lut_LC_6_14_5 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \tok.i6868_2_lut_3_lut_4_lut_LC_6_14_5  (
            .in0(N__36953),
            .in1(N__30063),
            .in2(N__19366),
            .in3(N__33950),
            .lcout(\tok.n6425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_325_LC_6_14_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_325_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_325_LC_6_14_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_325_LC_6_14_6  (
            .in0(N__20339),
            .in1(N__24329),
            .in2(N__19521),
            .in3(N__19435),
            .lcout(\tok.n248_adj_884 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6875_2_lut_3_lut_4_lut_LC_6_14_7 .C_ON=1'b0;
    defparam \tok.i6875_2_lut_3_lut_4_lut_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6875_2_lut_3_lut_4_lut_LC_6_14_7 .LUT_INIT=16'b0010001000000010;
    LogicCell40 \tok.i6875_2_lut_3_lut_4_lut_LC_6_14_7  (
            .in0(N__36954),
            .in1(N__33951),
            .in2(N__24433),
            .in3(N__23952),
            .lcout(\tok.n6346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i3_LC_7_2_0 .C_ON=1'b0;
    defparam \tok.tc_i3_LC_7_2_0 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i3_LC_7_2_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.tc_i3_LC_7_2_0  (
            .in0(N__19753),
            .in1(N__21264),
            .in2(_gnd_net_),
            .in3(N__22610),
            .lcout(tc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38453),
            .ce(),
            .sr(N__29169));
    defparam \tok.tc_i2_LC_7_2_1 .C_ON=1'b0;
    defparam \tok.tc_i2_LC_7_2_1 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i2_LC_7_2_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.tc_i2_LC_7_2_1  (
            .in0(N__21199),
            .in1(N__19752),
            .in2(_gnd_net_),
            .in3(N__22460),
            .lcout(tc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38453),
            .ce(),
            .sr(N__29169));
    defparam \tok.tc_i1_LC_7_2_2 .C_ON=1'b0;
    defparam \tok.tc_i1_LC_7_2_2 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i1_LC_7_2_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.tc_i1_LC_7_2_2  (
            .in0(N__19751),
            .in1(_gnd_net_),
            .in2(N__22723),
            .in3(N__24959),
            .lcout(tc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38453),
            .ce(),
            .sr(N__29169));
    defparam \tok.tc_i0_LC_7_2_3 .C_ON=1'b0;
    defparam \tok.tc_i0_LC_7_2_3 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i0_LC_7_2_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.tc_i0_LC_7_2_3  (
            .in0(N__19794),
            .in1(N__19750),
            .in2(_gnd_net_),
            .in3(N__21128),
            .lcout(tc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38453),
            .ce(),
            .sr(N__29169));
    defparam \tok.i2534_2_lut_LC_7_2_4 .C_ON=1'b0;
    defparam \tok.i2534_2_lut_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2534_2_lut_LC_7_2_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i2534_2_lut_LC_7_2_4  (
            .in0(N__35500),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33267),
            .lcout(\tok.n2557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_157_LC_7_3_0 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_157_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_157_LC_7_3_0 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_157_LC_7_3_0  (
            .in0(N__21004),
            .in1(N__33268),
            .in2(N__21646),
            .in3(N__31230),
            .lcout(),
            .ltout(\tok.n83_adj_756_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6644_2_lut_3_lut_LC_7_3_1 .C_ON=1'b0;
    defparam \tok.i6644_2_lut_3_lut_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6644_2_lut_3_lut_LC_7_3_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i6644_2_lut_3_lut_LC_7_3_1  (
            .in0(_gnd_net_),
            .in1(N__36316),
            .in2(N__19414),
            .in3(N__31935),
            .lcout(\tok.n6295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6609_4_lut_LC_7_3_2 .C_ON=1'b0;
    defparam \tok.ram.i6609_4_lut_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6609_4_lut_LC_7_3_2 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \tok.ram.i6609_4_lut_LC_7_3_2  (
            .in0(N__21055),
            .in1(N__22932),
            .in2(N__21010),
            .in3(N__22874),
            .lcout(),
            .ltout(\tok.ram.n6260_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1528_4_lut_LC_7_3_3 .C_ON=1'b0;
    defparam \tok.ram.i1528_4_lut_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1528_4_lut_LC_7_3_3 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.ram.i1528_4_lut_LC_7_3_3  (
            .in0(N__21008),
            .in1(N__22790),
            .in2(N__19573),
            .in3(N__31936),
            .lcout(),
            .ltout(\tok.n1565_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_158_LC_7_3_4 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_158_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_158_LC_7_3_4 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i27_4_lut_adj_158_LC_7_3_4  (
            .in0(N__19570),
            .in1(N__35501),
            .in2(N__19564),
            .in3(N__31231),
            .lcout(),
            .ltout(\tok.n13_adj_757_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_159_LC_7_3_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_159_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_159_LC_7_3_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_159_LC_7_3_5  (
            .in0(N__29710),
            .in1(N__25804),
            .in2(N__19561),
            .in3(N__21056),
            .lcout(n10_adj_906),
            .ltout(n10_adj_906_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_205_LC_7_3_6 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_205_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_205_LC_7_3_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \tok.i26_3_lut_adj_205_LC_7_3_6  (
            .in0(_gnd_net_),
            .in1(N__21029),
            .in2(N__19558),
            .in3(N__19748),
            .lcout(\tok.tc_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i4_LC_7_3_7 .C_ON=1'b0;
    defparam \tok.tc_i4_LC_7_3_7 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i4_LC_7_3_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.tc_i4_LC_7_3_7  (
            .in0(N__19749),
            .in1(_gnd_net_),
            .in2(N__21034),
            .in3(N__19537),
            .lcout(tc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38459),
            .ce(),
            .sr(N__29179));
    defparam \tok.i6857_4_lut_LC_7_4_0 .C_ON=1'b0;
    defparam \tok.i6857_4_lut_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6857_4_lut_LC_7_4_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \tok.i6857_4_lut_LC_7_4_0  (
            .in0(N__36251),
            .in1(N__19528),
            .in2(N__37138),
            .in3(N__31319),
            .lcout(\tok.n6622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i303_4_lut_LC_7_4_2 .C_ON=1'b0;
    defparam \tok.i303_4_lut_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i303_4_lut_LC_7_4_2 .LUT_INIT=16'b1000000110001001;
    LogicCell40 \tok.i303_4_lut_LC_7_4_2  (
            .in0(N__36250),
            .in1(N__32096),
            .in2(N__35523),
            .in3(N__31318),
            .lcout(),
            .ltout(\tok.n324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i307_4_lut_LC_7_4_3 .C_ON=1'b0;
    defparam \tok.i307_4_lut_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i307_4_lut_LC_7_4_3 .LUT_INIT=16'b1010101011110011;
    LogicCell40 \tok.i307_4_lut_LC_7_4_3  (
            .in0(N__19642),
            .in1(N__37130),
            .in2(N__19531),
            .in3(N__33265),
            .lcout(\tok.n239_adj_679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_63_LC_7_4_4 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_63_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_63_LC_7_4_4 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \tok.i1_3_lut_adj_63_LC_7_4_4  (
            .in0(N__35496),
            .in1(N__32095),
            .in2(_gnd_net_),
            .in3(N__31316),
            .lcout(\tok.n225_adj_678 ),
            .ltout(\tok.n225_adj_678_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6686_3_lut_4_lut_LC_7_4_5 .C_ON=1'b0;
    defparam \tok.i6686_3_lut_4_lut_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6686_3_lut_4_lut_LC_7_4_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \tok.i6686_3_lut_4_lut_LC_7_4_5  (
            .in0(N__31317),
            .in1(N__37129),
            .in2(N__19645),
            .in3(N__36249),
            .lcout(\tok.n6351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2596_rep_330_2_lut_LC_7_4_6 .C_ON=1'b0;
    defparam \tok.i2596_rep_330_2_lut_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2596_rep_330_2_lut_LC_7_4_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i2596_rep_330_2_lut_LC_7_4_6  (
            .in0(N__34059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32097),
            .lcout(),
            .ltout(\tok.n7456_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i283_4_lut_LC_7_4_7 .C_ON=1'b0;
    defparam \tok.i283_4_lut_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i283_4_lut_LC_7_4_7 .LUT_INIT=16'b1010101000001100;
    LogicCell40 \tok.i283_4_lut_LC_7_4_7  (
            .in0(N__19636),
            .in1(N__25727),
            .in2(N__19630),
            .in3(N__33266),
            .lcout(\tok.n176 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_4_lut_LC_7_5_0 .C_ON=1'b0;
    defparam \tok.i3_3_lut_4_lut_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_4_lut_LC_7_5_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i3_3_lut_4_lut_LC_7_5_0  (
            .in0(N__36232),
            .in1(N__34751),
            .in2(N__37099),
            .in3(N__32043),
            .lcout(\tok.n8_adj_686 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_adj_175_LC_7_5_1 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_adj_175_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_adj_175_LC_7_5_1 .LUT_INIT=16'b1111010011111100;
    LogicCell40 \tok.i1_3_lut_4_lut_adj_175_LC_7_5_1  (
            .in0(N__32045),
            .in1(N__20560),
            .in2(N__34104),
            .in3(N__33270),
            .lcout(\tok.n877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_62_LC_7_5_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_62_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_62_LC_7_5_2 .LUT_INIT=16'b1111111101000101;
    LogicCell40 \tok.i1_4_lut_adj_62_LC_7_5_2  (
            .in0(N__37134),
            .in1(N__19651),
            .in2(N__35505),
            .in3(N__34055),
            .lcout(\tok.n900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_121_LC_7_5_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_121_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_121_LC_7_5_3 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \tok.i1_4_lut_adj_121_LC_7_5_3  (
            .in0(N__34752),
            .in1(N__19600),
            .in2(N__21325),
            .in3(N__33269),
            .lcout(),
            .ltout(\tok.n237_adj_724_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_129_LC_7_5_4 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_129_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_129_LC_7_5_4 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i2_4_lut_adj_129_LC_7_5_4  (
            .in0(N__19579),
            .in1(N__20514),
            .in2(N__19594),
            .in3(N__31235),
            .lcout(\tok.n4893 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_273_LC_7_5_5 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_273_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_273_LC_7_5_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i1_3_lut_adj_273_LC_7_5_5  (
            .in0(N__32044),
            .in1(N__20559),
            .in2(_gnd_net_),
            .in3(N__35423),
            .lcout(\tok.n286 ),
            .ltout(\tok.n286_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i371_4_lut_LC_7_5_6 .C_ON=1'b0;
    defparam \tok.i371_4_lut_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i371_4_lut_LC_7_5_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \tok.i371_4_lut_LC_7_5_6  (
            .in0(N__33271),
            .in1(N__21316),
            .in2(N__19873),
            .in3(N__31236),
            .lcout(),
            .ltout(\tok.n394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_298_LC_7_5_7 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_298_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_298_LC_7_5_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \tok.i1_3_lut_adj_298_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(N__19860),
            .in2(N__19849),
            .in3(N__25120),
            .lcout(\tok.n6143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i7_LC_7_6_0 .C_ON=1'b0;
    defparam \tok.A_i7_LC_7_6_0 .SEQ_MODE=4'b1010;
    defparam \tok.A_i7_LC_7_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_i7_LC_7_6_0  (
            .in0(N__25449),
            .in1(N__25964),
            .in2(_gnd_net_),
            .in3(N__26527),
            .lcout(\tok.A_low_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38474),
            .ce(N__25635),
            .sr(N__29255));
    defparam \tok.i129_3_lut_LC_7_6_1 .C_ON=1'b0;
    defparam \tok.i129_3_lut_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i129_3_lut_LC_7_6_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.i129_3_lut_LC_7_6_1  (
            .in0(N__19716),
            .in1(N__21265),
            .in2(_gnd_net_),
            .in3(N__22620),
            .lcout(\tok.tc_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i129_3_lut_adj_209_LC_7_6_2 .C_ON=1'b0;
    defparam \tok.i129_3_lut_adj_209_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i129_3_lut_adj_209_LC_7_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.i129_3_lut_adj_209_LC_7_6_2  (
            .in0(N__24963),
            .in1(N__22719),
            .in2(_gnd_net_),
            .in3(N__19717),
            .lcout(\tok.tc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i129_3_lut_adj_211_LC_7_6_3 .C_ON=1'b0;
    defparam \tok.i129_3_lut_adj_211_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i129_3_lut_adj_211_LC_7_6_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.i129_3_lut_adj_211_LC_7_6_3  (
            .in0(N__19718),
            .in1(_gnd_net_),
            .in2(N__19795),
            .in3(N__21130),
            .lcout(\tok.tc_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_207_LC_7_6_4 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_207_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_207_LC_7_6_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \tok.i26_3_lut_adj_207_LC_7_6_4  (
            .in0(N__22464),
            .in1(_gnd_net_),
            .in2(N__21198),
            .in3(N__19719),
            .lcout(\tok.tc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_LC_7_6_5 .C_ON=1'b0;
    defparam \tok.i1_3_lut_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_LC_7_6_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \tok.i1_3_lut_LC_7_6_5  (
            .in0(N__25106),
            .in1(N__19942),
            .in2(_gnd_net_),
            .in3(N__36252),
            .lcout(\tok.n6140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6668_3_lut_LC_7_6_6 .C_ON=1'b0;
    defparam \tok.i6668_3_lut_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6668_3_lut_LC_7_6_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \tok.i6668_3_lut_LC_7_6_6  (
            .in0(N__35419),
            .in1(N__34753),
            .in2(_gnd_net_),
            .in3(N__33183),
            .lcout(\tok.n6331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6954_2_lut_3_lut_LC_7_6_7 .C_ON=1'b0;
    defparam \tok.i6954_2_lut_3_lut_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6954_2_lut_3_lut_LC_7_6_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \tok.i6954_2_lut_3_lut_LC_7_6_7  (
            .in0(N__34754),
            .in1(N__32059),
            .in2(_gnd_net_),
            .in3(N__31224),
            .lcout(\tok.n6582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1500_3_lut_LC_7_7_0 .C_ON=1'b0;
    defparam \tok.ram.i1500_3_lut_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1500_3_lut_LC_7_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.ram.i1500_3_lut_LC_7_7_0  (
            .in0(N__28483),
            .in1(N__22347),
            .in2(_gnd_net_),
            .in3(N__21991),
            .lcout(\tok.table_wr_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i127_4_lut_4_lut_LC_7_7_1 .C_ON=1'b0;
    defparam \tok.i127_4_lut_4_lut_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i127_4_lut_4_lut_LC_7_7_1 .LUT_INIT=16'b1001001111001111;
    LogicCell40 \tok.i127_4_lut_4_lut_LC_7_7_1  (
            .in0(N__33167),
            .in1(N__35396),
            .in2(N__31311),
            .in3(N__31979),
            .lcout(\tok.n127_adj_772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i336_4_lut_adj_141_LC_7_7_2 .C_ON=1'b0;
    defparam \tok.i336_4_lut_adj_141_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i336_4_lut_adj_141_LC_7_7_2 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \tok.i336_4_lut_adj_141_LC_7_7_2  (
            .in0(N__23355),
            .in1(N__20017),
            .in2(N__23746),
            .in3(N__31220),
            .lcout(),
            .ltout(\tok.n199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_142_LC_7_7_3 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_142_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_142_LC_7_7_3 .LUT_INIT=16'b1111001100110011;
    LogicCell40 \tok.i1_3_lut_adj_142_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__34612),
            .in2(N__19954),
            .in3(N__31981),
            .lcout(\tok.n262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2588_3_lut_LC_7_7_4 .C_ON=1'b0;
    defparam \tok.i2588_3_lut_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2588_3_lut_LC_7_7_4 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \tok.i2588_3_lut_LC_7_7_4  (
            .in0(N__31980),
            .in1(N__23993),
            .in2(_gnd_net_),
            .in3(N__33168),
            .lcout(\tok.n2611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i291_4_lut_4_lut_4_lut_LC_7_7_5 .C_ON=1'b0;
    defparam \tok.i291_4_lut_4_lut_4_lut_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i291_4_lut_4_lut_4_lut_LC_7_7_5 .LUT_INIT=16'b0000011100100010;
    LogicCell40 \tok.i291_4_lut_4_lut_4_lut_LC_7_7_5  (
            .in0(N__36215),
            .in1(N__34611),
            .in2(N__32112),
            .in3(N__35397),
            .lcout(\tok.n311_adj_721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_38_LC_7_7_6 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_38_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_38_LC_7_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i1_2_lut_adj_38_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__31216),
            .in2(_gnd_net_),
            .in3(N__33166),
            .lcout(\tok.n4_adj_648 ),
            .ltout(\tok.n4_adj_648_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i305_4_lut_4_lut_LC_7_7_7 .C_ON=1'b0;
    defparam \tok.i305_4_lut_4_lut_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i305_4_lut_4_lut_LC_7_7_7 .LUT_INIT=16'b0111000011001100;
    LogicCell40 \tok.i305_4_lut_4_lut_LC_7_7_7  (
            .in0(N__36214),
            .in1(N__34610),
            .in2(N__19945),
            .in3(N__31978),
            .lcout(\tok.n326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i304_4_lut_4_lut_adj_333_LC_7_8_0 .C_ON=1'b0;
    defparam \tok.i304_4_lut_4_lut_adj_333_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i304_4_lut_4_lut_adj_333_LC_7_8_0 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \tok.i304_4_lut_4_lut_adj_333_LC_7_8_0  (
            .in0(N__31239),
            .in1(N__19936),
            .in2(N__19905),
            .in3(N__31905),
            .lcout(\tok.n210_adj_784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_4_lut_adj_332_LC_7_8_1 .C_ON=1'b0;
    defparam \tok.i2_4_lut_4_lut_adj_332_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_4_lut_adj_332_LC_7_8_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \tok.i2_4_lut_4_lut_adj_332_LC_7_8_1  (
            .in0(N__31906),
            .in1(N__31240),
            .in2(N__23113),
            .in3(N__37112),
            .lcout(),
            .ltout(\tok.n4842_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_122_LC_7_8_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_122_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_122_LC_7_8_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \tok.i1_4_lut_adj_122_LC_7_8_2  (
            .in0(N__20437),
            .in1(N__20026),
            .in2(N__20110),
            .in3(N__22943),
            .lcout(\tok.n239_adj_727 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_rep_325_2_lut_LC_7_8_3 .C_ON=1'b0;
    defparam \tok.i1_rep_325_2_lut_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_rep_325_2_lut_LC_7_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i1_rep_325_2_lut_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__37111),
            .in2(_gnd_net_),
            .in3(N__31237),
            .lcout(),
            .ltout(\tok.n7451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6956_4_lut_LC_7_8_4 .C_ON=1'b0;
    defparam \tok.i6956_4_lut_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6956_4_lut_LC_7_8_4 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \tok.i6956_4_lut_LC_7_8_4  (
            .in0(N__34722),
            .in1(N__20088),
            .in2(N__20107),
            .in3(N__20104),
            .lcout(\tok.n6624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i297_4_lut_LC_7_8_5 .C_ON=1'b0;
    defparam \tok.i297_4_lut_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i297_4_lut_LC_7_8_5 .LUT_INIT=16'b0010000000101100;
    LogicCell40 \tok.i297_4_lut_LC_7_8_5  (
            .in0(N__20089),
            .in1(N__31238),
            .in2(N__37135),
            .in3(N__33581),
            .lcout(\tok.n164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6833_4_lut_LC_7_8_6 .C_ON=1'b0;
    defparam \tok.i6833_4_lut_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6833_4_lut_LC_7_8_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \tok.i6833_4_lut_LC_7_8_6  (
            .in0(N__34723),
            .in1(N__23216),
            .in2(N__35503),
            .in3(N__33031),
            .lcout(\tok.n6597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i335_4_lut_LC_7_8_7 .C_ON=1'b0;
    defparam \tok.i335_4_lut_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i335_4_lut_LC_7_8_7 .LUT_INIT=16'b0011001100001010;
    LogicCell40 \tok.i335_4_lut_LC_7_8_7  (
            .in0(N__20011),
            .in1(N__20488),
            .in2(N__19999),
            .in3(N__35415),
            .lcout(\tok.n247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_LC_7_9_1 .C_ON=1'b0;
    defparam \tok.i308_4_lut_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_LC_7_9_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \tok.i308_4_lut_LC_7_9_1  (
            .in0(N__37124),
            .in1(N__37386),
            .in2(N__26221),
            .in3(N__19987),
            .lcout(),
            .ltout(\tok.n242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_27_LC_7_9_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_27_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_27_LC_7_9_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_27_LC_7_9_2  (
            .in0(N__35377),
            .in1(N__37125),
            .in2(N__19978),
            .in3(N__20278),
            .lcout(\tok.n200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_26_LC_7_9_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_26_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_26_LC_7_9_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_26_LC_7_9_3  (
            .in0(N__20284),
            .in1(N__20321),
            .in2(N__24337),
            .in3(N__20259),
            .lcout(\tok.n248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6630_4_lut_LC_7_9_4 .C_ON=1'b0;
    defparam \tok.i6630_4_lut_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6630_4_lut_LC_7_9_4 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \tok.i6630_4_lut_LC_7_9_4  (
            .in0(N__37387),
            .in1(N__34129),
            .in2(N__26615),
            .in3(N__21796),
            .lcout(),
            .ltout(\tok.n6606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i8_LC_7_9_5 .C_ON=1'b0;
    defparam \tok.A_i8_LC_7_9_5 .SEQ_MODE=4'b1010;
    defparam \tok.A_i8_LC_7_9_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_i8_LC_7_9_5  (
            .in0(N__25467),
            .in1(_gnd_net_),
            .in2(N__20272),
            .in3(N__28329),
            .lcout(A_low_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38486),
            .ce(N__25651),
            .sr(N__29241));
    defparam \tok.i2_4_lut_LC_7_9_6 .C_ON=1'b0;
    defparam \tok.i2_4_lut_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_LC_7_9_6 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \tok.i2_4_lut_LC_7_9_6  (
            .in0(N__34005),
            .in1(N__27011),
            .in2(N__26616),
            .in3(N__20269),
            .lcout(),
            .ltout(\tok.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i13_LC_7_9_7 .C_ON=1'b0;
    defparam \tok.A_i13_LC_7_9_7 .SEQ_MODE=4'b1010;
    defparam \tok.A_i13_LC_7_9_7 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \tok.A_i13_LC_7_9_7  (
            .in0(N__25466),
            .in1(N__21688),
            .in2(N__20263),
            .in3(N__20260),
            .lcout(\tok.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38486),
            .ce(N__25651),
            .sr(N__29241));
    defparam \tok.i6591_2_lut_LC_7_10_0 .C_ON=1'b0;
    defparam \tok.i6591_2_lut_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6591_2_lut_LC_7_10_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i6591_2_lut_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__34030),
            .in2(_gnd_net_),
            .in3(N__29547),
            .lcout(\tok.n6344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_314_LC_7_10_1 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_314_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_314_LC_7_10_1 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \tok.i2_4_lut_adj_314_LC_7_10_1  (
            .in0(N__29549),
            .in1(N__26586),
            .in2(N__34100),
            .in3(N__20203),
            .lcout(),
            .ltout(\tok.n6_adj_878_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i11_LC_7_10_2 .C_ON=1'b0;
    defparam \tok.A_i11_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \tok.A_i11_LC_7_10_2 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \tok.A_i11_LC_7_10_2  (
            .in0(N__25479),
            .in1(N__20926),
            .in2(N__20194),
            .in3(N__20191),
            .lcout(\tok.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38490),
            .ce(N__25649),
            .sr(N__29270));
    defparam \tok.i2577_2_lut_LC_7_10_3 .C_ON=1'b0;
    defparam \tok.i2577_2_lut_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2577_2_lut_LC_7_10_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i2577_2_lut_LC_7_10_3  (
            .in0(N__34031),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30258),
            .lcout(),
            .ltout(\tok.n2600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i310_4_lut_adj_311_LC_7_10_4 .C_ON=1'b0;
    defparam \tok.i310_4_lut_adj_311_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i310_4_lut_adj_311_LC_7_10_4 .LUT_INIT=16'b0001101100001010;
    LogicCell40 \tok.i310_4_lut_adj_311_LC_7_10_4  (
            .in0(N__31072),
            .in1(N__33417),
            .in2(N__20473),
            .in3(N__29548),
            .lcout(\tok.n215_adj_876 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6777_4_lut_LC_7_10_5 .C_ON=1'b0;
    defparam \tok.i6777_4_lut_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6777_4_lut_LC_7_10_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \tok.i6777_4_lut_LC_7_10_5  (
            .in0(N__26583),
            .in1(N__30259),
            .in2(N__30547),
            .in3(N__20446),
            .lcout(),
            .ltout(\tok.n6610_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i6_LC_7_10_6 .C_ON=1'b0;
    defparam \tok.A_i6_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \tok.A_i6_LC_7_10_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_i6_LC_7_10_6  (
            .in0(N__25480),
            .in1(_gnd_net_),
            .in2(N__20470),
            .in3(N__22029),
            .lcout(\tok.A_low_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38490),
            .ce(N__25649),
            .sr(N__29270));
    defparam \tok.i310_4_lut_adj_82_LC_7_10_7 .C_ON=1'b0;
    defparam \tok.i310_4_lut_adj_82_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i310_4_lut_adj_82_LC_7_10_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.i310_4_lut_adj_82_LC_7_10_7  (
            .in0(N__33416),
            .in1(N__24179),
            .in2(N__20467),
            .in3(N__31071),
            .lcout(\tok.n215_adj_697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_LC_7_11_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_LC_7_11_0 .LUT_INIT=16'b0110001000000000;
    LogicCell40 \tok.i1_4_lut_4_lut_LC_7_11_0  (
            .in0(N__32956),
            .in1(N__35279),
            .in2(N__36138),
            .in3(N__34843),
            .lcout(),
            .ltout(\tok.n269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_110_LC_7_11_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_110_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_110_LC_7_11_1 .LUT_INIT=16'b1111100011111101;
    LogicCell40 \tok.i1_4_lut_adj_110_LC_7_11_1  (
            .in0(N__31069),
            .in1(N__26013),
            .in2(N__20458),
            .in3(N__20575),
            .lcout(\tok.n229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_193_LC_7_11_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_193_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_193_LC_7_11_2 .LUT_INIT=16'b0011000100110000;
    LogicCell40 \tok.i1_4_lut_adj_193_LC_7_11_2  (
            .in0(N__32957),
            .in1(N__33986),
            .in2(N__20455),
            .in3(N__21922),
            .lcout(\tok.n205_adj_789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6683_3_lut_4_lut_LC_7_11_3 .C_ON=1'b0;
    defparam \tok.i6683_3_lut_4_lut_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6683_3_lut_4_lut_LC_7_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \tok.i6683_3_lut_4_lut_LC_7_11_3  (
            .in0(N__35278),
            .in1(N__35918),
            .in2(N__20425),
            .in3(N__32955),
            .lcout(),
            .ltout(\tok.n6341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i311_4_lut_LC_7_11_4 .C_ON=1'b0;
    defparam \tok.i311_4_lut_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i311_4_lut_LC_7_11_4 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \tok.i311_4_lut_LC_7_11_4  (
            .in0(N__20573),
            .in1(N__27122),
            .in2(N__20347),
            .in3(N__31068),
            .lcout(\tok.n170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i5_1_lut_LC_7_11_5 .C_ON=1'b0;
    defparam \tok.inv_105_i5_1_lut_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i5_1_lut_LC_7_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i5_1_lut_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27262),
            .lcout(\tok.n321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_64_LC_7_11_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_64_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_64_LC_7_11_6 .LUT_INIT=16'b0000000011110100;
    LogicCell40 \tok.i1_4_lut_adj_64_LC_7_11_6  (
            .in0(N__20574),
            .in1(N__31956),
            .in2(N__20558),
            .in3(N__31070),
            .lcout(),
            .ltout(\tok.n238_adj_681_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_65_LC_7_11_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_65_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_65_LC_7_11_7 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \tok.i1_4_lut_adj_65_LC_7_11_7  (
            .in0(N__34844),
            .in1(N__20530),
            .in2(N__20518),
            .in3(N__20515),
            .lcout(\tok.n194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6870_2_lut_3_lut_4_lut_LC_7_12_0 .C_ON=1'b0;
    defparam \tok.i6870_2_lut_3_lut_4_lut_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6870_2_lut_3_lut_4_lut_LC_7_12_0 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \tok.i6870_2_lut_3_lut_4_lut_LC_7_12_0  (
            .in0(N__22191),
            .in1(N__33872),
            .in2(N__24463),
            .in3(N__37046),
            .lcout(\tok.n6396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i9_1_lut_LC_7_12_1 .C_ON=1'b0;
    defparam \tok.inv_105_i9_1_lut_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i9_1_lut_LC_7_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i9_1_lut_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22190),
            .lcout(\tok.n317_adj_659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2639_3_lut_LC_7_12_3 .C_ON=1'b0;
    defparam \tok.i2639_3_lut_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2639_3_lut_LC_7_12_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i2639_3_lut_LC_7_12_3  (
            .in0(N__37045),
            .in1(N__26831),
            .in2(_gnd_net_),
            .in3(N__34514),
            .lcout(\tok.n2663 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6100_2_lut_3_lut_LC_7_12_4 .C_ON=1'b0;
    defparam \tok.i6100_2_lut_3_lut_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6100_2_lut_3_lut_LC_7_12_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i6100_2_lut_3_lut_LC_7_12_4  (
            .in0(N__25376),
            .in1(N__33871),
            .in2(_gnd_net_),
            .in3(N__35127),
            .lcout(\tok.n6183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i6_LC_7_12_5 .C_ON=1'b0;
    defparam \tok.uart.sender_i6_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i6_LC_7_12_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i6_LC_7_12_5  (
            .in0(N__27205),
            .in1(N__37565),
            .in2(_gnd_net_),
            .in3(N__36555),
            .lcout(\tok.uart.sender_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38500),
            .ce(N__27170),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i5_LC_7_12_6 .C_ON=1'b0;
    defparam \tok.uart.sender_i5_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i5_LC_7_12_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \tok.uart.sender_i5_LC_7_12_6  (
            .in0(N__33632),
            .in1(_gnd_net_),
            .in2(N__37567),
            .in3(N__20479),
            .lcout(\tok.uart.sender_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38500),
            .ce(N__27170),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i4_LC_7_12_7 .C_ON=1'b0;
    defparam \tok.uart.sender_i4_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i4_LC_7_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i4_LC_7_12_7  (
            .in0(N__20869),
            .in1(N__37561),
            .in2(_gnd_net_),
            .in3(N__27544),
            .lcout(\tok.uart.sender_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38500),
            .ce(N__27170),
            .sr(_gnd_net_));
    defparam \tok.i6935_3_lut_4_lut_LC_7_13_0 .C_ON=1'b0;
    defparam \tok.i6935_3_lut_4_lut_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6935_3_lut_4_lut_LC_7_13_0 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \tok.i6935_3_lut_4_lut_LC_7_13_0  (
            .in0(N__27378),
            .in1(N__34054),
            .in2(N__24437),
            .in3(N__36148),
            .lcout(\tok.n6450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i310_4_lut_adj_251_LC_7_13_1 .C_ON=1'b0;
    defparam \tok.i310_4_lut_adj_251_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i310_4_lut_adj_251_LC_7_13_1 .LUT_INIT=16'b0000111100100010;
    LogicCell40 \tok.i310_4_lut_adj_251_LC_7_13_1  (
            .in0(N__22245),
            .in1(N__33479),
            .in2(N__20851),
            .in3(N__31090),
            .lcout(),
            .ltout(\tok.n215_adj_830_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6792_4_lut_LC_7_13_2 .C_ON=1'b0;
    defparam \tok.i6792_4_lut_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6792_4_lut_LC_7_13_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.i6792_4_lut_LC_7_13_2  (
            .in0(N__26938),
            .in1(N__20836),
            .in2(N__20830),
            .in3(N__35389),
            .lcout(),
            .ltout(\tok.n6605_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7003_4_lut_LC_7_13_3 .C_ON=1'b0;
    defparam \tok.i7003_4_lut_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.i7003_4_lut_LC_7_13_3 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \tok.i7003_4_lut_LC_7_13_3  (
            .in0(N__34483),
            .in1(N__35390),
            .in2(N__20827),
            .in3(N__20800),
            .lcout(\tok.n6604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i309_4_lut_adj_253_LC_7_13_4 .C_ON=1'b0;
    defparam \tok.i309_4_lut_adj_253_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i309_4_lut_adj_253_LC_7_13_4 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \tok.i309_4_lut_adj_253_LC_7_13_4  (
            .in0(N__20812),
            .in1(N__22244),
            .in2(N__24551),
            .in3(N__36149),
            .lcout(\tok.n179_adj_831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6747_3_lut_4_lut_LC_7_13_5 .C_ON=1'b0;
    defparam \tok.i6747_3_lut_4_lut_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6747_3_lut_4_lut_LC_7_13_5 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \tok.i6747_3_lut_4_lut_LC_7_13_5  (
            .in0(N__34482),
            .in1(N__31089),
            .in2(N__27392),
            .in3(N__20794),
            .lcout(),
            .ltout(\tok.n6462_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i300_4_lut_adj_245_LC_7_13_6 .C_ON=1'b0;
    defparam \tok.i300_4_lut_adj_245_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.i300_4_lut_adj_245_LC_7_13_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \tok.i300_4_lut_adj_245_LC_7_13_6  (
            .in0(N__36281),
            .in1(N__22243),
            .in2(N__20698),
            .in3(N__20691),
            .lcout(\tok.n206_adj_823 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i12_1_lut_LC_7_13_7 .C_ON=1'b0;
    defparam \tok.inv_105_i12_1_lut_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i12_1_lut_LC_7_13_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \tok.inv_105_i12_1_lut_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__23968),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i309_4_lut_adj_313_LC_7_14_0 .C_ON=1'b0;
    defparam \tok.i309_4_lut_adj_313_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \tok.i309_4_lut_adj_313_LC_7_14_0 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \tok.i309_4_lut_adj_313_LC_7_14_0  (
            .in0(N__36150),
            .in1(N__20956),
            .in2(N__29596),
            .in3(N__24540),
            .lcout(\tok.n179_adj_877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i309_4_lut_adj_83_LC_7_14_1 .C_ON=1'b0;
    defparam \tok.i309_4_lut_adj_83_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \tok.i309_4_lut_adj_83_LC_7_14_1 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \tok.i309_4_lut_adj_83_LC_7_14_1  (
            .in0(N__24541),
            .in1(N__36152),
            .in2(N__24180),
            .in3(N__20950),
            .lcout(\tok.n179_adj_698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6844_4_lut_LC_7_14_2 .C_ON=1'b0;
    defparam \tok.i6844_4_lut_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6844_4_lut_LC_7_14_2 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \tok.i6844_4_lut_LC_7_14_2  (
            .in0(N__35384),
            .in1(N__26931),
            .in2(N__22381),
            .in3(N__20944),
            .lcout(),
            .ltout(\tok.n6553_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6995_4_lut_LC_7_14_3 .C_ON=1'b0;
    defparam \tok.i6995_4_lut_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6995_4_lut_LC_7_14_3 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \tok.i6995_4_lut_LC_7_14_3  (
            .in0(N__34792),
            .in1(N__20935),
            .in2(N__20929),
            .in3(N__35386),
            .lcout(\tok.n6552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6948_4_lut_LC_7_14_4 .C_ON=1'b0;
    defparam \tok.i6948_4_lut_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6948_4_lut_LC_7_14_4 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \tok.i6948_4_lut_LC_7_14_4  (
            .in0(N__35388),
            .in1(N__20914),
            .in2(N__22357),
            .in3(N__34794),
            .lcout(\tok.n6537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6772_4_lut_LC_7_14_5 .C_ON=1'b0;
    defparam \tok.i6772_4_lut_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6772_4_lut_LC_7_14_5 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \tok.i6772_4_lut_LC_7_14_5  (
            .in0(N__24073),
            .in1(N__21892),
            .in2(N__26937),
            .in3(N__35385),
            .lcout(),
            .ltout(\tok.n6541_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6847_4_lut_LC_7_14_6 .C_ON=1'b0;
    defparam \tok.i6847_4_lut_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6847_4_lut_LC_7_14_6 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \tok.i6847_4_lut_LC_7_14_6  (
            .in0(N__35387),
            .in1(N__20875),
            .in2(N__20899),
            .in3(N__34793),
            .lcout(\tok.n6540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i309_4_lut_adj_59_LC_7_14_7 .C_ON=1'b0;
    defparam \tok.i309_4_lut_adj_59_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \tok.i309_4_lut_adj_59_LC_7_14_7 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i309_4_lut_adj_59_LC_7_14_7  (
            .in0(N__20884),
            .in1(N__36151),
            .in2(N__24554),
            .in3(N__32354),
            .lcout(\tok.n179_adj_673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i0_LC_8_1_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i0_LC_8_1_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i0_LC_8_1_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.C_stk.tail_i0_i0_LC_8_1_0  (
            .in0(N__24696),
            .in1(N__28733),
            .in2(_gnd_net_),
            .in3(N__21089),
            .lcout(\tok.C_stk.tail_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38454),
            .ce(N__28909),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i6146_3_lut_LC_8_1_1 .C_ON=1'b0;
    defparam \tok.C_stk.i6146_3_lut_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i6146_3_lut_LC_8_1_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i6146_3_lut_LC_8_1_1  (
            .in0(N__21069),
            .in1(N__28116),
            .in2(_gnd_net_),
            .in3(N__21171),
            .lcout(),
            .ltout(\tok.C_stk.n6230_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i0_LC_8_1_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i0_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i0_LC_8_1_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i0_LC_8_1_2  (
            .in0(N__28054),
            .in1(N__27929),
            .in2(N__21133),
            .in3(N__21129),
            .lcout(c_stk_r_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38454),
            .ce(N__28909),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i8_LC_8_1_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i8_LC_8_1_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i8_LC_8_1_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.C_stk.tail_i0_i8_LC_8_1_3  (
            .in0(N__28734),
            .in1(_gnd_net_),
            .in2(N__21073),
            .in3(N__24670),
            .lcout(tail_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38454),
            .ce(N__28909),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i4_LC_8_2_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i4_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i4_LC_8_2_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i4_LC_8_2_0  (
            .in0(N__28747),
            .in1(N__20977),
            .in2(_gnd_net_),
            .in3(N__21009),
            .lcout(\tok.C_stk.tail_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38460),
            .ce(N__28918),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i6155_3_lut_LC_8_2_1 .C_ON=1'b0;
    defparam \tok.C_stk.i6155_3_lut_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i6155_3_lut_LC_8_2_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i6155_3_lut_LC_8_2_1  (
            .in0(N__20985),
            .in1(N__28098),
            .in2(_gnd_net_),
            .in3(N__21061),
            .lcout(),
            .ltout(\tok.C_stk.n6239_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i4_LC_8_2_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i4_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i4_LC_8_2_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i4_LC_8_2_2  (
            .in0(N__27924),
            .in1(N__28047),
            .in2(N__21037),
            .in3(N__21033),
            .lcout(\tok.c_stk_r_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38460),
            .ce(N__28918),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i12_LC_8_2_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i12_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i12_LC_8_2_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i12_LC_8_2_3  (
            .in0(N__20986),
            .in1(_gnd_net_),
            .in2(N__20968),
            .in3(N__28742),
            .lcout(\tok.tail_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38460),
            .ce(N__28918),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i20_LC_8_2_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i20_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i20_LC_8_2_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i20_LC_8_2_4  (
            .in0(N__28743),
            .in1(N__21220),
            .in2(_gnd_net_),
            .in3(N__20976),
            .lcout(\tok.C_stk.tail_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38460),
            .ce(N__28918),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i28_LC_8_2_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i28_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i28_LC_8_2_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i28_LC_8_2_5  (
            .in0(N__20964),
            .in1(N__21211),
            .in2(_gnd_net_),
            .in3(N__28744),
            .lcout(\tok.tail_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38460),
            .ce(N__28918),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i36_LC_8_2_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i36_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i36_LC_8_2_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i36_LC_8_2_6  (
            .in0(N__28745),
            .in1(N__24870),
            .in2(_gnd_net_),
            .in3(N__21219),
            .lcout(\tok.C_stk.tail_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38460),
            .ce(N__28918),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i44_LC_8_2_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i44_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i44_LC_8_2_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i44_LC_8_2_7  (
            .in0(N__24751),
            .in1(N__21210),
            .in2(_gnd_net_),
            .in3(N__28746),
            .lcout(\tok.tail_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38460),
            .ce(N__28918),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_140_LC_8_3_0 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_140_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_140_LC_8_3_0 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \tok.i125_4_lut_adj_140_LC_8_3_0  (
            .in0(N__21562),
            .in1(N__33274),
            .in2(N__22435),
            .in3(N__31297),
            .lcout(),
            .ltout(\tok.n83_adj_723_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6979_2_lut_3_lut_LC_8_3_1 .C_ON=1'b0;
    defparam \tok.i6979_2_lut_3_lut_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6979_2_lut_3_lut_LC_8_3_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \tok.i6979_2_lut_3_lut_LC_8_3_1  (
            .in0(N__36315),
            .in1(_gnd_net_),
            .in2(N__21202),
            .in3(N__31879),
            .lcout(\tok.n6664 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_148_LC_8_3_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_148_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_148_LC_8_3_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_148_LC_8_3_2  (
            .in0(N__21292),
            .in1(N__29706),
            .in2(N__22501),
            .in3(N__25808),
            .lcout(n10_adj_908),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_181_LC_8_3_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_181_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_181_LC_8_3_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \tok.i1_2_lut_adj_181_LC_8_3_3  (
            .in0(N__33273),
            .in1(_gnd_net_),
            .in2(N__36325),
            .in3(_gnd_net_),
            .lcout(\tok.n2573 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_194_LC_8_3_4 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_194_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_194_LC_8_3_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i1_2_lut_adj_194_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__36311),
            .in2(_gnd_net_),
            .in3(N__33272),
            .lcout(\tok.n4_adj_726 ),
            .ltout(\tok.n4_adj_726_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i6600_4_lut_LC_8_3_5 .C_ON=1'b0;
    defparam \tok.ram.i6600_4_lut_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i6600_4_lut_LC_8_3_5 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \tok.ram.i6600_4_lut_LC_8_3_5  (
            .in0(N__22432),
            .in1(N__22497),
            .in2(N__21178),
            .in3(N__22870),
            .lcout(),
            .ltout(\tok.ram.n6257_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1564_4_lut_LC_8_3_6 .C_ON=1'b0;
    defparam \tok.ram.i1564_4_lut_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1564_4_lut_LC_8_3_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \tok.ram.i1564_4_lut_LC_8_3_6  (
            .in0(N__31880),
            .in1(N__22775),
            .in2(N__21175),
            .in3(N__22433),
            .lcout(),
            .ltout(\tok.n1600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_LC_8_3_7 .C_ON=1'b0;
    defparam \tok.i27_4_lut_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_LC_8_3_7 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \tok.i27_4_lut_LC_8_3_7  (
            .in0(N__31298),
            .in1(N__21301),
            .in2(N__21295),
            .in3(N__35331),
            .lcout(\tok.n13_adj_742 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6675_4_lut_LC_8_4_0 .C_ON=1'b0;
    defparam \tok.i6675_4_lut_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6675_4_lut_LC_8_4_0 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \tok.i6675_4_lut_LC_8_4_0  (
            .in0(N__22914),
            .in1(N__22583),
            .in2(N__22660),
            .in3(N__22868),
            .lcout(),
            .ltout(\tok.n6301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i124_4_lut_adj_152_LC_8_4_1 .C_ON=1'b0;
    defparam \tok.i124_4_lut_adj_152_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.i124_4_lut_adj_152_LC_8_4_1 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \tok.i124_4_lut_adj_152_LC_8_4_1  (
            .in0(N__22584),
            .in1(N__32122),
            .in2(N__21286),
            .in3(N__22791),
            .lcout(),
            .ltout(\tok.n80_adj_751_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i126_4_lut_adj_155_LC_8_4_2 .C_ON=1'b0;
    defparam \tok.i126_4_lut_adj_155_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i126_4_lut_adj_155_LC_8_4_2 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \tok.i126_4_lut_adj_155_LC_8_4_2  (
            .in0(N__31323),
            .in1(N__21277),
            .in2(N__21283),
            .in3(N__35330),
            .lcout(\tok.n89_adj_754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_149_LC_8_4_3 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_149_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_149_LC_8_4_3 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_149_LC_8_4_3  (
            .in0(N__22582),
            .in1(N__33275),
            .in2(N__21244),
            .in3(N__31320),
            .lcout(),
            .ltout(\tok.n83_adj_746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6647_2_lut_3_lut_LC_8_4_4 .C_ON=1'b0;
    defparam \tok.i6647_2_lut_3_lut_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6647_2_lut_3_lut_LC_8_4_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i6647_2_lut_3_lut_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(N__36253),
            .in2(N__21280),
            .in3(N__32121),
            .lcout(\tok.n6297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_156_LC_8_4_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_156_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_156_LC_8_4_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_156_LC_8_4_5  (
            .in0(N__21271),
            .in1(N__25807),
            .in2(N__29724),
            .in3(N__22659),
            .lcout(n92_adj_898),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i335_4_lut_adj_135_LC_8_4_6 .C_ON=1'b0;
    defparam \tok.i335_4_lut_adj_135_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i335_4_lut_adj_135_LC_8_4_6 .LUT_INIT=16'b1111111001010100;
    LogicCell40 \tok.i335_4_lut_adj_135_LC_8_4_6  (
            .in0(N__31321),
            .in1(N__21243),
            .in2(N__33300),
            .in3(N__21487),
            .lcout(\tok.n2700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_3_lut_LC_8_4_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_3_lut_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_3_lut_LC_8_4_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \tok.i1_4_lut_3_lut_LC_8_4_7  (
            .in0(N__21486),
            .in1(N__33279),
            .in2(_gnd_net_),
            .in3(N__31322),
            .lcout(\tok.n236_adj_737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_4_lut_LC_8_5_0 .C_ON=1'b0;
    defparam \tok.i2_2_lut_4_lut_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_4_lut_LC_8_5_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \tok.i2_2_lut_4_lut_LC_8_5_0  (
            .in0(N__35490),
            .in1(N__37091),
            .in2(N__34113),
            .in3(N__36233),
            .lcout(\tok.n14_adj_683 ),
            .ltout(\tok.n14_adj_683_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_adj_67_LC_8_5_1 .C_ON=1'b0;
    defparam \tok.i2_2_lut_adj_67_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_adj_67_LC_8_5_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \tok.i2_2_lut_adj_67_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21370),
            .in3(N__21381),
            .lcout(\tok.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.stall_I_0_400_i15_2_lut_LC_8_5_2 .C_ON=1'b0;
    defparam \tok.stall_I_0_400_i15_2_lut_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.stall_I_0_400_i15_2_lut_LC_8_5_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \tok.stall_I_0_400_i15_2_lut_LC_8_5_2  (
            .in0(N__35492),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37093),
            .lcout(),
            .ltout(\tok.n15_adj_807_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_222_LC_8_5_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_222_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_222_LC_8_5_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i1_4_lut_adj_222_LC_8_5_3  (
            .in0(N__23119),
            .in1(N__21367),
            .in2(N__21352),
            .in3(N__33485),
            .lcout(\tok.n903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i406_4_lut_LC_8_5_4 .C_ON=1'b0;
    defparam \tok.C_stk.i406_4_lut_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i406_4_lut_LC_8_5_4 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \tok.C_stk.i406_4_lut_LC_8_5_4  (
            .in0(N__21382),
            .in1(N__23002),
            .in2(N__21337),
            .in3(N__28004),
            .lcout(\tok.C_stk.n449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_111_LC_8_5_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_111_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_111_LC_8_5_5 .LUT_INIT=16'b0000000000111011;
    LogicCell40 \tok.i1_4_lut_adj_111_LC_8_5_5  (
            .in0(N__36235),
            .in1(N__35493),
            .in2(N__26131),
            .in3(N__37097),
            .lcout(\tok.n278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6855_4_lut_4_lut_LC_8_5_6 .C_ON=1'b0;
    defparam \tok.i6855_4_lut_4_lut_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6855_4_lut_4_lut_LC_8_5_6 .LUT_INIT=16'b1000000111111111;
    LogicCell40 \tok.i6855_4_lut_4_lut_LC_8_5_6  (
            .in0(N__35491),
            .in1(N__36234),
            .in2(N__32126),
            .in3(N__37092),
            .lcout(\tok.n6621 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i362_4_lut_4_lut_LC_8_5_7 .C_ON=1'b0;
    defparam \tok.i362_4_lut_4_lut_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i362_4_lut_4_lut_LC_8_5_7 .LUT_INIT=16'b1100000000100010;
    LogicCell40 \tok.i362_4_lut_4_lut_LC_8_5_7  (
            .in0(N__32106),
            .in1(N__34790),
            .in2(N__36310),
            .in3(N__37098),
            .lcout(\tok.n241_adj_747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6829_4_lut_LC_8_6_0 .C_ON=1'b0;
    defparam \tok.i6829_4_lut_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6829_4_lut_LC_8_6_0 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \tok.i6829_4_lut_LC_8_6_0  (
            .in0(N__31877),
            .in1(N__22039),
            .in2(N__34759),
            .in3(N__21451),
            .lcout(\tok.n6593 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_137_LC_8_6_1 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_137_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_137_LC_8_6_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i2_3_lut_adj_137_LC_8_6_1  (
            .in0(N__31161),
            .in1(N__21480),
            .in2(_gnd_net_),
            .in3(N__36254),
            .lcout(\tok.n4925 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6726_2_lut_LC_8_6_2 .C_ON=1'b0;
    defparam \tok.i6726_2_lut_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6726_2_lut_LC_8_6_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i6726_2_lut_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__21445),
            .in2(_gnd_net_),
            .in3(N__33165),
            .lcout(),
            .ltout(\tok.n6578_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6840_4_lut_LC_8_6_3 .C_ON=1'b0;
    defparam \tok.i6840_4_lut_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6840_4_lut_LC_8_6_3 .LUT_INIT=16'b0010001010100000;
    LogicCell40 \tok.i6840_4_lut_LC_8_6_3  (
            .in0(N__21406),
            .in1(N__21433),
            .in2(N__21418),
            .in3(N__31876),
            .lcout(\tok.n6581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_219_LC_8_6_4 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_219_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_219_LC_8_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i1_2_lut_adj_219_LC_8_6_4  (
            .in0(N__34606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31160),
            .lcout(\tok.n4_adj_739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6953_4_lut_LC_8_6_5 .C_ON=1'b0;
    defparam \tok.i6953_4_lut_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6953_4_lut_LC_8_6_5 .LUT_INIT=16'b1111111110110001;
    LogicCell40 \tok.i6953_4_lut_LC_8_6_5  (
            .in0(N__31163),
            .in1(N__21400),
            .in2(N__23143),
            .in3(N__36255),
            .lcout(\tok.n6580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_4_lut_LC_8_6_6 .C_ON=1'b0;
    defparam \tok.i1_2_lut_4_lut_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_4_lut_LC_8_6_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \tok.i1_2_lut_4_lut_LC_8_6_6  (
            .in0(N__31875),
            .in1(N__33164),
            .in2(N__34758),
            .in3(N__31159),
            .lcout(\tok.n4_adj_684 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_228_LC_8_6_7 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_228_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_228_LC_8_6_7 .LUT_INIT=16'b0001000000100000;
    LogicCell40 \tok.i5_4_lut_adj_228_LC_8_6_7  (
            .in0(N__31162),
            .in1(N__25238),
            .in2(N__22081),
            .in3(N__31878),
            .lcout(\tok.n273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_107_LC_8_7_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_107_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_107_LC_8_7_0 .LUT_INIT=16'b1100010001000100;
    LogicCell40 \tok.i1_4_lut_adj_107_LC_8_7_0  (
            .in0(N__23302),
            .in1(N__31174),
            .in2(N__36303),
            .in3(N__23742),
            .lcout(\tok.n251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6854_2_lut_LC_8_7_1 .C_ON=1'b0;
    defparam \tok.i6854_2_lut_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6854_2_lut_LC_8_7_1 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \tok.i6854_2_lut_LC_8_7_1  (
            .in0(N__34614),
            .in1(N__28207),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\tok.n6620_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i296_4_lut_LC_8_7_2 .C_ON=1'b0;
    defparam \tok.i296_4_lut_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i296_4_lut_LC_8_7_2 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.i296_4_lut_LC_8_7_2  (
            .in0(N__36206),
            .in1(N__23741),
            .in2(N__21373),
            .in3(N__33185),
            .lcout(),
            .ltout(\tok.n167_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_124_LC_8_7_3 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_124_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_124_LC_8_7_3 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \tok.i1_3_lut_adj_124_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__21580),
            .in2(N__21574),
            .in3(N__24318),
            .lcout(\tok.n179_adj_730 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_165_LC_8_7_4 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_165_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_165_LC_8_7_4 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \tok.i308_4_lut_adj_165_LC_8_7_4  (
            .in0(N__21520),
            .in1(N__21571),
            .in2(N__36304),
            .in3(N__33186),
            .lcout(\tok.n186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i288_4_lut_4_lut_LC_8_7_5 .C_ON=1'b0;
    defparam \tok.i288_4_lut_4_lut_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i288_4_lut_4_lut_LC_8_7_5 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \tok.i288_4_lut_4_lut_LC_8_7_5  (
            .in0(N__31173),
            .in1(N__23259),
            .in2(N__21561),
            .in3(N__32071),
            .lcout(),
            .ltout(\tok.n209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6959_3_lut_LC_8_7_6 .C_ON=1'b0;
    defparam \tok.i6959_3_lut_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6959_3_lut_LC_8_7_6 .LUT_INIT=16'b0001000000010000;
    LogicCell40 \tok.i6959_3_lut_LC_8_7_6  (
            .in0(N__37113),
            .in1(N__34613),
            .in2(N__21535),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\tok.n6625_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_120_LC_8_7_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_120_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_120_LC_8_7_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \tok.i1_4_lut_adj_120_LC_8_7_7  (
            .in0(N__33184),
            .in1(N__35494),
            .in2(N__21532),
            .in3(N__21529),
            .lcout(\tok.n162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i320_4_lut_4_lut_4_lut_adj_85_LC_8_8_0 .C_ON=1'b0;
    defparam \tok.i320_4_lut_4_lut_4_lut_adj_85_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i320_4_lut_4_lut_4_lut_adj_85_LC_8_8_0 .LUT_INIT=16'b1000010110000000;
    LogicCell40 \tok.i320_4_lut_4_lut_4_lut_adj_85_LC_8_8_0  (
            .in0(N__31165),
            .in1(N__28225),
            .in2(N__32116),
            .in3(N__27022),
            .lcout(),
            .ltout(\tok.n168_adj_700_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6621_4_lut_LC_8_8_1 .C_ON=1'b0;
    defparam \tok.i6621_4_lut_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6621_4_lut_LC_8_8_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i6621_4_lut_LC_8_8_1  (
            .in0(N__32460),
            .in1(N__36341),
            .in2(N__21523),
            .in3(N__27346),
            .lcout(\tok.n6569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2525_2_lut_4_lut_LC_8_8_2 .C_ON=1'b0;
    defparam \tok.i2525_2_lut_4_lut_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2525_2_lut_4_lut_LC_8_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i2525_2_lut_4_lut_LC_8_8_2  (
            .in0(N__32034),
            .in1(N__34750),
            .in2(N__36256),
            .in3(N__33287),
            .lcout(\tok.n2548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i309_4_lut_LC_8_8_3 .C_ON=1'b0;
    defparam \tok.i309_4_lut_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i309_4_lut_LC_8_8_3 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \tok.i309_4_lut_LC_8_8_3  (
            .in0(N__27023),
            .in1(N__36102),
            .in2(N__21502),
            .in3(N__24556),
            .lcout(),
            .ltout(\tok.n179_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6997_4_lut_LC_8_8_4 .C_ON=1'b0;
    defparam \tok.i6997_4_lut_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6997_4_lut_LC_8_8_4 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \tok.i6997_4_lut_LC_8_8_4  (
            .in0(N__26875),
            .in1(N__35442),
            .in2(N__21691),
            .in3(N__34846),
            .lcout(\tok.n6546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i304_4_lut_4_lut_adj_315_LC_8_8_5 .C_ON=1'b0;
    defparam \tok.i304_4_lut_4_lut_adj_315_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i304_4_lut_4_lut_adj_315_LC_8_8_5 .LUT_INIT=16'b1010101000110000;
    LogicCell40 \tok.i304_4_lut_4_lut_adj_315_LC_8_8_5  (
            .in0(N__21607),
            .in1(N__32041),
            .in2(N__21682),
            .in3(N__31167),
            .lcout(\tok.n210_adj_816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i304_4_lut_4_lut_adj_317_LC_8_8_6 .C_ON=1'b0;
    defparam \tok.i304_4_lut_4_lut_adj_317_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i304_4_lut_4_lut_adj_317_LC_8_8_6 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \tok.i304_4_lut_4_lut_adj_317_LC_8_8_6  (
            .in0(N__31166),
            .in1(N__21642),
            .in2(N__32117),
            .in3(N__21859),
            .lcout(\tok.n210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_66_LC_8_8_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_66_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_66_LC_8_8_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i1_2_lut_adj_66_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__32033),
            .in2(_gnd_net_),
            .in3(N__31164),
            .lcout(\tok.n5_adj_682 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_234_LC_8_9_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_234_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_234_LC_8_9_0 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \tok.i1_4_lut_adj_234_LC_8_9_0  (
            .in0(N__26305),
            .in1(N__21586),
            .in2(N__32251),
            .in3(N__36098),
            .lcout(\tok.n258_adj_814 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i303_4_lut_adj_235_LC_8_9_1 .C_ON=1'b0;
    defparam \tok.i303_4_lut_adj_235_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i303_4_lut_adj_235_LC_8_9_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \tok.i303_4_lut_adj_235_LC_8_9_1  (
            .in0(N__35374),
            .in1(N__26410),
            .in2(N__23629),
            .in3(N__25894),
            .lcout(),
            .ltout(\tok.n252_adj_815_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_240_LC_8_9_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_240_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_240_LC_8_9_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_240_LC_8_9_2  (
            .in0(N__35376),
            .in1(N__21616),
            .in2(N__21610),
            .in3(N__34845),
            .lcout(\tok.n4_adj_818 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_adj_226_LC_8_9_3 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_226_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_226_LC_8_9_3 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \tok.i314_4_lut_adj_226_LC_8_9_3  (
            .in0(N__32247),
            .in1(N__21606),
            .in2(N__26392),
            .in3(N__37122),
            .lcout(\tok.n255_adj_808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_218_LC_8_9_4 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_218_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_218_LC_8_9_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_218_LC_8_9_4  (
            .in0(N__34821),
            .in1(N__36097),
            .in2(_gnd_net_),
            .in3(N__35373),
            .lcout(\tok.n872 ),
            .ltout(\tok.n872_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i306_4_lut_adj_239_LC_8_9_5 .C_ON=1'b0;
    defparam \tok.i306_4_lut_adj_239_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i306_4_lut_adj_239_LC_8_9_5 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \tok.i306_4_lut_adj_239_LC_8_9_5  (
            .in0(N__21814),
            .in1(N__37123),
            .in2(N__21808),
            .in3(N__23878),
            .lcout(),
            .ltout(\tok.n174_adj_817_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_242_LC_8_9_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_242_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_242_LC_8_9_6 .LUT_INIT=16'b0011001100010000;
    LogicCell40 \tok.i1_4_lut_adj_242_LC_8_9_6  (
            .in0(N__33217),
            .in1(N__34040),
            .in2(N__21805),
            .in3(N__21802),
            .lcout(\tok.n205_adj_820 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6888_2_lut_LC_8_10_0 .C_ON=1'b0;
    defparam \tok.i6888_2_lut_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6888_2_lut_LC_8_10_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i6888_2_lut_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__34035),
            .in2(_gnd_net_),
            .in3(N__26736),
            .lcout(\tok.n6365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_274_LC_8_10_1 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_274_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_274_LC_8_10_1 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \tok.i2_4_lut_adj_274_LC_8_10_1  (
            .in0(N__26585),
            .in1(N__26738),
            .in2(N__34101),
            .in3(N__21790),
            .lcout(),
            .ltout(\tok.n6_adj_843_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i10_LC_8_10_2 .C_ON=1'b0;
    defparam \tok.A_i10_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \tok.A_i10_LC_8_10_2 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \tok.A_i10_LC_8_10_2  (
            .in0(N__24574),
            .in1(N__25477),
            .in2(N__21781),
            .in3(N__21778),
            .lcout(\tok.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38496),
            .ce(N__25645),
            .sr(N__29261));
    defparam \tok.i6920_2_lut_LC_8_10_3 .C_ON=1'b0;
    defparam \tok.i6920_2_lut_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6920_2_lut_LC_8_10_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \tok.i6920_2_lut_LC_8_10_3  (
            .in0(N__34036),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27293),
            .lcout(),
            .ltout(\tok.n6440_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i310_4_lut_adj_271_LC_8_10_4 .C_ON=1'b0;
    defparam \tok.i310_4_lut_adj_271_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i310_4_lut_adj_271_LC_8_10_4 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.i310_4_lut_adj_271_LC_8_10_4  (
            .in0(N__33429),
            .in1(N__26737),
            .in2(N__21697),
            .in3(N__31213),
            .lcout(\tok.n215_adj_841 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6794_4_lut_LC_8_10_5 .C_ON=1'b0;
    defparam \tok.i6794_4_lut_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6794_4_lut_LC_8_10_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \tok.i6794_4_lut_LC_8_10_5  (
            .in0(N__26584),
            .in1(N__27294),
            .in2(N__23062),
            .in3(N__21865),
            .lcout(),
            .ltout(\tok.n6612_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i5_LC_8_10_6 .C_ON=1'b0;
    defparam \tok.A_i5_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \tok.A_i5_LC_8_10_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \tok.A_i5_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__25478),
            .in2(N__21694),
            .in3(N__23856),
            .lcout(\tok.A_low_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38496),
            .ce(N__25645),
            .sr(N__29261));
    defparam \tok.i310_4_lut_adj_58_LC_8_10_7 .C_ON=1'b0;
    defparam \tok.i310_4_lut_adj_58_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i310_4_lut_adj_58_LC_8_10_7 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \tok.i310_4_lut_adj_58_LC_8_10_7  (
            .in0(N__31212),
            .in1(N__33428),
            .in2(N__21901),
            .in3(N__32372),
            .lcout(\tok.n215_adj_672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_170_LC_8_11_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_170_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_170_LC_8_11_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_170_LC_8_11_0  (
            .in0(N__21823),
            .in1(N__35372),
            .in2(N__34791),
            .in3(N__21880),
            .lcout(),
            .ltout(\tok.n4_adj_769_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_171_LC_8_11_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_171_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_171_LC_8_11_1 .LUT_INIT=16'b0011000100110000;
    LogicCell40 \tok.i1_4_lut_adj_171_LC_8_11_1  (
            .in0(N__33291),
            .in1(N__33980),
            .in2(N__21868),
            .in3(N__23752),
            .lcout(\tok.n205_adj_770 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_231_LC_8_11_2 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_231_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_231_LC_8_11_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_231_LC_8_11_2  (
            .in0(N__35764),
            .in1(N__31955),
            .in2(_gnd_net_),
            .in3(N__31211),
            .lcout(\tok.n190 ),
            .ltout(\tok.n190_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_adj_161_LC_8_11_3 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_161_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_161_LC_8_11_3 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \tok.i314_4_lut_adj_161_LC_8_11_3  (
            .in0(N__26384),
            .in1(N__21858),
            .in2(N__21835),
            .in3(N__36797),
            .lcout(),
            .ltout(\tok.n255_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_166_LC_8_11_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_166_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_166_LC_8_11_4 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \tok.i1_4_lut_adj_166_LC_8_11_4  (
            .in0(N__35766),
            .in1(N__21832),
            .in2(N__21826),
            .in3(N__26315),
            .lcout(\tok.n258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6939_3_lut_4_lut_LC_8_11_5 .C_ON=1'b0;
    defparam \tok.i6939_3_lut_4_lut_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6939_3_lut_4_lut_LC_8_11_5 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \tok.i6939_3_lut_4_lut_LC_8_11_5  (
            .in0(N__22240),
            .in1(N__33979),
            .in2(N__24460),
            .in3(N__35765),
            .lcout(\tok.n6390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6787_2_lut_3_lut_LC_8_11_6 .C_ON=1'b0;
    defparam \tok.i6787_2_lut_3_lut_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6787_2_lut_3_lut_LC_8_11_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \tok.i6787_2_lut_3_lut_LC_8_11_6  (
            .in0(N__27541),
            .in1(N__35370),
            .in2(_gnd_net_),
            .in3(N__31210),
            .lcout(),
            .ltout(\tok.n6508_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i305_4_lut_adj_202_LC_8_11_7 .C_ON=1'b0;
    defparam \tok.i305_4_lut_adj_202_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i305_4_lut_adj_202_LC_8_11_7 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \tok.i305_4_lut_adj_202_LC_8_11_7  (
            .in0(N__35371),
            .in1(N__23400),
            .in2(N__21817),
            .in3(N__35763),
            .lcout(\tok.n213_adj_795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_98_i6_3_lut_LC_8_12_0 .C_ON=1'b0;
    defparam \tok.or_98_i6_3_lut_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.or_98_i6_3_lut_LC_8_12_0 .LUT_INIT=16'b1010111111111010;
    LogicCell40 \tok.or_98_i6_3_lut_LC_8_12_0  (
            .in0(N__27543),
            .in1(_gnd_net_),
            .in2(N__36322),
            .in3(N__37063),
            .lcout(),
            .ltout(\tok.n207_adj_771_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i305_4_lut_LC_8_12_1 .C_ON=1'b0;
    defparam \tok.i305_4_lut_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i305_4_lut_LC_8_12_1 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \tok.i305_4_lut_LC_8_12_1  (
            .in0(N__22057),
            .in1(N__36279),
            .in2(N__22042),
            .in3(N__35375),
            .lcout(\tok.n213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6836_3_lut_4_lut_LC_8_12_2 .C_ON=1'b0;
    defparam \tok.i6836_3_lut_4_lut_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6836_3_lut_4_lut_LC_8_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \tok.i6836_3_lut_4_lut_LC_8_12_2  (
            .in0(N__36554),
            .in1(N__33064),
            .in2(N__36320),
            .in3(N__30954),
            .lcout(\tok.n6583 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i318_4_lut_adj_179_LC_8_12_3 .C_ON=1'b0;
    defparam \tok.i318_4_lut_adj_179_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i318_4_lut_adj_179_LC_8_12_3 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.i318_4_lut_adj_179_LC_8_12_3  (
            .in0(N__22028),
            .in1(N__34523),
            .in2(N__23677),
            .in3(N__36280),
            .lcout(),
            .ltout(\tok.n207_adj_776_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6823_4_lut_4_lut_LC_8_12_4 .C_ON=1'b0;
    defparam \tok.i6823_4_lut_4_lut_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6823_4_lut_4_lut_LC_8_12_4 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \tok.i6823_4_lut_4_lut_LC_8_12_4  (
            .in0(N__31897),
            .in1(N__21946),
            .in2(N__21940),
            .in3(N__24287),
            .lcout(),
            .ltout(\tok.n6529_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i306_4_lut_adj_188_LC_8_12_5 .C_ON=1'b0;
    defparam \tok.i306_4_lut_adj_188_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i306_4_lut_adj_188_LC_8_12_5 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \tok.i306_4_lut_adj_188_LC_8_12_5  (
            .in0(N__37064),
            .in1(N__24223),
            .in2(N__21937),
            .in3(N__21934),
            .lcout(\tok.n174_adj_785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2641_2_lut_3_lut_LC_8_12_6 .C_ON=1'b0;
    defparam \tok.i2641_2_lut_3_lut_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2641_2_lut_3_lut_LC_8_12_6 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \tok.i2641_2_lut_3_lut_LC_8_12_6  (
            .in0(N__27542),
            .in1(_gnd_net_),
            .in2(N__36321),
            .in3(N__33065),
            .lcout(\tok.n2665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_261_LC_8_12_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_261_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_261_LC_8_12_7 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_261_LC_8_12_7  (
            .in0(N__30955),
            .in1(_gnd_net_),
            .in2(N__33223),
            .in3(N__31896),
            .lcout(\tok.n847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i369_4_lut_LC_8_13_0 .C_ON=1'b0;
    defparam \tok.i369_4_lut_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.i369_4_lut_LC_8_13_0 .LUT_INIT=16'b1111000000010001;
    LogicCell40 \tok.i369_4_lut_LC_8_13_0  (
            .in0(N__26504),
            .in1(N__30533),
            .in2(N__22264),
            .in3(N__36147),
            .lcout(\tok.n229_adj_861 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6662_3_lut_LC_8_13_1 .C_ON=1'b0;
    defparam \tok.i6662_3_lut_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6662_3_lut_LC_8_13_1 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \tok.i6662_3_lut_LC_8_13_1  (
            .in0(N__35379),
            .in1(_gnd_net_),
            .in2(N__34102),
            .in3(N__31086),
            .lcout(\tok.n6320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6895_2_lut_LC_8_13_2 .C_ON=1'b0;
    defparam \tok.i6895_2_lut_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6895_2_lut_LC_8_13_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \tok.i6895_2_lut_LC_8_13_2  (
            .in0(N__22228),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34045),
            .lcout(),
            .ltout(\tok.n6380_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i310_4_lut_adj_46_LC_8_13_3 .C_ON=1'b0;
    defparam \tok.i310_4_lut_adj_46_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.i310_4_lut_adj_46_LC_8_13_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.i310_4_lut_adj_46_LC_8_13_3  (
            .in0(N__33475),
            .in1(N__32220),
            .in2(N__22108),
            .in3(N__31087),
            .lcout(),
            .ltout(\tok.n215_adj_656_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6745_4_lut_LC_8_13_4 .C_ON=1'b0;
    defparam \tok.i6745_4_lut_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6745_4_lut_LC_8_13_4 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.i6745_4_lut_LC_8_13_4  (
            .in0(N__26932),
            .in1(N__24565),
            .in2(N__22105),
            .in3(N__35380),
            .lcout(\tok.n6544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i338_4_lut_LC_8_13_5 .C_ON=1'b0;
    defparam \tok.i338_4_lut_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.i338_4_lut_LC_8_13_5 .LUT_INIT=16'b0100000001110011;
    LogicCell40 \tok.i338_4_lut_LC_8_13_5  (
            .in0(N__33219),
            .in1(N__34842),
            .in2(N__22093),
            .in3(N__22102),
            .lcout(\tok.n256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_225_LC_8_13_6 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_225_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_225_LC_8_13_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i1_2_lut_adj_225_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__34041),
            .in2(_gnd_net_),
            .in3(N__35378),
            .lcout(\tok.n4_adj_719 ),
            .ltout(\tok.n4_adj_719_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_227_LC_8_13_7 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_227_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_227_LC_8_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \tok.i4_4_lut_adj_227_LC_8_13_7  (
            .in0(N__33218),
            .in1(N__34841),
            .in2(N__22084),
            .in3(N__36571),
            .lcout(\tok.n10_adj_809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i309_4_lut_adj_330_LC_8_14_0 .C_ON=1'b0;
    defparam \tok.i309_4_lut_adj_330_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \tok.i309_4_lut_adj_330_LC_8_14_0 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i309_4_lut_adj_330_LC_8_14_0  (
            .in0(N__22066),
            .in1(N__36145),
            .in2(N__24555),
            .in3(N__23988),
            .lcout(\tok.n179_adj_888 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6938_3_lut_4_lut_LC_8_14_1 .C_ON=1'b0;
    defparam \tok.i6938_3_lut_4_lut_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6938_3_lut_4_lut_LC_8_14_1 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \tok.i6938_3_lut_4_lut_LC_8_14_1  (
            .in0(N__36146),
            .in1(N__24452),
            .in2(N__34103),
            .in3(N__37465),
            .lcout(),
            .ltout(\tok.n6404_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6821_4_lut_LC_8_14_2 .C_ON=1'b0;
    defparam \tok.i6821_4_lut_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6821_4_lut_LC_8_14_2 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \tok.i6821_4_lut_LC_8_14_2  (
            .in0(N__35382),
            .in1(N__26927),
            .in2(N__22402),
            .in3(N__23890),
            .lcout(),
            .ltout(\tok.n6550_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6999_4_lut_LC_8_14_3 .C_ON=1'b0;
    defparam \tok.i6999_4_lut_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6999_4_lut_LC_8_14_3 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \tok.i6999_4_lut_LC_8_14_3  (
            .in0(N__22399),
            .in1(N__35383),
            .in2(N__22393),
            .in3(N__34795),
            .lcout(\tok.n6549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6863_2_lut_3_lut_4_lut_LC_8_14_4 .C_ON=1'b0;
    defparam \tok.i6863_2_lut_3_lut_4_lut_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6863_2_lut_3_lut_4_lut_LC_8_14_4 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \tok.i6863_2_lut_3_lut_4_lut_LC_8_14_4  (
            .in0(N__34046),
            .in1(N__37065),
            .in2(N__24461),
            .in3(N__30323),
            .lcout(\tok.n6442 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6937_3_lut_4_lut_LC_8_14_5 .C_ON=1'b0;
    defparam \tok.i6937_3_lut_4_lut_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6937_3_lut_4_lut_LC_8_14_5 .LUT_INIT=16'b0000000010100010;
    LogicCell40 \tok.i6937_3_lut_4_lut_LC_8_14_5  (
            .in0(N__36143),
            .in1(N__24448),
            .in2(N__30074),
            .in3(N__34047),
            .lcout(\tok.n6419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6674_3_lut_4_lut_LC_8_14_6 .C_ON=1'b0;
    defparam \tok.i6674_3_lut_4_lut_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6674_3_lut_4_lut_LC_8_14_6 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \tok.i6674_3_lut_4_lut_LC_8_14_6  (
            .in0(N__34048),
            .in1(N__36144),
            .in2(N__24462),
            .in3(N__23987),
            .lcout(),
            .ltout(\tok.n6337_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6771_4_lut_LC_8_14_7 .C_ON=1'b0;
    defparam \tok.i6771_4_lut_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6771_4_lut_LC_8_14_7 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \tok.i6771_4_lut_LC_8_14_7  (
            .in0(N__26926),
            .in1(N__22372),
            .in2(N__22360),
            .in3(N__35381),
            .lcout(\tok.n6538 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i5_LC_9_1_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i5_LC_9_1_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i5_LC_9_1_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i5_LC_9_1_0  (
            .in0(N__28753),
            .in1(N__22540),
            .in2(_gnd_net_),
            .in3(N__22278),
            .lcout(\tok.C_stk.tail_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38461),
            .ce(N__28919),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i6152_3_lut_LC_9_1_1 .C_ON=1'b0;
    defparam \tok.C_stk.i6152_3_lut_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i6152_3_lut_LC_9_1_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i6152_3_lut_LC_9_1_1  (
            .in0(N__22548),
            .in1(N__28122),
            .in2(_gnd_net_),
            .in3(N__22348),
            .lcout(),
            .ltout(\tok.C_stk.n6236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i5_LC_9_1_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i5_LC_9_1_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i5_LC_9_1_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i5_LC_9_1_2  (
            .in0(N__28051),
            .in1(N__27940),
            .in2(N__22318),
            .in3(N__22315),
            .lcout(\tok.c_stk_r_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38461),
            .ce(N__28919),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i13_LC_9_1_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i13_LC_9_1_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i13_LC_9_1_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i13_LC_9_1_3  (
            .in0(N__22549),
            .in1(_gnd_net_),
            .in2(N__22531),
            .in3(N__28748),
            .lcout(\tok.tail_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38461),
            .ce(N__28919),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i21_LC_9_1_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i21_LC_9_1_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i21_LC_9_1_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i21_LC_9_1_4  (
            .in0(N__28749),
            .in1(N__22519),
            .in2(_gnd_net_),
            .in3(N__22539),
            .lcout(\tok.C_stk.tail_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38461),
            .ce(N__28919),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i29_LC_9_1_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i29_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i29_LC_9_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i29_LC_9_1_5  (
            .in0(N__22527),
            .in1(N__22510),
            .in2(_gnd_net_),
            .in3(N__28750),
            .lcout(\tok.tail_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38461),
            .ce(N__28919),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i37_LC_9_1_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i37_LC_9_1_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i37_LC_9_1_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i37_LC_9_1_6  (
            .in0(N__28751),
            .in1(N__24618),
            .in2(_gnd_net_),
            .in3(N__22518),
            .lcout(\tok.C_stk.tail_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38461),
            .ce(N__28919),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i45_LC_9_1_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i45_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i45_LC_9_1_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i45_LC_9_1_7  (
            .in0(N__25033),
            .in1(N__22509),
            .in2(_gnd_net_),
            .in3(N__28752),
            .lcout(\tok.tail_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38461),
            .ce(N__28919),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i2_LC_9_2_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i2_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i2_LC_9_2_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i2_LC_9_2_0  (
            .in0(N__28739),
            .in1(N__22699),
            .in2(_gnd_net_),
            .in3(N__22434),
            .lcout(\tok.C_stk.tail_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38465),
            .ce(N__28905),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i6161_3_lut_LC_9_2_1 .C_ON=1'b0;
    defparam \tok.C_stk.i6161_3_lut_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i6161_3_lut_LC_9_2_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i6161_3_lut_LC_9_2_1  (
            .in0(N__22410),
            .in1(N__28103),
            .in2(_gnd_net_),
            .in3(N__22496),
            .lcout(),
            .ltout(\tok.C_stk.n6245_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i2_LC_9_2_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i2_LC_9_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i2_LC_9_2_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i2_LC_9_2_2  (
            .in0(N__28050),
            .in1(N__27933),
            .in2(N__22468),
            .in3(N__22465),
            .lcout(\tok.c_stk_r_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38465),
            .ce(N__28905),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i10_LC_9_2_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i10_LC_9_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i10_LC_9_2_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i10_LC_9_2_3  (
            .in0(N__22411),
            .in1(_gnd_net_),
            .in2(N__22690),
            .in3(N__28736),
            .lcout(\tok.tail_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38465),
            .ce(N__28905),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i18_LC_9_2_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i18_LC_9_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i18_LC_9_2_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i18_LC_9_2_4  (
            .in0(N__28737),
            .in1(N__22678),
            .in2(_gnd_net_),
            .in3(N__22698),
            .lcout(\tok.C_stk.tail_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38465),
            .ce(N__28905),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i26_LC_9_2_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i26_LC_9_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i26_LC_9_2_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i26_LC_9_2_5  (
            .in0(N__22686),
            .in1(N__22669),
            .in2(_gnd_net_),
            .in3(N__28738),
            .lcout(\tok.tail_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38465),
            .ce(N__28905),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i34_LC_9_2_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i34_LC_9_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i34_LC_9_2_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i34_LC_9_2_6  (
            .in0(N__28740),
            .in1(N__24856),
            .in2(_gnd_net_),
            .in3(N__22677),
            .lcout(\tok.C_stk.tail_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38465),
            .ce(N__28905),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i42_LC_9_2_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i42_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i42_LC_9_2_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i42_LC_9_2_7  (
            .in0(N__27781),
            .in1(N__22668),
            .in2(_gnd_net_),
            .in3(N__28741),
            .lcout(\tok.tail_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38465),
            .ce(N__28905),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i3_LC_9_3_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i3_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i3_LC_9_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i3_LC_9_3_0  (
            .in0(N__28679),
            .in1(N__22558),
            .in2(_gnd_net_),
            .in3(N__22585),
            .lcout(\tok.C_stk.tail_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38470),
            .ce(N__28921),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i6158_3_lut_LC_9_3_1 .C_ON=1'b0;
    defparam \tok.C_stk.i6158_3_lut_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i6158_3_lut_LC_9_3_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.C_stk.i6158_3_lut_LC_9_3_1  (
            .in0(N__28102),
            .in1(N__22566),
            .in2(_gnd_net_),
            .in3(N__22655),
            .lcout(),
            .ltout(\tok.C_stk.n6242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i3_LC_9_3_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i3_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i3_LC_9_3_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i3_LC_9_3_2  (
            .in0(N__28049),
            .in1(N__27925),
            .in2(N__22624),
            .in3(N__22621),
            .lcout(\tok.c_stk_r_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38470),
            .ce(N__28921),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i11_LC_9_3_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i11_LC_9_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i11_LC_9_3_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i11_LC_9_3_3  (
            .in0(N__22972),
            .in1(N__22567),
            .in2(_gnd_net_),
            .in3(N__28675),
            .lcout(\tok.C_stk.tail_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38470),
            .ce(N__28921),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i19_LC_9_3_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i19_LC_9_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i19_LC_9_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i19_LC_9_3_4  (
            .in0(N__28676),
            .in1(N__22963),
            .in2(_gnd_net_),
            .in3(N__22557),
            .lcout(\tok.C_stk.tail_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38470),
            .ce(N__28921),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i27_LC_9_3_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i27_LC_9_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i27_LC_9_3_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i27_LC_9_3_5  (
            .in0(N__22971),
            .in1(N__22954),
            .in2(_gnd_net_),
            .in3(N__28677),
            .lcout(\tok.C_stk.tail_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38470),
            .ce(N__28921),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i35_LC_9_3_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i35_LC_9_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i35_LC_9_3_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.C_stk.tail_i0_i35_LC_9_3_6  (
            .in0(N__28678),
            .in1(N__22962),
            .in2(_gnd_net_),
            .in3(N__24636),
            .lcout(\tok.C_stk.tail_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38470),
            .ce(N__28921),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i43_LC_9_3_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i43_LC_9_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i43_LC_9_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i43_LC_9_3_7  (
            .in0(N__24840),
            .in1(N__22953),
            .in2(_gnd_net_),
            .in3(N__28680),
            .lcout(\tok.C_stk.tail_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38470),
            .ce(N__28921),
            .sr(_gnd_net_));
    defparam \tok.i6605_4_lut_LC_9_4_0 .C_ON=1'b0;
    defparam \tok.i6605_4_lut_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6605_4_lut_LC_9_4_0 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.i6605_4_lut_LC_9_4_0  (
            .in0(N__22915),
            .in1(N__24995),
            .in2(N__24934),
            .in3(N__22869),
            .lcout(),
            .ltout(\tok.n6291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i124_4_lut_adj_133_LC_9_4_1 .C_ON=1'b0;
    defparam \tok.i124_4_lut_adj_133_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.i124_4_lut_adj_133_LC_9_4_1 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \tok.i124_4_lut_adj_133_LC_9_4_1  (
            .in0(N__32120),
            .in1(N__22779),
            .in2(N__22744),
            .in3(N__24933),
            .lcout(),
            .ltout(\tok.n80_adj_735_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i126_4_lut_adj_136_LC_9_4_2 .C_ON=1'b0;
    defparam \tok.i126_4_lut_adj_136_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i126_4_lut_adj_136_LC_9_4_2 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \tok.i126_4_lut_adj_136_LC_9_4_2  (
            .in0(N__35517),
            .in1(N__22735),
            .in2(N__22741),
            .in3(N__31328),
            .lcout(\tok.n89_adj_736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_132_LC_9_4_3 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_132_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_132_LC_9_4_3 .LUT_INIT=16'b0101000010001000;
    LogicCell40 \tok.i125_4_lut_adj_132_LC_9_4_3  (
            .in0(N__31327),
            .in1(N__24929),
            .in2(N__23296),
            .in3(N__33264),
            .lcout(),
            .ltout(\tok.n83_adj_725_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6641_2_lut_3_lut_LC_9_4_4 .C_ON=1'b0;
    defparam \tok.i6641_2_lut_3_lut_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6641_2_lut_3_lut_LC_9_4_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i6641_2_lut_3_lut_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(N__36299),
            .in2(N__22738),
            .in3(N__32119),
            .lcout(\tok.n6287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_139_LC_9_4_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_139_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_139_LC_9_4_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_139_LC_9_4_5  (
            .in0(N__24996),
            .in1(N__25797),
            .in2(N__29723),
            .in3(N__22729),
            .lcout(n92),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i307_3_lut_3_lut_3_lut_LC_9_4_6 .C_ON=1'b0;
    defparam \tok.i307_3_lut_3_lut_3_lut_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i307_3_lut_3_lut_3_lut_LC_9_4_6 .LUT_INIT=16'b0011001111101110;
    LogicCell40 \tok.i307_3_lut_3_lut_3_lut_LC_9_4_6  (
            .in0(N__33263),
            .in1(N__32118),
            .in2(_gnd_net_),
            .in3(N__31326),
            .lcout(\tok.n180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_147_LC_9_4_7 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_147_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_147_LC_9_4_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i2_4_lut_adj_147_LC_9_4_7  (
            .in0(N__31329),
            .in1(N__34820),
            .in2(N__26511),
            .in3(N__36533),
            .lcout(\tok.n4926 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2664_4_lut_LC_9_5_0 .C_ON=1'b0;
    defparam \tok.i2664_4_lut_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2664_4_lut_LC_9_5_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i2664_4_lut_LC_9_5_0  (
            .in0(N__33283),
            .in1(N__36296),
            .in2(N__34839),
            .in3(N__35516),
            .lcout(),
            .ltout(\tok.n2692_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i359_4_lut_LC_9_5_1 .C_ON=1'b0;
    defparam \tok.i359_4_lut_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i359_4_lut_LC_9_5_1 .LUT_INIT=16'b0000111110001000;
    LogicCell40 \tok.i359_4_lut_LC_9_5_1  (
            .in0(N__23008),
            .in1(N__25875),
            .in2(N__23023),
            .in3(N__31303),
            .lcout(\tok.n217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_rep_28_2_lut_LC_9_5_2 .C_ON=1'b0;
    defparam \tok.i1_rep_28_2_lut_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_rep_28_2_lut_LC_9_5_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i1_rep_28_2_lut_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__35515),
            .in2(_gnd_net_),
            .in3(N__34785),
            .lcout(\tok.n7154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_LC_9_5_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_LC_9_5_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.i1_2_lut_3_lut_LC_9_5_3  (
            .in0(N__36295),
            .in1(N__32098),
            .in2(_gnd_net_),
            .in3(N__33282),
            .lcout(\tok.n815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_rep_332_2_lut_LC_9_5_4 .C_ON=1'b0;
    defparam \tok.i1_rep_332_2_lut_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_rep_332_2_lut_LC_9_5_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i1_rep_332_2_lut_LC_9_5_4  (
            .in0(N__32099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37110),
            .lcout(\tok.n7458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_3_lut_4_lut_LC_9_5_6 .C_ON=1'b0;
    defparam \tok.i2_2_lut_3_lut_4_lut_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_3_lut_4_lut_LC_9_5_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \tok.i2_2_lut_3_lut_4_lut_LC_9_5_6  (
            .in0(N__31302),
            .in1(N__34786),
            .in2(N__33301),
            .in3(N__32107),
            .lcout(\tok.n6_adj_701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_138_LC_9_5_7 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_138_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_138_LC_9_5_7 .LUT_INIT=16'b0000110000001101;
    LogicCell40 \tok.i2_4_lut_adj_138_LC_9_5_7  (
            .in0(N__22996),
            .in1(N__22990),
            .in2(N__33489),
            .in3(N__32100),
            .lcout(\tok.n239_adj_738 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_4_lut_LC_9_6_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_4_lut_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_4_lut_LC_9_6_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_4_lut_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__34106),
            .in2(_gnd_net_),
            .in3(N__36298),
            .lcout(\tok.n864 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2679_3_lut_3_lut_LC_9_6_1 .C_ON=1'b0;
    defparam \tok.i2679_3_lut_3_lut_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2679_3_lut_3_lut_LC_9_6_1 .LUT_INIT=16'b1011101101110111;
    LogicCell40 \tok.i2679_3_lut_3_lut_LC_9_6_1  (
            .in0(N__32123),
            .in1(N__33288),
            .in2(_gnd_net_),
            .in3(N__31249),
            .lcout(\tok.n2679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_336_LC_9_6_2 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_336_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_336_LC_9_6_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i1_2_lut_adj_336_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__36297),
            .in2(_gnd_net_),
            .in3(N__34797),
            .lcout(\tok.n5_adj_821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_334_LC_9_6_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_334_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_334_LC_9_6_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_334_LC_9_6_3  (
            .in0(N__34105),
            .in1(N__25368),
            .in2(_gnd_net_),
            .in3(N__29408),
            .lcout(\tok.n17 ),
            .ltout(\tok.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_243_LC_9_6_4 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_243_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_243_LC_9_6_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \tok.i2_4_lut_adj_243_LC_9_6_4  (
            .in0(N__23106),
            .in1(N__23092),
            .in2(N__23086),
            .in3(N__25737),
            .lcout(\tok.n2559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6809_4_lut_LC_9_6_5 .C_ON=1'b0;
    defparam \tok.i6809_4_lut_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6809_4_lut_LC_9_6_5 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \tok.i6809_4_lut_LC_9_6_5  (
            .in0(N__32551),
            .in1(N__32601),
            .in2(N__23083),
            .in3(N__27393),
            .lcout(),
            .ltout(\tok.n6562_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i315_4_lut_LC_9_6_6 .C_ON=1'b0;
    defparam \tok.i315_4_lut_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i315_4_lut_LC_9_6_6 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \tok.i315_4_lut_LC_9_6_6  (
            .in0(N__35520),
            .in1(N__23074),
            .in2(N__23065),
            .in3(N__34799),
            .lcout(\tok.n338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6867_4_lut_LC_9_6_7 .C_ON=1'b0;
    defparam \tok.i6867_4_lut_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6867_4_lut_LC_9_6_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \tok.i6867_4_lut_LC_9_6_7  (
            .in0(N__34798),
            .in1(N__23470),
            .in2(N__25110),
            .in3(N__35521),
            .lcout(\tok.n6637 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_123_LC_9_7_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_123_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_123_LC_9_7_0 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \tok.i1_4_lut_adj_123_LC_9_7_0  (
            .in0(N__23047),
            .in1(N__29458),
            .in2(N__23227),
            .in3(N__35468),
            .lcout(),
            .ltout(\tok.n197_adj_729_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_125_LC_9_7_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_125_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_125_LC_9_7_1 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \tok.i1_4_lut_adj_125_LC_9_7_1  (
            .in0(N__36219),
            .in1(N__23041),
            .in2(N__23314),
            .in3(N__23311),
            .lcout(\tok.n203_adj_731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2521_2_lut_LC_9_7_2 .C_ON=1'b0;
    defparam \tok.i2521_2_lut_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2521_2_lut_LC_9_7_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i2521_2_lut_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__23549),
            .in2(_gnd_net_),
            .in3(N__34800),
            .lcout(\tok.n2544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_3_lut_LC_9_7_3 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_3_lut_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_3_lut_LC_9_7_3 .LUT_INIT=16'b0101010110100000;
    LogicCell40 \tok.i1_3_lut_4_lut_3_lut_LC_9_7_3  (
            .in0(N__35467),
            .in1(_gnd_net_),
            .in2(N__36305),
            .in3(N__33290),
            .lcout(\tok.n256_adj_749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2598_rep_349_2_lut_LC_9_7_4 .C_ON=1'b0;
    defparam \tok.i2598_rep_349_2_lut_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2598_rep_349_2_lut_LC_9_7_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i2598_rep_349_2_lut_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__37137),
            .in2(_gnd_net_),
            .in3(N__34802),
            .lcout(),
            .ltout(\tok.n7475_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6981_4_lut_4_lut_LC_9_7_5 .C_ON=1'b0;
    defparam \tok.i6981_4_lut_4_lut_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6981_4_lut_4_lut_LC_9_7_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \tok.i6981_4_lut_4_lut_LC_9_7_5  (
            .in0(N__35466),
            .in1(N__23295),
            .in2(N__23263),
            .in3(N__32125),
            .lcout(\tok.n6645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6984_4_lut_LC_9_7_6 .C_ON=1'b0;
    defparam \tok.i6984_4_lut_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6984_4_lut_LC_9_7_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \tok.i6984_4_lut_LC_9_7_6  (
            .in0(N__23260),
            .in1(N__37136),
            .in2(N__23239),
            .in3(N__34801),
            .lcout(\tok.n6628 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i337_4_lut_adj_145_LC_9_7_7 .C_ON=1'b0;
    defparam \tok.i337_4_lut_adj_145_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i337_4_lut_adj_145_LC_9_7_7 .LUT_INIT=16'b0000110001010101;
    LogicCell40 \tok.i337_4_lut_adj_145_LC_9_7_7  (
            .in0(N__23217),
            .in1(N__32124),
            .in2(N__37891),
            .in3(N__33289),
            .lcout(\tok.n241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_112_LC_9_8_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_112_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_112_LC_9_8_0 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \tok.i1_4_lut_adj_112_LC_9_8_0  (
            .in0(N__36287),
            .in1(N__27129),
            .in2(N__37126),
            .in3(N__23329),
            .lcout(),
            .ltout(\tok.n284_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_113_LC_9_8_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_113_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_113_LC_9_8_1 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \tok.i1_4_lut_adj_113_LC_9_8_1  (
            .in0(N__36230),
            .in1(N__23131),
            .in2(N__23122),
            .in3(N__26023),
            .lcout(),
            .ltout(\tok.n244_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_116_LC_9_8_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_116_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_116_LC_9_8_2 .LUT_INIT=16'b0011001111110010;
    LogicCell40 \tok.i1_4_lut_adj_116_LC_9_8_2  (
            .in0(N__25672),
            .in1(N__27461),
            .in2(N__23380),
            .in3(N__34076),
            .lcout(),
            .ltout(\tok.n4_adj_720_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i2_LC_9_8_3 .C_ON=1'b0;
    defparam \tok.A_i2_LC_9_8_3 .SEQ_MODE=4'b1010;
    defparam \tok.A_i2_LC_9_8_3 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \tok.A_i2_LC_9_8_3  (
            .in0(N__25481),
            .in1(N__23553),
            .in2(N__23377),
            .in3(N__27577),
            .lcout(\tok.A_low_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38491),
            .ce(N__25607),
            .sr(N__29204));
    defparam \tok.inv_105_i2_1_lut_LC_9_8_4 .C_ON=1'b0;
    defparam \tok.inv_105_i2_1_lut_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i2_1_lut_LC_9_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i2_1_lut_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27457),
            .lcout(\tok.n145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_108_LC_9_8_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_108_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_108_LC_9_8_5 .LUT_INIT=16'b1111111100001101;
    LogicCell40 \tok.i1_4_lut_adj_108_LC_9_8_5  (
            .in0(N__27090),
            .in1(N__36285),
            .in2(N__34813),
            .in3(N__23365),
            .lcout(),
            .ltout(\tok.n4_adj_714_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_4_lut_adj_316_LC_9_8_6 .C_ON=1'b0;
    defparam \tok.i2_4_lut_4_lut_adj_316_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_4_lut_adj_316_LC_9_8_6 .LUT_INIT=16'b0011000000110010;
    LogicCell40 \tok.i2_4_lut_4_lut_adj_316_LC_9_8_6  (
            .in0(N__36286),
            .in1(N__23359),
            .in2(N__23332),
            .in3(N__32042),
            .lcout(\tok.n218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6795_2_lut_4_lut_LC_9_8_7 .C_ON=1'b0;
    defparam \tok.i6795_2_lut_4_lut_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6795_2_lut_4_lut_LC_9_8_7 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \tok.i6795_2_lut_4_lut_LC_9_8_7  (
            .in0(N__34075),
            .in1(N__37069),
            .in2(N__27509),
            .in3(N__36284),
            .lcout(\tok.n6525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i57_4_lut_3_lut_LC_9_9_0 .C_ON=1'b0;
    defparam \tok.i57_4_lut_3_lut_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i57_4_lut_3_lut_LC_9_9_0 .LUT_INIT=16'b0101101010100000;
    LogicCell40 \tok.i57_4_lut_3_lut_LC_9_9_0  (
            .in0(N__31206),
            .in1(_gnd_net_),
            .in2(N__33281),
            .in3(N__31973),
            .lcout(\tok.n39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6628_4_lut_4_lut_LC_9_9_1 .C_ON=1'b0;
    defparam \tok.i6628_4_lut_4_lut_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6628_4_lut_4_lut_LC_9_9_1 .LUT_INIT=16'b1000000100000000;
    LogicCell40 \tok.i6628_4_lut_4_lut_LC_9_9_1  (
            .in0(N__31974),
            .in1(N__33196),
            .in2(N__36323),
            .in3(N__31207),
            .lcout(),
            .ltout(\tok.n6269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i58_4_lut_LC_9_9_2 .C_ON=1'b0;
    defparam \tok.i58_4_lut_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i58_4_lut_LC_9_9_2 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \tok.i58_4_lut_LC_9_9_2  (
            .in0(N__23323),
            .in1(N__35455),
            .in2(N__23317),
            .in3(N__36293),
            .lcout(\tok.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_104_LC_9_9_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_104_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_104_LC_9_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i1_2_lut_adj_104_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__31958),
            .in2(_gnd_net_),
            .in3(N__33192),
            .lcout(\tok.n6_adj_676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6765_4_lut_LC_9_9_4 .C_ON=1'b0;
    defparam \tok.i6765_4_lut_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6765_4_lut_LC_9_9_4 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \tok.i6765_4_lut_LC_9_9_4  (
            .in0(N__31960),
            .in1(N__23653),
            .in2(N__23617),
            .in3(N__23638),
            .lcout(\tok.n6486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6783_4_lut_LC_9_9_5 .C_ON=1'b0;
    defparam \tok.i6783_4_lut_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6783_4_lut_LC_9_9_5 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.i6783_4_lut_LC_9_9_5  (
            .in0(N__23612),
            .in1(N__23581),
            .in2(N__23569),
            .in3(N__31959),
            .lcout(\tok.n6510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i336_4_lut_LC_9_9_6 .C_ON=1'b0;
    defparam \tok.i336_4_lut_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i336_4_lut_LC_9_9_6 .LUT_INIT=16'b0000010110001000;
    LogicCell40 \tok.i336_4_lut_LC_9_9_6  (
            .in0(N__31208),
            .in1(N__27471),
            .in2(N__23554),
            .in3(N__37073),
            .lcout(\tok.n208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6824_4_lut_4_lut_4_lut_LC_9_9_7 .C_ON=1'b0;
    defparam \tok.i6824_4_lut_4_lut_4_lut_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6824_4_lut_4_lut_4_lut_LC_9_9_7 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \tok.i6824_4_lut_4_lut_4_lut_LC_9_9_7  (
            .in0(N__34697),
            .in1(N__33197),
            .in2(N__32094),
            .in3(N__31209),
            .lcout(\tok.n6589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i17_4_lut_LC_9_10_0 .C_ON=1'b0;
    defparam \tok.i17_4_lut_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i17_4_lut_LC_9_10_0 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \tok.i17_4_lut_LC_9_10_0  (
            .in0(N__34062),
            .in1(N__33635),
            .in2(N__32605),
            .in3(N__32077),
            .lcout(),
            .ltout(\tok.n6_adj_728_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_128_LC_9_10_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_128_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_128_LC_9_10_1 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \tok.i1_4_lut_adj_128_LC_9_10_1  (
            .in0(N__23440),
            .in1(N__32550),
            .in2(N__23428),
            .in3(N__34063),
            .lcout(),
            .ltout(\tok.n200_adj_732_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_130_LC_9_10_2 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_130_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_130_LC_9_10_2 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \tok.i2_4_lut_adj_130_LC_9_10_2  (
            .in0(N__35519),
            .in1(N__34107),
            .in2(N__23425),
            .in3(N__23422),
            .lcout(\tok.n6_adj_733 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6778_2_lut_LC_9_10_3 .C_ON=1'b0;
    defparam \tok.i6778_2_lut_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6778_2_lut_LC_9_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i6778_2_lut_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__32469),
            .in2(_gnd_net_),
            .in3(N__23401),
            .lcout(\tok.n6501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6769_3_lut_LC_9_10_4 .C_ON=1'b0;
    defparam \tok.i6769_3_lut_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6769_3_lut_LC_9_10_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \tok.i6769_3_lut_LC_9_10_4  (
            .in0(N__34061),
            .in1(N__33634),
            .in2(_gnd_net_),
            .in3(N__31130),
            .lcout(\tok.n6484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i318_4_lut_adj_230_LC_9_10_5 .C_ON=1'b0;
    defparam \tok.i318_4_lut_adj_230_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i318_4_lut_adj_230_LC_9_10_5 .LUT_INIT=16'b1100111000000010;
    LogicCell40 \tok.i318_4_lut_adj_230_LC_9_10_5  (
            .in0(N__28334),
            .in1(N__36292),
            .in2(N__34803),
            .in3(N__23675),
            .lcout(),
            .ltout(\tok.n207_adj_811_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6834_4_lut_4_lut_LC_9_10_6 .C_ON=1'b0;
    defparam \tok.i6834_4_lut_4_lut_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6834_4_lut_4_lut_LC_9_10_6 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \tok.i6834_4_lut_4_lut_LC_9_10_6  (
            .in0(N__24324),
            .in1(N__23863),
            .in2(N__23881),
            .in3(N__32076),
            .lcout(\tok.n6481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i305_4_lut_adj_229_LC_9_10_7 .C_ON=1'b0;
    defparam \tok.i305_4_lut_adj_229_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i305_4_lut_adj_229_LC_9_10_7 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \tok.i305_4_lut_adj_229_LC_9_10_7  (
            .in0(N__32407),
            .in1(N__35518),
            .in2(N__23872),
            .in3(N__36291),
            .lcout(\tok.n213_adj_810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i318_4_lut_LC_9_11_0 .C_ON=1'b0;
    defparam \tok.i318_4_lut_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i318_4_lut_LC_9_11_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \tok.i318_4_lut_LC_9_11_0  (
            .in0(N__35779),
            .in1(N__34682),
            .in2(N__23857),
            .in3(N__23676),
            .lcout(),
            .ltout(\tok.n207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6822_4_lut_LC_9_11_1 .C_ON=1'b0;
    defparam \tok.i6822_4_lut_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6822_4_lut_LC_9_11_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i6822_4_lut_LC_9_11_1  (
            .in0(N__24323),
            .in1(N__27058),
            .in2(N__23767),
            .in3(N__24472),
            .lcout(),
            .ltout(\tok.n6572_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i306_4_lut_LC_9_11_2 .C_ON=1'b0;
    defparam \tok.i306_4_lut_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i306_4_lut_LC_9_11_2 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \tok.i306_4_lut_LC_9_11_2  (
            .in0(N__24219),
            .in1(N__23764),
            .in2(N__23755),
            .in3(N__36796),
            .lcout(\tok.n174_adj_768 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_3_lut_LC_9_11_3 .C_ON=1'b0;
    defparam \tok.i2_2_lut_3_lut_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_3_lut_LC_9_11_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \tok.i2_2_lut_3_lut_LC_9_11_3  (
            .in0(N__34680),
            .in1(N__23732),
            .in2(_gnd_net_),
            .in3(N__31943),
            .lcout(\tok.n26_adj_763 ),
            .ltout(\tok.n26_adj_763_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i318_4_lut_adj_203_LC_9_11_4 .C_ON=1'b0;
    defparam \tok.i318_4_lut_adj_203_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i318_4_lut_adj_203_LC_9_11_4 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \tok.i318_4_lut_adj_203_LC_9_11_4  (
            .in0(N__25993),
            .in1(N__35767),
            .in2(N__23656),
            .in3(N__34681),
            .lcout(),
            .ltout(\tok.n207_adj_796_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6816_4_lut_4_lut_LC_9_11_5 .C_ON=1'b0;
    defparam \tok.i6816_4_lut_4_lut_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6816_4_lut_4_lut_LC_9_11_5 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \tok.i6816_4_lut_4_lut_LC_9_11_5  (
            .in0(N__24322),
            .in1(N__24232),
            .in2(N__24226),
            .in3(N__31944),
            .lcout(),
            .ltout(\tok.n6505_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i306_4_lut_adj_214_LC_9_11_6 .C_ON=1'b0;
    defparam \tok.i306_4_lut_adj_214_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i306_4_lut_adj_214_LC_9_11_6 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \tok.i306_4_lut_adj_214_LC_9_11_6  (
            .in0(N__24218),
            .in1(N__24028),
            .in2(N__24202),
            .in3(N__36795),
            .lcout(\tok.n174_adj_803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_4_lut_4_lut_LC_9_11_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_4_lut_4_lut_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_4_lut_4_lut_LC_9_11_7 .LUT_INIT=16'b0000011100000110;
    LogicCell40 \tok.i1_2_lut_4_lut_4_lut_LC_9_11_7  (
            .in0(N__31112),
            .in1(N__31942),
            .in2(N__34796),
            .in3(N__33198),
            .lcout(\tok.n867 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i320_4_lut_4_lut_4_lut_LC_9_12_0 .C_ON=1'b0;
    defparam \tok.i320_4_lut_4_lut_4_lut_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i320_4_lut_4_lut_4_lut_LC_9_12_0 .LUT_INIT=16'b1100000000100010;
    LogicCell40 \tok.i320_4_lut_4_lut_4_lut_LC_9_12_0  (
            .in0(N__24169),
            .in1(N__31885),
            .in2(N__37645),
            .in3(N__30787),
            .lcout(\tok.n168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6943_3_lut_4_lut_LC_9_12_1 .C_ON=1'b0;
    defparam \tok.i6943_3_lut_4_lut_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6943_3_lut_4_lut_LC_9_12_1 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \tok.i6943_3_lut_4_lut_LC_9_12_1  (
            .in0(N__36229),
            .in1(N__24454),
            .in2(N__34096),
            .in3(N__29619),
            .lcout(\tok.n6360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i304_4_lut_4_lut_LC_9_12_2 .C_ON=1'b0;
    defparam \tok.i304_4_lut_4_lut_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i304_4_lut_4_lut_LC_9_12_2 .LUT_INIT=16'b1010101000110000;
    LogicCell40 \tok.i304_4_lut_4_lut_LC_9_12_2  (
            .in0(N__26349),
            .in1(N__31884),
            .in2(N__24061),
            .in3(N__30786),
            .lcout(\tok.n210_adj_802 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i10_1_lut_LC_9_12_3 .C_ON=1'b0;
    defparam \tok.inv_105_i10_1_lut_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i10_1_lut_LC_9_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i10_1_lut_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26758),
            .lcout(\tok.n316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6909_2_lut_LC_9_12_4 .C_ON=1'b0;
    defparam \tok.i6909_2_lut_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6909_2_lut_LC_9_12_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.i6909_2_lut_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__30058),
            .in2(_gnd_net_),
            .in3(N__34026),
            .lcout(),
            .ltout(\tok.n6409_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i310_4_lut_adj_329_LC_9_12_5 .C_ON=1'b0;
    defparam \tok.i310_4_lut_adj_329_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i310_4_lut_adj_329_LC_9_12_5 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \tok.i310_4_lut_adj_329_LC_9_12_5  (
            .in0(N__30788),
            .in1(N__33484),
            .in2(N__24004),
            .in3(N__23999),
            .lcout(\tok.n215_adj_887 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i309_4_lut_adj_272_LC_9_13_0 .C_ON=1'b0;
    defparam \tok.i309_4_lut_adj_272_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.i309_4_lut_adj_272_LC_9_13_0 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i309_4_lut_adj_272_LC_9_13_0  (
            .in0(N__24604),
            .in1(N__36154),
            .in2(N__24552),
            .in3(N__26768),
            .lcout(\tok.n179_adj_842 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6936_3_lut_4_lut_LC_9_13_1 .C_ON=1'b0;
    defparam \tok.i6936_3_lut_4_lut_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6936_3_lut_4_lut_LC_9_13_1 .LUT_INIT=16'b0010000000100010;
    LogicCell40 \tok.i6936_3_lut_4_lut_LC_9_13_1  (
            .in0(N__36155),
            .in1(N__34070),
            .in2(N__30345),
            .in3(N__24441),
            .lcout(),
            .ltout(\tok.n6433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6655_4_lut_LC_9_13_2 .C_ON=1'b0;
    defparam \tok.i6655_4_lut_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6655_4_lut_LC_9_13_2 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \tok.i6655_4_lut_LC_9_13_2  (
            .in0(N__35457),
            .in1(N__26933),
            .in2(N__24598),
            .in3(N__24595),
            .lcout(),
            .ltout(\tok.n6602_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6987_4_lut_LC_9_13_3 .C_ON=1'b0;
    defparam \tok.i6987_4_lut_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.i6987_4_lut_LC_9_13_3 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \tok.i6987_4_lut_LC_9_13_3  (
            .in0(N__34675),
            .in1(N__24583),
            .in2(N__24577),
            .in3(N__35459),
            .lcout(\tok.n6601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6940_3_lut_4_lut_LC_9_13_4 .C_ON=1'b0;
    defparam \tok.i6940_3_lut_4_lut_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6940_3_lut_4_lut_LC_9_13_4 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \tok.i6940_3_lut_4_lut_LC_9_13_4  (
            .in0(N__34069),
            .in1(N__36153),
            .in2(N__24459),
            .in3(N__26767),
            .lcout(\tok.n6375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i309_4_lut_adj_47_LC_9_13_5 .C_ON=1'b0;
    defparam \tok.i309_4_lut_adj_47_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.i309_4_lut_adj_47_LC_9_13_5 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \tok.i309_4_lut_adj_47_LC_9_13_5  (
            .in0(N__36156),
            .in1(N__24343),
            .in2(N__24553),
            .in3(N__32231),
            .lcout(),
            .ltout(\tok.n179_adj_657_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6980_4_lut_LC_9_13_6 .C_ON=1'b0;
    defparam \tok.i6980_4_lut_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6980_4_lut_LC_9_13_6 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \tok.i6980_4_lut_LC_9_13_6  (
            .in0(N__35458),
            .in1(N__24493),
            .in2(N__24487),
            .in3(N__34676),
            .lcout(\tok.n6543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i305_3_lut_LC_9_13_7 .C_ON=1'b0;
    defparam \tok.i305_3_lut_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.i305_3_lut_LC_9_13_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.i305_3_lut_LC_9_13_7  (
            .in0(N__30532),
            .in1(N__35456),
            .in2(_gnd_net_),
            .in3(N__31088),
            .lcout(\tok.n464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6874_2_lut_3_lut_4_lut_LC_9_14_2 .C_ON=1'b0;
    defparam \tok.i6874_2_lut_3_lut_4_lut_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6874_2_lut_3_lut_4_lut_LC_9_14_2 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \tok.i6874_2_lut_3_lut_4_lut_LC_9_14_2  (
            .in0(N__34071),
            .in1(N__37127),
            .in2(N__24458),
            .in3(N__26792),
            .lcout(\tok.n6382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i40_LC_11_1_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i40_LC_11_1_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i40_LC_11_1_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i40_LC_11_1_0  (
            .in0(N__24801),
            .in1(N__24681),
            .in2(_gnd_net_),
            .in3(N__28692),
            .lcout(tail_40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38466),
            .ce(N__28920),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i32_LC_11_1_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i32_LC_11_1_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i32_LC_11_1_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i32_LC_11_1_2  (
            .in0(N__24706),
            .in1(N__24651),
            .in2(_gnd_net_),
            .in3(N__28691),
            .lcout(\tok.C_stk.tail_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38466),
            .ce(N__28920),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i48_LC_11_1_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i48_LC_11_1_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i48_LC_11_1_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i48_LC_11_1_3  (
            .in0(N__28693),
            .in1(N__24784),
            .in2(_gnd_net_),
            .in3(N__24705),
            .lcout(tail_48_adj_900),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38466),
            .ce(N__28920),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i16_LC_11_1_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i16_LC_11_1_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i16_LC_11_1_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i16_LC_11_1_4  (
            .in0(N__24652),
            .in1(N__24697),
            .in2(_gnd_net_),
            .in3(N__28689),
            .lcout(\tok.C_stk.tail_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38466),
            .ce(N__28920),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i24_LC_11_1_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i24_LC_11_1_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i24_LC_11_1_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i24_LC_11_1_6  (
            .in0(N__24682),
            .in1(N__24663),
            .in2(_gnd_net_),
            .in3(N__28690),
            .lcout(tail_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38466),
            .ce(N__28920),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i49_LC_11_2_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i49_LC_11_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i49_LC_11_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i49_LC_11_2_0  (
            .in0(N__24766),
            .in1(N__25186),
            .in2(_gnd_net_),
            .in3(N__28623),
            .lcout(tail_49_adj_899),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38471),
            .ce(N__28889),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i51_LC_11_2_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i51_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i51_LC_11_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i51_LC_11_2_2  (
            .in0(N__24817),
            .in1(N__24640),
            .in2(_gnd_net_),
            .in3(N__28625),
            .lcout(tail_51),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38471),
            .ce(N__28889),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i54_LC_11_2_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i54_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i54_LC_11_2_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i54_LC_11_2_3  (
            .in0(N__28628),
            .in1(N__24721),
            .in2(_gnd_net_),
            .in3(N__28134),
            .lcout(\tok.tail_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38471),
            .ce(N__28889),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i53_LC_11_2_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i53_LC_11_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i53_LC_11_2_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i53_LC_11_2_4  (
            .in0(N__25012),
            .in1(N__24622),
            .in2(_gnd_net_),
            .in3(N__28627),
            .lcout(\tok.tail_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38471),
            .ce(N__28889),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i52_LC_11_2_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i52_LC_11_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i52_LC_11_2_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i52_LC_11_2_5  (
            .in0(N__28626),
            .in1(N__24733),
            .in2(_gnd_net_),
            .in3(N__24871),
            .lcout(\tok.tail_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38471),
            .ce(N__28889),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i50_LC_11_2_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i50_LC_11_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i50_LC_11_2_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i50_LC_11_2_6  (
            .in0(N__24855),
            .in1(N__27760),
            .in2(_gnd_net_),
            .in3(N__28624),
            .lcout(\tok.tail_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38471),
            .ce(N__28889),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i55_LC_11_2_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i55_LC_11_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i55_LC_11_2_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i55_LC_11_2_7  (
            .in0(N__28629),
            .in1(N__28501),
            .in2(_gnd_net_),
            .in3(N__28939),
            .lcout(\tok.tail_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38471),
            .ce(N__28889),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i59_LC_11_3_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i59_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i59_LC_11_3_0 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \tok.C_stk.tail_i0_i59_LC_11_3_0  (
            .in0(N__28607),
            .in1(N__24816),
            .in2(N__24841),
            .in3(N__28834),
            .lcout(tail_59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38475),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i56_LC_11_3_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i56_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i56_LC_11_3_1 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \tok.C_stk.tail_i0_i56_LC_11_3_1  (
            .in0(N__28832),
            .in1(N__24780),
            .in2(N__24805),
            .in3(N__28606),
            .lcout(tail_56),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38475),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2545_2_lut_4_lut_LC_11_3_2 .C_ON=1'b0;
    defparam \tok.i2545_2_lut_4_lut_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2545_2_lut_4_lut_LC_11_3_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \tok.i2545_2_lut_4_lut_LC_11_3_2  (
            .in0(N__25068),
            .in1(N__25050),
            .in2(N__29838),
            .in3(N__25247),
            .lcout(C_stk_delta_1),
            .ltout(C_stk_delta_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i57_LC_11_3_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i57_LC_11_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i57_LC_11_3_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \tok.C_stk.tail_i0_i57_LC_11_3_3  (
            .in0(N__28833),
            .in1(N__25209),
            .in2(N__24769),
            .in3(N__24762),
            .lcout(tail_57),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38475),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i60_LC_11_3_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i60_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i60_LC_11_3_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \tok.C_stk.tail_i0_i60_LC_11_3_4  (
            .in0(N__28608),
            .in1(N__24732),
            .in2(N__24750),
            .in3(N__28830),
            .lcout(\tok.tail_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38475),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i62_LC_11_3_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i62_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i62_LC_11_3_5 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \tok.C_stk.tail_i0_i62_LC_11_3_5  (
            .in0(N__28831),
            .in1(N__24717),
            .in2(N__28159),
            .in3(N__28610),
            .lcout(\tok.tail_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38475),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i427_2_lut_4_lut_LC_11_3_6 .C_ON=1'b0;
    defparam \tok.i427_2_lut_4_lut_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.i427_2_lut_4_lut_LC_11_3_6 .LUT_INIT=16'b0011001110110011;
    LogicCell40 \tok.i427_2_lut_4_lut_LC_11_3_6  (
            .in0(N__25069),
            .in1(N__25051),
            .in2(N__29839),
            .in3(N__25248),
            .lcout(rd_7__N_373),
            .ltout(rd_7__N_373_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i61_LC_11_3_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i61_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i61_LC_11_3_7 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \tok.C_stk.tail_i0_i61_LC_11_3_7  (
            .in0(N__25029),
            .in1(N__25011),
            .in2(N__25015),
            .in3(N__28609),
            .lcout(\tok.tail_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38475),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i1_LC_11_4_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i1_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i1_LC_11_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i1_LC_11_4_0  (
            .in0(N__28618),
            .in1(N__24901),
            .in2(_gnd_net_),
            .in3(N__24928),
            .lcout(\tok.C_stk.tail_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38480),
            .ce(N__28873),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i6164_3_lut_LC_11_4_1 .C_ON=1'b0;
    defparam \tok.C_stk.i6164_3_lut_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i6164_3_lut_LC_11_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i6164_3_lut_LC_11_4_1  (
            .in0(N__24909),
            .in1(N__28117),
            .in2(_gnd_net_),
            .in3(N__25000),
            .lcout(),
            .ltout(\tok.C_stk.n6248_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i1_LC_11_4_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i1_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i1_LC_11_4_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i1_LC_11_4_2  (
            .in0(N__28053),
            .in1(N__27941),
            .in2(N__24970),
            .in3(N__24967),
            .lcout(c_stk_r_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38480),
            .ce(N__28873),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i9_LC_11_4_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i9_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i9_LC_11_4_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i9_LC_11_4_3  (
            .in0(N__24910),
            .in1(_gnd_net_),
            .in2(N__24892),
            .in3(N__28622),
            .lcout(tail_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38480),
            .ce(N__28873),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i17_LC_11_4_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i17_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i17_LC_11_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i17_LC_11_4_4  (
            .in0(N__28617),
            .in1(N__24880),
            .in2(_gnd_net_),
            .in3(N__24900),
            .lcout(\tok.C_stk.tail_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38480),
            .ce(N__28873),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i25_LC_11_4_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i25_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i25_LC_11_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i25_LC_11_4_5  (
            .in0(N__24888),
            .in1(N__25195),
            .in2(_gnd_net_),
            .in3(N__28619),
            .lcout(tail_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38480),
            .ce(N__28873),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i33_LC_11_4_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i33_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i33_LC_11_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.C_stk.tail_i0_i33_LC_11_4_6  (
            .in0(N__28620),
            .in1(N__24879),
            .in2(_gnd_net_),
            .in3(N__25185),
            .lcout(\tok.C_stk.tail_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38480),
            .ce(N__28873),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i41_LC_11_4_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i41_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i41_LC_11_4_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i41_LC_11_4_7  (
            .in0(N__25210),
            .in1(N__25194),
            .in2(_gnd_net_),
            .in3(N__28621),
            .lcout(tail_41),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38480),
            .ce(N__28873),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_144_LC_11_5_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_144_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_144_LC_11_5_0 .LUT_INIT=16'b1010000011111100;
    LogicCell40 \tok.i1_4_lut_adj_144_LC_11_5_0  (
            .in0(N__25171),
            .in1(N__36318),
            .in2(N__34838),
            .in3(N__37095),
            .lcout(\tok.n265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_134_LC_11_5_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_134_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_134_LC_11_5_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i1_2_lut_adj_134_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__35507),
            .in2(_gnd_net_),
            .in3(N__33252),
            .lcout(\tok.n156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i338_4_lut_adj_143_LC_11_5_2 .C_ON=1'b0;
    defparam \tok.i338_4_lut_adj_143_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i338_4_lut_adj_143_LC_11_5_2 .LUT_INIT=16'b0000001110100000;
    LogicCell40 \tok.i338_4_lut_adj_143_LC_11_5_2  (
            .in0(N__31300),
            .in1(N__36319),
            .in2(N__33298),
            .in3(N__34811),
            .lcout(),
            .ltout(\tok.n211_adj_741_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_3_lut_LC_11_5_3 .C_ON=1'b0;
    defparam \tok.i1_3_lut_3_lut_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_3_lut_LC_11_5_3 .LUT_INIT=16'b0101010111110101;
    LogicCell40 \tok.i1_3_lut_3_lut_LC_11_5_3  (
            .in0(N__37096),
            .in1(_gnd_net_),
            .in2(N__25165),
            .in3(N__32133),
            .lcout(),
            .ltout(\tok.n277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_150_LC_11_5_4 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_150_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_150_LC_11_5_4 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \tok.i2_4_lut_adj_150_LC_11_5_4  (
            .in0(N__31301),
            .in1(N__35509),
            .in2(N__25162),
            .in3(N__25159),
            .lcout(\tok.n6_adj_748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i361_4_lut_LC_11_5_5 .C_ON=1'b0;
    defparam \tok.i361_4_lut_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i361_4_lut_LC_11_5_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \tok.i361_4_lut_LC_11_5_5  (
            .in0(N__26863),
            .in1(N__32132),
            .in2(N__25138),
            .in3(N__33253),
            .lcout(),
            .ltout(\tok.n238_adj_855_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_295_LC_11_5_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_295_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_295_LC_11_5_6 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \tok.i1_4_lut_adj_295_LC_11_5_6  (
            .in0(N__35508),
            .in1(N__36317),
            .in2(N__25123),
            .in3(N__25075),
            .lcout(\tok.n4_adj_859 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_289_LC_11_5_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_289_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_289_LC_11_5_7 .LUT_INIT=16'b1101010111011101;
    LogicCell40 \tok.i1_4_lut_adj_289_LC_11_5_7  (
            .in0(N__37094),
            .in1(N__34781),
            .in2(N__25111),
            .in3(N__31299),
            .lcout(\tok.n298_adj_856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_i0_LC_11_6_0 .C_ON=1'b0;
    defparam \tok.depth_i0_LC_11_6_0 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i0_LC_11_6_0 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \tok.depth_i0_LC_11_6_0  (
            .in0(N__29346),
            .in1(_gnd_net_),
            .in2(N__29818),
            .in3(_gnd_net_),
            .lcout(\tok.depth_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38487),
            .ce(),
            .sr(N__29168));
    defparam \tok.i1_2_lut_adj_288_LC_11_6_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_288_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_288_LC_11_6_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.i1_2_lut_adj_288_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__29814),
            .in2(_gnd_net_),
            .in3(N__29345),
            .lcout(),
            .ltout(\tok.n53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7015_4_lut_LC_11_6_2 .C_ON=1'b0;
    defparam \tok.i7015_4_lut_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i7015_4_lut_LC_11_6_2 .LUT_INIT=16'b0011001100110111;
    LogicCell40 \tok.i7015_4_lut_LC_11_6_2  (
            .in0(N__25378),
            .in1(N__25409),
            .in2(N__25654),
            .in3(N__29305),
            .lcout(\tok.n992 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_3__I_0_389_i2_2_lut_LC_11_6_3 .C_ON=1'b0;
    defparam \tok.depth_3__I_0_389_i2_2_lut_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.depth_3__I_0_389_i2_2_lut_LC_11_6_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.depth_3__I_0_389_i2_2_lut_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__29759),
            .in2(_gnd_net_),
            .in3(N__28979),
            .lcout(),
            .ltout(\tok.n2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_287_LC_11_6_4 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_287_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_287_LC_11_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i4_4_lut_adj_287_LC_11_6_4  (
            .in0(N__31312),
            .in1(N__26500),
            .in2(N__25522),
            .in3(N__25216),
            .lcout(\tok.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2566_2_lut_LC_11_6_5 .C_ON=1'b0;
    defparam \tok.i2566_2_lut_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2566_2_lut_LC_11_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i2566_2_lut_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__29344),
            .in2(_gnd_net_),
            .in3(N__29395),
            .lcout(\tok.n174 ),
            .ltout(\tok.n174_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_i2_LC_11_6_6 .C_ON=1'b0;
    defparam \tok.depth_i2_LC_11_6_6 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i2_LC_11_6_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \tok.depth_i2_LC_11_6_6  (
            .in0(N__28980),
            .in1(_gnd_net_),
            .in2(N__25381),
            .in3(N__29287),
            .lcout(\tok.depth_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38487),
            .ce(),
            .sr(N__29168));
    defparam \tok.i6106_2_lut_LC_11_6_7 .C_ON=1'b0;
    defparam \tok.i6106_2_lut_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6106_2_lut_LC_11_6_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i6106_2_lut_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__25377),
            .in2(_gnd_net_),
            .in3(N__29396),
            .lcout(\tok.n6189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_118_LC_11_7_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_118_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_118_LC_11_7_0 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_adj_118_LC_11_7_0  (
            .in0(N__37087),
            .in1(N__35506),
            .in2(N__29851),
            .in3(N__36301),
            .lcout(\tok.n6_adj_722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i965_3_lut_3_lut_LC_11_7_1 .C_ON=1'b0;
    defparam \tok.i965_3_lut_3_lut_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i965_3_lut_3_lut_LC_11_7_1 .LUT_INIT=16'b0111011101100110;
    LogicCell40 \tok.i965_3_lut_3_lut_LC_11_7_1  (
            .in0(N__36300),
            .in1(N__32092),
            .in2(_gnd_net_),
            .in3(N__33249),
            .lcout(),
            .ltout(\tok.n10_adj_773_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_174_LC_11_7_2 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_174_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_174_LC_11_7_2 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \tok.i2_4_lut_adj_174_LC_11_7_2  (
            .in0(N__33250),
            .in1(N__25828),
            .in2(N__25819),
            .in3(N__31307),
            .lcout(),
            .ltout(\tok.n6146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_178_LC_11_7_3 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_178_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_178_LC_11_7_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i4_4_lut_adj_178_LC_11_7_3  (
            .in0(N__25660),
            .in1(N__28973),
            .in2(N__25816),
            .in3(N__37086),
            .lcout(\tok.n86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i349_4_lut_4_lut_LC_11_7_4 .C_ON=1'b0;
    defparam \tok.i349_4_lut_4_lut_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i349_4_lut_4_lut_LC_11_7_4 .LUT_INIT=16'b1000010100000101;
    LogicCell40 \tok.i349_4_lut_4_lut_LC_11_7_4  (
            .in0(N__33251),
            .in1(N__36302),
            .in2(N__37128),
            .in3(N__31308),
            .lcout(),
            .ltout(\tok.n369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_109_LC_11_7_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_109_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_109_LC_11_7_5 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \tok.i1_4_lut_adj_109_LC_11_7_5  (
            .in0(N__31309),
            .in1(N__25738),
            .in2(N__25705),
            .in3(N__34812),
            .lcout(),
            .ltout(\tok.n233_adj_716_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_114_LC_11_7_6 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_114_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_114_LC_11_7_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \tok.i2_4_lut_adj_114_LC_11_7_6  (
            .in0(N__32093),
            .in1(N__25702),
            .in2(N__25690),
            .in3(N__25687),
            .lcout(\tok.n6156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_adj_177_LC_11_7_7 .C_ON=1'b0;
    defparam \tok.i2_2_lut_adj_177_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_adj_177_LC_11_7_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i2_2_lut_adj_177_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__29847),
            .in2(_gnd_net_),
            .in3(N__29757),
            .lcout(\tok.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6858_4_lut_LC_11_8_0 .C_ON=1'b0;
    defparam \tok.i6858_4_lut_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6858_4_lut_LC_11_8_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \tok.i6858_4_lut_LC_11_8_0  (
            .in0(N__26496),
            .in1(N__26842),
            .in2(N__26074),
            .in3(N__31314),
            .lcout(\tok.n6639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6753_2_lut_LC_11_8_1 .C_ON=1'b0;
    defparam \tok.i6753_2_lut_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6753_2_lut_LC_11_8_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \tok.i6753_2_lut_LC_11_8_1  (
            .in0(N__28189),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32115),
            .lcout(),
            .ltout(\tok.n6653_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6982_4_lut_LC_11_8_2 .C_ON=1'b0;
    defparam \tok.i6982_4_lut_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6982_4_lut_LC_11_8_2 .LUT_INIT=16'b0010001010100000;
    LogicCell40 \tok.i6982_4_lut_LC_11_8_2  (
            .in0(N__26130),
            .in1(N__26098),
            .in2(N__26080),
            .in3(N__34809),
            .lcout(),
            .ltout(\tok.n6646_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i341_4_lut_LC_11_8_3 .C_ON=1'b0;
    defparam \tok.i341_4_lut_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i341_4_lut_LC_11_8_3 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \tok.i341_4_lut_LC_11_8_3  (
            .in0(N__35514),
            .in1(N__27091),
            .in2(N__26077),
            .in3(N__33190),
            .lcout(\tok.n280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_221_LC_11_8_4 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_221_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_221_LC_11_8_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i1_2_lut_adj_221_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__34808),
            .in2(_gnd_net_),
            .in3(N__35510),
            .lcout(\tok.n6167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6989_4_lut_LC_11_8_5 .C_ON=1'b0;
    defparam \tok.i6989_4_lut_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6989_4_lut_LC_11_8_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \tok.i6989_4_lut_LC_11_8_5  (
            .in0(N__31315),
            .in1(N__26065),
            .in2(N__26053),
            .in3(N__33191),
            .lcout(),
            .ltout(\tok.n6638_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6963_4_lut_LC_11_8_6 .C_ON=1'b0;
    defparam \tok.i6963_4_lut_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6963_4_lut_LC_11_8_6 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \tok.i6963_4_lut_LC_11_8_6  (
            .in0(N__26038),
            .in1(N__26032),
            .in2(N__26026),
            .in3(N__37068),
            .lcout(\tok.n6636 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i345_3_lut_LC_11_8_7 .C_ON=1'b0;
    defparam \tok.i345_3_lut_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i345_3_lut_LC_11_8_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \tok.i345_3_lut_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__31313),
            .in2(N__35524),
            .in3(N__26014),
            .lcout(\tok.n367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i317_4_lut_adj_210_LC_11_9_0 .C_ON=1'b0;
    defparam \tok.i317_4_lut_adj_210_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i317_4_lut_adj_210_LC_11_9_0 .LUT_INIT=16'b0001000110100000;
    LogicCell40 \tok.i317_4_lut_adj_210_LC_11_9_0  (
            .in0(N__36988),
            .in1(N__30026),
            .in2(N__25992),
            .in3(N__31188),
            .lcout(),
            .ltout(\tok.n177_adj_799_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i303_4_lut_adj_213_LC_11_9_1 .C_ON=1'b0;
    defparam \tok.i303_4_lut_adj_213_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i303_4_lut_adj_213_LC_11_9_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \tok.i303_4_lut_adj_213_LC_11_9_1  (
            .in0(N__25882),
            .in1(N__25840),
            .in2(N__25831),
            .in3(N__35485),
            .lcout(),
            .ltout(\tok.n252_adj_801_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_215_LC_11_9_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_215_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_215_LC_11_9_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_215_LC_11_9_2  (
            .in0(N__35486),
            .in1(N__26266),
            .in2(N__26395),
            .in3(N__34816),
            .lcout(\tok.n4_adj_804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_223_LC_11_9_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_223_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_223_LC_11_9_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \tok.i1_2_lut_adj_223_LC_11_9_3  (
            .in0(N__34815),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36986),
            .lcout(\tok.n5_adj_745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i314_4_lut_adj_198_LC_11_9_4 .C_ON=1'b0;
    defparam \tok.i314_4_lut_adj_198_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i314_4_lut_adj_198_LC_11_9_4 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \tok.i314_4_lut_adj_198_LC_11_9_4  (
            .in0(N__36987),
            .in1(N__26445),
            .in2(N__26391),
            .in3(N__26350),
            .lcout(),
            .ltout(\tok.n255_adj_793_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_212_LC_11_9_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_212_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_212_LC_11_9_5 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \tok.i1_4_lut_adj_212_LC_11_9_5  (
            .in0(N__26446),
            .in1(N__26287),
            .in2(N__26269),
            .in3(N__36258),
            .lcout(\tok.n258_adj_800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_263_LC_11_9_6 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_263_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_263_LC_11_9_6 .LUT_INIT=16'b1000000000001000;
    LogicCell40 \tok.i2_4_lut_adj_263_LC_11_9_6  (
            .in0(N__36985),
            .in1(N__34814),
            .in2(N__29412),
            .in3(N__31187),
            .lcout(),
            .ltout(\tok.n6162_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_264_LC_11_9_7 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_264_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_264_LC_11_9_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \tok.i4_4_lut_adj_264_LC_11_9_7  (
            .in0(N__26483),
            .in1(N__26259),
            .in2(N__26236),
            .in3(N__36257),
            .lcout(\tok.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_LC_11_10_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_LC_11_10_0 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_LC_11_10_0  (
            .in0(N__34094),
            .in1(N__35488),
            .in2(N__32594),
            .in3(N__27536),
            .lcout(),
            .ltout(\tok.n865_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6776_4_lut_LC_11_10_1 .C_ON=1'b0;
    defparam \tok.i6776_4_lut_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6776_4_lut_LC_11_10_1 .LUT_INIT=16'b1010000010101000;
    LogicCell40 \tok.i6776_4_lut_LC_11_10_1  (
            .in0(N__32547),
            .in1(N__30027),
            .in2(N__26233),
            .in3(N__32585),
            .lcout(\tok.n6496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_3_lut_adj_260_LC_11_10_2 .C_ON=1'b0;
    defparam \tok.i2_2_lut_3_lut_adj_260_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_3_lut_adj_260_LC_11_10_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i2_2_lut_3_lut_adj_260_LC_11_10_2  (
            .in0(N__36259),
            .in1(N__34817),
            .in2(_gnd_net_),
            .in3(N__33257),
            .lcout(\tok.n222 ),
            .ltout(\tok.n222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i11_3_lut_4_lut_LC_11_10_3 .C_ON=1'b0;
    defparam \tok.i11_3_lut_4_lut_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i11_3_lut_4_lut_LC_11_10_3 .LUT_INIT=16'b0111010011111100;
    LogicCell40 \tok.i11_3_lut_4_lut_LC_11_10_3  (
            .in0(N__34818),
            .in1(N__27083),
            .in2(N__26230),
            .in3(N__36260),
            .lcout(\tok.n245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_208_LC_11_10_4 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_208_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_208_LC_11_10_4 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \tok.i308_4_lut_adj_208_LC_11_10_4  (
            .in0(N__36261),
            .in1(N__29890),
            .in2(N__26641),
            .in3(N__33258),
            .lcout(),
            .ltout(\tok.n186_adj_798_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i315_4_lut_adj_216_LC_11_10_5 .C_ON=1'b0;
    defparam \tok.i315_4_lut_adj_216_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i315_4_lut_adj_216_LC_11_10_5 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \tok.i315_4_lut_adj_216_LC_11_10_5  (
            .in0(N__34819),
            .in1(N__35489),
            .in2(N__26629),
            .in3(N__26626),
            .lcout(),
            .ltout(\tok.n338_adj_805_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6759_4_lut_LC_11_10_6 .C_ON=1'b0;
    defparam \tok.i6759_4_lut_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6759_4_lut_LC_11_10_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \tok.i6759_4_lut_LC_11_10_6  (
            .in0(N__30028),
            .in1(N__26608),
            .in2(N__26530),
            .in3(N__26416),
            .lcout(\tok.n6608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_286_LC_11_10_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_286_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_286_LC_11_10_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.i1_2_lut_adj_286_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__37043),
            .in2(_gnd_net_),
            .in3(N__31229),
            .lcout(\tok.n4_adj_712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_36_LC_11_11_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_36_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_36_LC_11_11_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_36_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__31744),
            .in2(_gnd_net_),
            .in3(N__33102),
            .lcout(\tok.n219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_256_LC_11_11_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_256_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_256_LC_11_11_1 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_adj_256_LC_11_11_1  (
            .in0(N__31745),
            .in1(N__31225),
            .in2(N__27558),
            .in3(N__35481),
            .lcout(\tok.n190_adj_792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_217_LC_11_11_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_217_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_217_LC_11_11_2 .LUT_INIT=16'b0100010101000100;
    LogicCell40 \tok.i1_4_lut_adj_217_LC_11_11_2  (
            .in0(N__34078),
            .in1(N__26434),
            .in2(N__33299),
            .in3(N__26425),
            .lcout(\tok.n205_adj_806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i317_4_lut_adj_233_LC_11_11_3 .C_ON=1'b0;
    defparam \tok.i317_4_lut_adj_233_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i317_4_lut_adj_233_LC_11_11_3 .LUT_INIT=16'b0000001110100000;
    LogicCell40 \tok.i317_4_lut_adj_233_LC_11_11_3  (
            .in0(N__28338),
            .in1(N__37455),
            .in2(N__36936),
            .in3(N__31226),
            .lcout(\tok.n177_adj_813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_220_LC_11_11_4 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_220_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_220_LC_11_11_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_220_LC_11_11_4  (
            .in0(N__33259),
            .in1(_gnd_net_),
            .in2(N__31957),
            .in3(N__36784),
            .lcout(\tok.n821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2575_2_lut_LC_11_11_5 .C_ON=1'b0;
    defparam \tok.i2575_2_lut_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2575_2_lut_LC_11_11_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i2575_2_lut_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__34077),
            .in2(_gnd_net_),
            .in3(N__37456),
            .lcout(),
            .ltout(\tok.n2598_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i310_4_lut_LC_11_11_6 .C_ON=1'b0;
    defparam \tok.i310_4_lut_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i310_4_lut_LC_11_11_6 .LUT_INIT=16'b0001101100001010;
    LogicCell40 \tok.i310_4_lut_LC_11_11_6  (
            .in0(N__31227),
            .in1(N__33467),
            .in2(N__27046),
            .in3(N__27037),
            .lcout(),
            .ltout(\tok.n215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6831_4_lut_LC_11_11_7 .C_ON=1'b0;
    defparam \tok.i6831_4_lut_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6831_4_lut_LC_11_11_7 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \tok.i6831_4_lut_LC_11_11_7  (
            .in0(N__26947),
            .in1(N__26906),
            .in2(N__26878),
            .in3(N__35482),
            .lcout(\tok.n6547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6966_2_lut_LC_11_12_0 .C_ON=1'b0;
    defparam \tok.i6966_2_lut_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6966_2_lut_LC_11_12_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.i6966_2_lut_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__26856),
            .in2(_gnd_net_),
            .in3(N__26838),
            .lcout(),
            .ltout(\tok.n6650_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i337_4_lut_LC_11_12_1 .C_ON=1'b0;
    defparam \tok.i337_4_lut_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i337_4_lut_LC_11_12_1 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \tok.i337_4_lut_LC_11_12_1  (
            .in0(N__35356),
            .in1(N__27609),
            .in2(N__26806),
            .in3(N__26779),
            .lcout(),
            .ltout(\tok.n211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6969_3_lut_LC_11_12_2 .C_ON=1'b0;
    defparam \tok.i6969_3_lut_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6969_3_lut_LC_11_12_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \tok.i6969_3_lut_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__34698),
            .in2(N__26671),
            .in3(N__34053),
            .lcout(\tok.n6641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_105_LC_11_12_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_105_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_105_LC_11_12_3 .LUT_INIT=16'b0001000001010100;
    LogicCell40 \tok.i1_4_lut_adj_105_LC_11_12_3  (
            .in0(N__35357),
            .in1(N__34699),
            .in2(N__26668),
            .in3(N__33233),
            .lcout(),
            .ltout(\tok.n260_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_106_LC_11_12_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_106_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_106_LC_11_12_4 .LUT_INIT=16'b0000000011110010;
    LogicCell40 \tok.i1_4_lut_adj_106_LC_11_12_4  (
            .in0(N__34700),
            .in1(N__37067),
            .in2(N__26644),
            .in3(N__27540),
            .lcout(),
            .ltout(\tok.n266_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_115_LC_11_12_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_115_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_115_LC_11_12_5 .LUT_INIT=16'b1111010111111100;
    LogicCell40 \tok.i1_4_lut_adj_115_LC_11_12_5  (
            .in0(N__27400),
            .in1(N__27619),
            .in2(N__27613),
            .in3(N__36177),
            .lcout(),
            .ltout(\tok.n4_adj_718_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_318_LC_11_12_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_318_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_318_LC_11_12_6 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_318_LC_11_12_6  (
            .in0(N__27610),
            .in1(N__27592),
            .in2(N__27580),
            .in3(N__32078),
            .lcout(\tok.n221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i344_4_lut_LC_11_12_7 .C_ON=1'b0;
    defparam \tok.i344_4_lut_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i344_4_lut_LC_11_12_7 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \tok.i344_4_lut_LC_11_12_7  (
            .in0(N__34052),
            .in1(N__37066),
            .in2(N__27559),
            .in3(N__33232),
            .lcout(\tok.n2637 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i7_LC_11_13_0 .C_ON=1'b0;
    defparam \tok.uart.sender_i7_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i7_LC_11_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.sender_i7_LC_11_13_0  (
            .in0(N__37534),
            .in1(N__27190),
            .in2(_gnd_net_),
            .in3(N__27382),
            .lcout(\tok.uart.sender_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38506),
            .ce(N__27178),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i8_LC_11_13_1 .C_ON=1'b0;
    defparam \tok.uart.sender_i8_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i8_LC_11_13_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i8_LC_11_13_1  (
            .in0(N__27184),
            .in1(N__37535),
            .in2(_gnd_net_),
            .in3(N__30346),
            .lcout(\tok.uart.sender_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38506),
            .ce(N__27178),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i9_LC_11_13_2 .C_ON=1'b0;
    defparam \tok.uart.sender_i9_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i9_LC_11_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.sender_i9_LC_11_13_2  (
            .in0(N__37536),
            .in1(N__37299),
            .in2(_gnd_net_),
            .in3(N__30062),
            .lcout(\tok.uart.sender_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38506),
            .ce(N__27178),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_126_LC_11_13_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_126_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_126_LC_11_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_126_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__34764),
            .in2(_gnd_net_),
            .in3(N__33124),
            .lcout(\tok.n274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_68_LC_11_13_5 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_68_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_68_LC_11_13_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_68_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__32079),
            .in2(_gnd_net_),
            .in3(N__31228),
            .lcout(\tok.n185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_rep_284_2_lut_2_lut_LC_11_13_7 .C_ON=1'b0;
    defparam \tok.i1_rep_284_2_lut_2_lut_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_rep_284_2_lut_2_lut_LC_11_13_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.i1_rep_284_2_lut_2_lut_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__36282),
            .in2(_gnd_net_),
            .in3(N__32080),
            .lcout(\tok.n7410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.reset_I_0_1_lut_LC_12_1_0 .C_ON=1'b0;
    defparam \tok.reset_I_0_1_lut_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \tok.reset_I_0_1_lut_LC_12_1_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \tok.reset_I_0_1_lut_LC_12_1_0  (
            .in0(N__27787),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.reset_N_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i58_LC_12_2_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i58_LC_12_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i58_LC_12_2_3 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \tok.C_stk.tail_i0_i58_LC_12_2_3  (
            .in0(N__27759),
            .in1(N__28835),
            .in2(N__27777),
            .in3(N__28674),
            .lcout(\tok.tail_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38476),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i6_LC_12_3_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i6_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i6_LC_12_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i6_LC_12_3_0  (
            .in0(N__28616),
            .in1(N__27649),
            .in2(_gnd_net_),
            .in3(N__27672),
            .lcout(\tok.C_stk.tail_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38481),
            .ce(N__28910),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i6149_3_lut_LC_12_3_1 .C_ON=1'b0;
    defparam \tok.C_stk.i6149_3_lut_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i6149_3_lut_LC_12_3_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i6149_3_lut_LC_12_3_1  (
            .in0(N__27657),
            .in1(N__28123),
            .in2(_gnd_net_),
            .in3(N__27748),
            .lcout(),
            .ltout(\tok.C_stk.n6233_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i6_LC_12_3_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i6_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i6_LC_12_3_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.C_stk.head_i0_i6_LC_12_3_2  (
            .in0(N__28048),
            .in1(N__27943),
            .in2(N__27718),
            .in3(N__27715),
            .lcout(\tok.c_stk_r_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38481),
            .ce(N__28910),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i14_LC_12_3_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i14_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i14_LC_12_3_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i14_LC_12_3_3  (
            .in0(N__27658),
            .in1(_gnd_net_),
            .in2(N__27640),
            .in3(N__28611),
            .lcout(\tok.tail_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38481),
            .ce(N__28910),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i22_LC_12_3_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i22_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i22_LC_12_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i22_LC_12_3_4  (
            .in0(N__28612),
            .in1(N__27628),
            .in2(_gnd_net_),
            .in3(N__27648),
            .lcout(\tok.C_stk.tail_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38481),
            .ce(N__28910),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i30_LC_12_3_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i30_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i30_LC_12_3_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i30_LC_12_3_5  (
            .in0(N__27636),
            .in1(N__28144),
            .in2(_gnd_net_),
            .in3(N__28613),
            .lcout(\tok.tail_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38481),
            .ce(N__28910),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i38_LC_12_3_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i38_LC_12_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i38_LC_12_3_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i38_LC_12_3_6  (
            .in0(N__28614),
            .in1(N__28135),
            .in2(_gnd_net_),
            .in3(N__27627),
            .lcout(\tok.C_stk.tail_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38481),
            .ce(N__28910),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i46_LC_12_3_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i46_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i46_LC_12_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i46_LC_12_3_7  (
            .in0(N__28158),
            .in1(N__28143),
            .in2(_gnd_net_),
            .in3(N__28615),
            .lcout(\tok.tail_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38481),
            .ce(N__28910),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i7_LC_12_4_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i7_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i7_LC_12_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i7_LC_12_4_0  (
            .in0(N__28665),
            .in1(N__27826),
            .in2(_gnd_net_),
            .in3(N__27853),
            .lcout(\tok.C_stk.tail_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38484),
            .ce(N__28917),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i6143_3_lut_LC_12_4_1 .C_ON=1'b0;
    defparam \tok.C_stk.i6143_3_lut_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i6143_3_lut_LC_12_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.C_stk.i6143_3_lut_LC_12_4_1  (
            .in0(N__27834),
            .in1(N__28118),
            .in2(_gnd_net_),
            .in3(N__28380),
            .lcout(),
            .ltout(\tok.C_stk.n6227_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i7_LC_12_4_2 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i7_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i7_LC_12_4_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.C_stk.head_i0_i7_LC_12_4_2  (
            .in0(N__28052),
            .in1(N__27978),
            .in2(N__27946),
            .in3(N__27942),
            .lcout(\tok.c_stk_r_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38484),
            .ce(N__28917),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i15_LC_12_4_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i15_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i15_LC_12_4_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i15_LC_12_4_3  (
            .in0(N__27835),
            .in1(_gnd_net_),
            .in2(N__27817),
            .in3(N__28660),
            .lcout(\tok.tail_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38484),
            .ce(N__28917),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i23_LC_12_4_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i23_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i23_LC_12_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i23_LC_12_4_4  (
            .in0(N__28661),
            .in1(N__27805),
            .in2(_gnd_net_),
            .in3(N__27825),
            .lcout(\tok.C_stk.tail_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38484),
            .ce(N__28917),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i31_LC_12_4_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i31_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i31_LC_12_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i31_LC_12_4_5  (
            .in0(N__27813),
            .in1(N__27796),
            .in2(_gnd_net_),
            .in3(N__28662),
            .lcout(\tok.tail_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38484),
            .ce(N__28917),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i39_LC_12_4_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i39_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i39_LC_12_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i39_LC_12_4_6  (
            .in0(N__28663),
            .in1(N__28935),
            .in2(_gnd_net_),
            .in3(N__27804),
            .lcout(\tok.C_stk.tail_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38484),
            .ce(N__28917),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i47_LC_12_4_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i47_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i47_LC_12_4_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i47_LC_12_4_7  (
            .in0(N__28776),
            .in1(N__27795),
            .in2(_gnd_net_),
            .in3(N__28664),
            .lcout(\tok.tail_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38484),
            .ce(N__28917),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i63_LC_12_5_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i63_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i63_LC_12_5_1 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \tok.C_stk.tail_i0_i63_LC_12_5_1  (
            .in0(N__28862),
            .in1(N__28494),
            .in2(N__28780),
            .in3(N__28735),
            .lcout(\tok.tail_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1608_3_lut_LC_12_5_2 .C_ON=1'b0;
    defparam \tok.ram.i1608_3_lut_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1608_3_lut_LC_12_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.ram.i1608_3_lut_LC_12_5_2  (
            .in0(N__28472),
            .in1(N__28381),
            .in2(_gnd_net_),
            .in3(N__28339),
            .lcout(\tok.table_wr_data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i1_LC_12_5_3 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i1_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i1_LC_12_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i1_LC_12_5_3  (
            .in0(N__28174),
            .in1(N__37808),
            .in2(_gnd_net_),
            .in3(N__38217),
            .lcout(capture_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i4_LC_12_5_4 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i4_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i4_LC_12_5_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i4_LC_12_5_4  (
            .in0(N__37270),
            .in1(N__37790),
            .in2(_gnd_net_),
            .in3(N__28221),
            .lcout(uart_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i2_LC_12_5_5 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i2_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i2_LC_12_5_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.uart.rx_data_i0_i2_LC_12_5_5  (
            .in0(N__37789),
            .in1(_gnd_net_),
            .in2(N__37288),
            .in3(N__28203),
            .lcout(uart_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i1_LC_12_5_6 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i1_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i1_LC_12_5_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i1_LC_12_5_6  (
            .in0(N__28173),
            .in1(N__37788),
            .in2(_gnd_net_),
            .in3(N__28188),
            .lcout(uart_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i2_LC_12_5_7 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i2_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i2_LC_12_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i2_LC_12_5_7  (
            .in0(N__37284),
            .in1(N__28172),
            .in2(_gnd_net_),
            .in3(N__38218),
            .lcout(capture_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38488),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_87_LC_12_6_0 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_87_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_87_LC_12_6_0 .LUT_INIT=16'b1100100101101100;
    LogicCell40 \tok.i2_4_lut_adj_87_LC_12_6_0  (
            .in0(N__29285),
            .in1(N__29753),
            .in2(N__28981),
            .in3(N__29297),
            .lcout(\tok.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_i1_LC_12_6_1 .C_ON=1'b0;
    defparam \tok.depth_i1_LC_12_6_1 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i1_LC_12_6_1 .LUT_INIT=16'b1001111101100000;
    LogicCell40 \tok.depth_i1_LC_12_6_1  (
            .in0(N__29401),
            .in1(N__29798),
            .in2(N__29359),
            .in3(N__29873),
            .lcout(\tok.depth_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38492),
            .ce(),
            .sr(N__29116));
    defparam \tok.i2_4_lut_4_lut_LC_12_6_2 .C_ON=1'b0;
    defparam \tok.i2_4_lut_4_lut_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_4_lut_LC_12_6_2 .LUT_INIT=16'b1010011001101010;
    LogicCell40 \tok.i2_4_lut_4_lut_LC_12_6_2  (
            .in0(N__29872),
            .in1(N__29355),
            .in2(N__29811),
            .in3(N__29400),
            .lcout(\tok.n52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_72_LC_12_6_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_72_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_72_LC_12_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_adj_72_LC_12_6_3  (
            .in0(N__28971),
            .in1(N__29794),
            .in2(N__29760),
            .in3(N__29870),
            .lcout(\tok.A_stk_delta_1__N_4 ),
            .ltout(\tok.A_stk_delta_1__N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_252_LC_12_6_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_252_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_252_LC_12_6_4 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_252_LC_12_6_4  (
            .in0(N__29871),
            .in1(N__29813),
            .in2(N__29362),
            .in3(N__29354),
            .lcout(\tok.n4_adj_702 ),
            .ltout(\tok.n4_adj_702_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_LC_12_6_5 .C_ON=1'b0;
    defparam \tok.i2_3_lut_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_LC_12_6_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \tok.i2_3_lut_LC_12_6_5  (
            .in0(N__29298),
            .in1(_gnd_net_),
            .in2(N__29323),
            .in3(N__28977),
            .lcout(),
            .ltout(\tok.n51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_LC_12_6_6 .C_ON=1'b0;
    defparam \tok.i3_3_lut_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_LC_12_6_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \tok.i3_3_lut_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__29320),
            .in2(N__29314),
            .in3(N__29311),
            .lcout(\tok.n8_adj_854 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_i3_LC_12_6_7 .C_ON=1'b0;
    defparam \tok.depth_i3_LC_12_6_7 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i3_LC_12_6_7 .LUT_INIT=16'b1011010011010010;
    LogicCell40 \tok.depth_i3_LC_12_6_7  (
            .in0(N__29299),
            .in1(N__29286),
            .in2(N__29761),
            .in3(N__28978),
            .lcout(\tok.depth_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38492),
            .ce(),
            .sr(N__29116));
    defparam \tok.i1_4_lut_adj_151_LC_12_7_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_151_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_151_LC_12_7_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \tok.i1_4_lut_adj_151_LC_12_7_0  (
            .in0(N__29008),
            .in1(N__28999),
            .in2(N__32134),
            .in3(N__34763),
            .lcout(\tok.n215_adj_750 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6129_2_lut_LC_12_7_1 .C_ON=1'b0;
    defparam \tok.i6129_2_lut_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6129_2_lut_LC_12_7_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i6129_2_lut_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__28972),
            .in2(_gnd_net_),
            .in3(N__29875),
            .lcout(\tok.n6213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_4_lut_adj_335_LC_12_7_2 .C_ON=1'b0;
    defparam \tok.i2_3_lut_4_lut_adj_335_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_4_lut_adj_335_LC_12_7_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i2_3_lut_4_lut_adj_335_LC_12_7_2  (
            .in0(N__29874),
            .in1(N__34108),
            .in2(N__29812),
            .in3(N__34760),
            .lcout(\tok.n741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_199_LC_12_7_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_199_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_199_LC_12_7_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_199_LC_12_7_3  (
            .in0(N__34761),
            .in1(_gnd_net_),
            .in2(N__34114),
            .in3(N__37084),
            .lcout(\tok.n806 ),
            .ltout(\tok.n806_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_173_LC_12_7_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_173_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_173_LC_12_7_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \tok.i1_4_lut_adj_173_LC_12_7_4  (
            .in0(N__29802),
            .in1(N__29770),
            .in2(N__29764),
            .in3(N__29758),
            .lcout(\tok.n748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i299_4_lut_adj_119_LC_12_7_5 .C_ON=1'b0;
    defparam \tok.i299_4_lut_adj_119_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i299_4_lut_adj_119_LC_12_7_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.i299_4_lut_adj_119_LC_12_7_5  (
            .in0(N__34762),
            .in1(N__29626),
            .in2(N__29476),
            .in3(N__31310),
            .lcout(),
            .ltout(\tok.n158_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6851_3_lut_4_lut_LC_12_7_6 .C_ON=1'b0;
    defparam \tok.i6851_3_lut_4_lut_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6851_3_lut_4_lut_LC_12_7_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \tok.i6851_3_lut_4_lut_LC_12_7_6  (
            .in0(N__37085),
            .in1(N__32127),
            .in2(N__29461),
            .in3(N__33280),
            .lcout(\tok.n6627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i8_LC_12_7_7 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i8_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i8_LC_12_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.uart.capture_i0_i8_LC_12_7_7  (
            .in0(N__38208),
            .in1(N__37661),
            .in2(_gnd_net_),
            .in3(N__37870),
            .lcout(capture_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38497),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_LC_12_8_0 .C_ON=1'b0;
    defparam \tok.i3_4_lut_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_LC_12_8_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \tok.i3_4_lut_LC_12_8_0  (
            .in0(N__29428),
            .in1(N__37720),
            .in2(N__29422),
            .in3(N__30146),
            .lcout(\tok.uart_stall_N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_373_i9_2_lut_LC_12_8_1 .C_ON=1'b0;
    defparam \tok.T_7__I_0_373_i9_2_lut_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_373_i9_2_lut_LC_12_8_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \tok.T_7__I_0_373_i9_2_lut_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__33244),
            .in2(_gnd_net_),
            .in3(N__30937),
            .lcout(\tok.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_i10_2_lut_LC_12_8_2 .C_ON=1'b0;
    defparam \tok.T_7__I_0_i10_2_lut_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_i10_2_lut_LC_12_8_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.T_7__I_0_i10_2_lut_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__34807),
            .in2(_gnd_net_),
            .in3(N__32113),
            .lcout(\tok.n10 ),
            .ltout(\tok.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7025_2_lut_3_lut_4_lut_LC_12_8_3 .C_ON=1'b0;
    defparam \tok.i7025_2_lut_3_lut_4_lut_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i7025_2_lut_3_lut_4_lut_LC_12_8_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \tok.i7025_2_lut_3_lut_4_lut_LC_12_8_3  (
            .in0(N__30148),
            .in1(N__33248),
            .in2(N__30172),
            .in3(N__30939),
            .lcout(\tok.write_flag ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i4_4_lut_adj_21_LC_12_8_4 .C_ON=1'b0;
    defparam \tok.uart.i4_4_lut_adj_21_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i4_4_lut_adj_21_LC_12_8_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.uart.i4_4_lut_adj_21_LC_12_8_4  (
            .in0(N__30938),
            .in1(N__37721),
            .in2(N__33297),
            .in3(N__30147),
            .lcout(),
            .ltout(\tok.uart.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i7042_3_lut_LC_12_8_5 .C_ON=1'b0;
    defparam \tok.uart.i7042_3_lut_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i7042_3_lut_LC_12_8_5 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \tok.uart.i7042_3_lut_LC_12_8_5  (
            .in0(N__32114),
            .in1(_gnd_net_),
            .in2(N__30094),
            .in3(N__34810),
            .lcout(n23),
            .ltout(n23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i7022_2_lut_3_lut_LC_12_8_6 .C_ON=1'b0;
    defparam \tok.uart.i7022_2_lut_3_lut_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i7022_2_lut_3_lut_LC_12_8_6 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \tok.uart.i7022_2_lut_3_lut_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__37616),
            .in2(N__30091),
            .in3(N__37722),
            .lcout(\tok.uart.n1013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_3_lut_adj_25_LC_12_8_7 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_3_lut_adj_25_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_3_lut_adj_25_LC_12_8_7 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \tok.uart.i1_2_lut_3_lut_adj_25_LC_12_8_7  (
            .in0(N__37723),
            .in1(_gnd_net_),
            .in2(N__37623),
            .in3(N__37500),
            .lcout(\tok.uart.n994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i320_4_lut_4_lut_4_lut_adj_102_LC_12_9_0 .C_ON=1'b0;
    defparam \tok.i320_4_lut_4_lut_4_lut_adj_102_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i320_4_lut_4_lut_4_lut_adj_102_LC_12_9_0 .LUT_INIT=16'b1000010110000000;
    LogicCell40 \tok.i320_4_lut_4_lut_4_lut_adj_102_LC_12_9_0  (
            .in0(N__31305),
            .in1(N__29883),
            .in2(N__32131),
            .in3(N__32378),
            .lcout(),
            .ltout(\tok.n168_adj_710_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6945_4_lut_LC_12_9_1 .C_ON=1'b0;
    defparam \tok.i6945_4_lut_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6945_4_lut_LC_12_9_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i6945_4_lut_LC_12_9_1  (
            .in0(N__32476),
            .in1(N__36364),
            .in2(N__30088),
            .in3(N__30064),
            .lcout(\tok.n6502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i6_LC_12_9_2 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i6_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i6_LC_12_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.uart.rx_data_i0_i6_LC_12_9_2  (
            .in0(N__37791),
            .in1(N__37152),
            .in2(_gnd_net_),
            .in3(N__29884),
            .lcout(uart_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38503),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i7_LC_12_9_3 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i7_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i7_LC_12_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.uart.capture_i0_i7_LC_12_9_3  (
            .in0(N__37151),
            .in1(N__37668),
            .in2(_gnd_net_),
            .in3(N__38184),
            .lcout(capture_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38503),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_105_i15_1_lut_LC_12_9_4 .C_ON=1'b0;
    defparam \tok.inv_105_i15_1_lut_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.inv_105_i15_1_lut_LC_12_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_105_i15_1_lut_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32377),
            .lcout(\tok.n311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_adj_204_LC_12_9_5 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_adj_204_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_adj_204_LC_12_9_5 .LUT_INIT=16'b0101101001001000;
    LogicCell40 \tok.i1_3_lut_4_lut_adj_204_LC_12_9_5  (
            .in0(N__33607),
            .in1(N__32087),
            .in2(N__34112),
            .in3(N__31304),
            .lcout(\tok.n190_adj_797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i320_4_lut_4_lut_4_lut_adj_75_LC_12_9_7 .C_ON=1'b0;
    defparam \tok.i320_4_lut_4_lut_4_lut_adj_75_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i320_4_lut_4_lut_4_lut_adj_75_LC_12_9_7 .LUT_INIT=16'b1100000000100010;
    LogicCell40 \tok.i320_4_lut_4_lut_4_lut_adj_75_LC_12_9_7  (
            .in0(N__32230),
            .in1(N__32091),
            .in2(N__37834),
            .in3(N__31306),
            .lcout(\tok.n168_adj_690 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6949_4_lut_LC_12_10_0 .C_ON=1'b0;
    defparam \tok.i6949_4_lut_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6949_4_lut_LC_12_10_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i6949_4_lut_LC_12_10_0  (
            .in0(N__32470),
            .in1(N__36374),
            .in2(N__30577),
            .in3(N__30314),
            .lcout(),
            .ltout(\tok.n6526_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_180_LC_12_10_1 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_180_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_180_LC_12_10_1 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i308_4_lut_adj_180_LC_12_10_1  (
            .in0(N__30568),
            .in1(N__36269),
            .in2(N__30553),
            .in3(N__33294),
            .lcout(),
            .ltout(\tok.n186_adj_777_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i315_4_lut_adj_190_LC_12_10_2 .C_ON=1'b0;
    defparam \tok.i315_4_lut_adj_190_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i315_4_lut_adj_190_LC_12_10_2 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \tok.i315_4_lut_adj_190_LC_12_10_2  (
            .in0(N__30178),
            .in1(N__35487),
            .in2(N__30550),
            .in3(N__34779),
            .lcout(\tok.n338_adj_787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_61_LC_12_10_4 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_61_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_61_LC_12_10_4 .LUT_INIT=16'b0001000000100000;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_adj_61_LC_12_10_4  (
            .in0(N__30525),
            .in1(N__34095),
            .in2(N__32593),
            .in3(N__37044),
            .lcout(),
            .ltout(\tok.n866_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6793_4_lut_LC_12_10_5 .C_ON=1'b0;
    defparam \tok.i6793_4_lut_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6793_4_lut_LC_12_10_5 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \tok.i6793_4_lut_LC_12_10_5  (
            .in0(N__30313),
            .in1(N__32549),
            .in2(N__30181),
            .in3(N__32581),
            .lcout(\tok.n6520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i271_2_lut_LC_12_11_0 .C_ON=1'b0;
    defparam \tok.i271_2_lut_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i271_2_lut_LC_12_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i271_2_lut_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__35951),
            .in2(_gnd_net_),
            .in3(N__36753),
            .lcout(\tok.n317 ),
            .ltout(\tok.n317_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_98_i8_3_lut_4_lut_LC_12_11_1 .C_ON=1'b0;
    defparam \tok.or_98_i8_3_lut_4_lut_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.or_98_i8_3_lut_4_lut_LC_12_11_1 .LUT_INIT=16'b1111111110101001;
    LogicCell40 \tok.or_98_i8_3_lut_4_lut_LC_12_11_1  (
            .in0(N__34092),
            .in1(N__35483),
            .in2(N__36559),
            .in3(N__36549),
            .lcout(\tok.n205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6934_4_lut_LC_12_11_2 .C_ON=1'b0;
    defparam \tok.i6934_4_lut_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i6934_4_lut_LC_12_11_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i6934_4_lut_LC_12_11_2  (
            .in0(N__36388),
            .in1(N__32472),
            .in2(N__36376),
            .in3(N__37476),
            .lcout(),
            .ltout(\tok.n6478_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i308_4_lut_adj_232_LC_12_11_3 .C_ON=1'b0;
    defparam \tok.i308_4_lut_adj_232_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i308_4_lut_adj_232_LC_12_11_3 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \tok.i308_4_lut_adj_232_LC_12_11_3  (
            .in0(N__35952),
            .in1(N__32386),
            .in2(N__35527),
            .in3(N__33293),
            .lcout(),
            .ltout(\tok.n186_adj_812_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i315_4_lut_adj_241_LC_12_11_4 .C_ON=1'b0;
    defparam \tok.i315_4_lut_adj_241_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i315_4_lut_adj_241_LC_12_11_4 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \tok.i315_4_lut_adj_241_LC_12_11_4  (
            .in0(N__35484),
            .in1(N__32482),
            .in2(N__34849),
            .in3(N__34778),
            .lcout(\tok.n338_adj_819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_290_LC_12_11_5 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_290_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_4_lut_adj_290_LC_12_11_5 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \tok.i1_2_lut_3_lut_4_lut_adj_290_LC_12_11_5  (
            .in0(N__34093),
            .in1(N__33644),
            .in2(N__33483),
            .in3(N__33292),
            .lcout(),
            .ltout(\tok.n863_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6758_4_lut_LC_12_11_6 .C_ON=1'b0;
    defparam \tok.i6758_4_lut_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i6758_4_lut_LC_12_11_6 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \tok.i6758_4_lut_LC_12_11_6  (
            .in0(N__32586),
            .in1(N__32548),
            .in2(N__32485),
            .in3(N__37475),
            .lcout(\tok.n6472 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6760_2_lut_LC_12_11_7 .C_ON=1'b0;
    defparam \tok.i6760_2_lut_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6760_2_lut_LC_12_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i6760_2_lut_LC_12_11_7  (
            .in0(N__32471),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32400),
            .lcout(\tok.n6477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i7_LC_12_12_5 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i7_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i7_LC_12_12_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i7_LC_12_12_5  (
            .in0(N__37669),
            .in1(N__37795),
            .in2(_gnd_net_),
            .in3(N__37641),
            .lcout(uart_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38507),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i10_LC_12_13_3 .C_ON=1'b0;
    defparam \tok.uart.sender_i10_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i10_LC_12_13_3 .LUT_INIT=16'b1111111000110010;
    LogicCell40 \tok.uart.sender_i10_LC_12_13_3  (
            .in0(N__37627),
            .in1(N__37515),
            .in2(N__37303),
            .in3(N__37474),
            .lcout(sender_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38509),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i3_LC_13_5_0 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i3_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i3_LC_13_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i3_LC_13_5_0  (
            .in0(N__37911),
            .in1(N__37283),
            .in2(_gnd_net_),
            .in3(N__38214),
            .lcout(capture_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38493),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_3_lut_LC_13_5_1 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_3_lut_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_3_lut_LC_13_5_1 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \tok.uart.i1_2_lut_3_lut_LC_13_5_1  (
            .in0(N__37787),
            .in1(N__37190),
            .in2(_gnd_net_),
            .in3(N__37242),
            .lcout(\tok.uart.n922 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i4_LC_13_5_4 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i4_LC_13_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i4_LC_13_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i4_LC_13_5_4  (
            .in0(N__37266),
            .in1(N__37910),
            .in2(_gnd_net_),
            .in3(N__38215),
            .lcout(capture_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38493),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i5_LC_13_5_5 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i5_LC_13_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i5_LC_13_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.capture_i0_i5_LC_13_5_5  (
            .in0(N__38216),
            .in1(N__37855),
            .in2(_gnd_net_),
            .in3(N__37265),
            .lcout(capture_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38493),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.valid_54_LC_13_6_0 .C_ON=1'b0;
    defparam \tok.uart.valid_54_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.valid_54_LC_13_6_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \tok.uart.valid_54_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__37191),
            .in2(_gnd_net_),
            .in3(N__37252),
            .lcout(\tok.uart_rx_valid ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38498),
            .ce(N__37171),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i6_LC_13_7_0 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i6_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i6_LC_13_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.uart.capture_i0_i6_LC_13_7_0  (
            .in0(N__38206),
            .in1(N__37847),
            .in2(_gnd_net_),
            .in3(N__37159),
            .lcout(capture_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38501),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i0_LC_13_7_1 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i0_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i0_LC_13_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i0_LC_13_7_1  (
            .in0(N__37815),
            .in1(N__37924),
            .in2(_gnd_net_),
            .in3(N__38205),
            .lcout(capture_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38501),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i2_3_lut_adj_24_LC_13_7_2 .C_ON=1'b0;
    defparam \tok.uart.i2_3_lut_adj_24_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_3_lut_adj_24_LC_13_7_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \tok.uart.i2_3_lut_adj_24_LC_13_7_2  (
            .in0(N__37923),
            .in1(N__37868),
            .in2(_gnd_net_),
            .in3(N__37984),
            .lcout(rx_data_7__N_510),
            .ltout(rx_data_7__N_510_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i3_LC_13_7_3 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i3_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i3_LC_13_7_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \tok.uart.rx_data_i0_i3_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__37915),
            .in2(N__37894),
            .in3(N__37884),
            .lcout(uart_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38501),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i9_LC_13_7_4 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i9_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i9_LC_13_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.capture_i0_i9_LC_13_7_4  (
            .in0(N__38207),
            .in1(N__38010),
            .in2(_gnd_net_),
            .in3(N__37869),
            .lcout(capture_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38501),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i5_LC_13_7_5 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i5_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i5_LC_13_7_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.uart.rx_data_i0_i5_LC_13_7_5  (
            .in0(N__37780),
            .in1(_gnd_net_),
            .in2(N__37854),
            .in3(N__37830),
            .lcout(uart_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38501),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i0_LC_13_7_6 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i0_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i0_LC_13_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i0_LC_13_7_6  (
            .in0(N__37816),
            .in1(N__37779),
            .in2(_gnd_net_),
            .in3(N__37737),
            .lcout(uart_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38501),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i2_4_lut_LC_13_8_0 .C_ON=1'b0;
    defparam \tok.uart.i2_4_lut_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_4_lut_LC_13_8_0 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \tok.uart.i2_4_lut_LC_13_8_0  (
            .in0(N__37707),
            .in1(N__38046),
            .in2(N__37699),
            .in3(N__37681),
            .lcout(\tok.uart_tx_busy ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sentbits_143__i3_LC_13_8_1 .C_ON=1'b0;
    defparam \tok.uart.sentbits_143__i3_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_143__i3_LC_13_8_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \tok.uart.sentbits_143__i3_LC_13_8_1  (
            .in0(N__37684),
            .in1(N__37698),
            .in2(N__38056),
            .in3(N__37708),
            .lcout(\tok.uart.sentbits_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38504),
            .ce(N__38032),
            .sr(N__38020));
    defparam \tok.uart.sentbits_143__i2_LC_13_8_2 .C_ON=1'b0;
    defparam \tok.uart.sentbits_143__i2_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_143__i2_LC_13_8_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \tok.uart.sentbits_143__i2_LC_13_8_2  (
            .in0(N__37697),
            .in1(N__38051),
            .in2(_gnd_net_),
            .in3(N__37683),
            .lcout(\tok.uart.sentbits_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38504),
            .ce(N__38032),
            .sr(N__38020));
    defparam \tok.uart.sentbits_143__i1_LC_13_8_3 .C_ON=1'b0;
    defparam \tok.uart.sentbits_143__i1_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_143__i1_LC_13_8_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \tok.uart.sentbits_143__i1_LC_13_8_3  (
            .in0(N__37682),
            .in1(_gnd_net_),
            .in2(N__38055),
            .in3(_gnd_net_),
            .lcout(\tok.uart.sentbits_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38504),
            .ce(N__38032),
            .sr(N__38020));
    defparam \tok.uart.sentbits_143__i0_LC_13_8_4 .C_ON=1'b0;
    defparam \tok.uart.sentbits_143__i0_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_143__i0_LC_13_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.uart.sentbits_143__i0_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38047),
            .lcout(\tok.uart.sentbits_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38504),
            .ce(N__38032),
            .sr(N__38020));
    defparam \tok.uart.i3_4_lut_LC_13_8_5 .C_ON=1'b0;
    defparam \tok.uart.i3_4_lut_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i3_4_lut_LC_13_8_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \tok.uart.i3_4_lut_LC_13_8_5  (
            .in0(N__38232),
            .in1(N__37962),
            .in2(N__38011),
            .in3(N__37941),
            .lcout(\tok.uart.n809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i3_4_lut_adj_23_LC_13_8_6 .C_ON=1'b0;
    defparam \tok.uart.i3_4_lut_adj_23_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i3_4_lut_adj_23_LC_13_8_6 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \tok.uart.i3_4_lut_adj_23_LC_13_8_6  (
            .in0(N__37940),
            .in1(N__38231),
            .in2(N__37966),
            .in3(N__38629),
            .lcout(\tok.uart.n4977 ),
            .ltout(\tok.uart.n4977_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rxstop_I_0_60_4_lut_LC_13_8_7 .C_ON=1'b0;
    defparam \tok.uart.rxstop_I_0_60_4_lut_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.uart.rxstop_I_0_60_4_lut_LC_13_8_7 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \tok.uart.rxstop_I_0_60_4_lut_LC_13_8_7  (
            .in0(N__38115),
            .in1(N__38128),
            .in2(N__37978),
            .in3(N__38652),
            .lcout(bytephase_5__N_509),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.bytephase__i0_LC_13_9_0 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i0_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i0_LC_13_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i0_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__38076),
            .in2(_gnd_net_),
            .in3(N__37975),
            .lcout(\tok.uart.bytephase_0 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\tok.uart.n4819 ),
            .clk(N__38505),
            .ce(N__38140),
            .sr(N__38158));
    defparam \tok.uart.bytephase__i1_LC_13_9_1 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i1_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i1_LC_13_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i1_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__38653),
            .in2(_gnd_net_),
            .in3(N__37972),
            .lcout(\tok.uart.bytephase_1 ),
            .ltout(),
            .carryin(\tok.uart.n4819 ),
            .carryout(\tok.uart.n4820 ),
            .clk(N__38505),
            .ce(N__38140),
            .sr(N__38158));
    defparam \tok.uart.bytephase__i2_LC_13_9_2 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i2_LC_13_9_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i2_LC_13_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i2_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__38092),
            .in2(_gnd_net_),
            .in3(N__37969),
            .lcout(\tok.uart.bytephase_2 ),
            .ltout(),
            .carryin(\tok.uart.n4820 ),
            .carryout(\tok.uart.n4821 ),
            .clk(N__38505),
            .ce(N__38140),
            .sr(N__38158));
    defparam \tok.uart.bytephase__i3_LC_13_9_3 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i3_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i3_LC_13_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i3_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__37961),
            .in2(_gnd_net_),
            .in3(N__37945),
            .lcout(\tok.uart.bytephase_3 ),
            .ltout(),
            .carryin(\tok.uart.n4821 ),
            .carryout(\tok.uart.n4822 ),
            .clk(N__38505),
            .ce(N__38140),
            .sr(N__38158));
    defparam \tok.uart.bytephase__i4_LC_13_9_4 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i4_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i4_LC_13_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i4_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__37942),
            .in2(_gnd_net_),
            .in3(N__37927),
            .lcout(\tok.uart.bytephase_4 ),
            .ltout(),
            .carryin(\tok.uart.n4822 ),
            .carryout(\tok.uart.n4823 ),
            .clk(N__38505),
            .ce(N__38140),
            .sr(N__38158));
    defparam \tok.uart.bytephase__i5_LC_13_9_5 .C_ON=1'b0;
    defparam \tok.uart.bytephase__i5_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i5_LC_13_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i5_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__38233),
            .in2(_gnd_net_),
            .in3(N__38236),
            .lcout(\tok.uart.bytephase_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38505),
            .ce(N__38140),
            .sr(N__38158));
    defparam \tok.uart.i2_3_lut_LC_13_10_0 .C_ON=1'b0;
    defparam \tok.uart.i2_3_lut_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_3_lut_LC_13_10_0 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \tok.uart.i2_3_lut_LC_13_10_0  (
            .in0(N__38650),
            .in1(_gnd_net_),
            .in2(N__38077),
            .in3(N__38100),
            .lcout(n4928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_LC_13_10_1 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_LC_13_10_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.uart.i1_2_lut_LC_13_10_1  (
            .in0(N__38520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38571),
            .lcout(),
            .ltout(\tok.uart.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i4_4_lut_LC_13_10_2 .C_ON=1'b0;
    defparam \tok.uart.i4_4_lut_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i4_4_lut_LC_13_10_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.uart.i4_4_lut_LC_13_10_2  (
            .in0(N__38605),
            .in1(N__38619),
            .in2(N__38164),
            .in3(N__38134),
            .lcout(n746),
            .ltout(n746_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_13_10_3.C_ON=1'b0;
    defparam i1_2_lut_LC_13_10_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_13_10_3.LUT_INIT=16'b1111111100001111;
    LogicCell40 i1_2_lut_LC_13_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38161),
            .in3(N__38157),
            .lcout(n974),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i6127_3_lut_LC_13_10_4 .C_ON=1'b0;
    defparam \tok.uart.i6127_3_lut_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i6127_3_lut_LC_13_10_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \tok.uart.i6127_3_lut_LC_13_10_4  (
            .in0(N__38586),
            .in1(_gnd_net_),
            .in2(N__38557),
            .in3(N__38538),
            .lcout(\tok.uart.n6211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_adj_22_LC_13_10_5 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_adj_22_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_adj_22_LC_13_10_5 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \tok.uart.i1_2_lut_adj_22_LC_13_10_5  (
            .in0(N__38091),
            .in1(N__38072),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.uart.n2356 ),
            .ltout(\tok.uart.n2356_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rxrst_I_0_3_lut_4_lut_LC_13_10_6 .C_ON=1'b0;
    defparam \tok.uart.rxrst_I_0_3_lut_4_lut_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.rxrst_I_0_3_lut_4_lut_LC_13_10_6 .LUT_INIT=16'b0000010011111111;
    LogicCell40 \tok.uart.rxrst_I_0_3_lut_4_lut_LC_13_10_6  (
            .in0(N__38651),
            .in1(N__38119),
            .in2(N__38104),
            .in3(N__38101),
            .lcout(\tok.uart.rxclkcounter_6__N_476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_3_lut_adj_20_LC_13_10_7 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_3_lut_adj_20_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_3_lut_adj_20_LC_13_10_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.uart.i1_2_lut_3_lut_adj_20_LC_13_10_7  (
            .in0(N__38090),
            .in1(N__38071),
            .in2(_gnd_net_),
            .in3(N__38649),
            .lcout(\tok.uart.n2357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rxclkcounter_144__i0_LC_13_11_0 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_144__i0_LC_13_11_0 .SEQ_MODE=4'b1001;
    defparam \tok.uart.rxclkcounter_144__i0_LC_13_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_144__i0_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__38620),
            .in2(_gnd_net_),
            .in3(N__38608),
            .lcout(\tok.uart.rxclkcounter_0 ),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\tok.uart.n4824 ),
            .clk(N__38508),
            .ce(),
            .sr(N__38251));
    defparam \tok.uart.rxclkcounter_144__i1_LC_13_11_1 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_144__i1_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_144__i1_LC_13_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_144__i1_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__38604),
            .in2(_gnd_net_),
            .in3(N__38590),
            .lcout(\tok.uart.rxclkcounter_1 ),
            .ltout(),
            .carryin(\tok.uart.n4824 ),
            .carryout(\tok.uart.n4825 ),
            .clk(N__38508),
            .ce(),
            .sr(N__38251));
    defparam \tok.uart.rxclkcounter_144__i2_LC_13_11_2 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_144__i2_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_144__i2_LC_13_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_144__i2_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__38587),
            .in2(_gnd_net_),
            .in3(N__38575),
            .lcout(\tok.uart.rxclkcounter_2 ),
            .ltout(),
            .carryin(\tok.uart.n4825 ),
            .carryout(\tok.uart.n4826 ),
            .clk(N__38508),
            .ce(),
            .sr(N__38251));
    defparam \tok.uart.rxclkcounter_144__i3_LC_13_11_3 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_144__i3_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_144__i3_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_144__i3_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__38572),
            .in2(_gnd_net_),
            .in3(N__38560),
            .lcout(\tok.uart.rxclkcounter_3 ),
            .ltout(),
            .carryin(\tok.uart.n4826 ),
            .carryout(\tok.uart.n4827 ),
            .clk(N__38508),
            .ce(),
            .sr(N__38251));
    defparam \tok.uart.rxclkcounter_144__i4_LC_13_11_4 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_144__i4_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_144__i4_LC_13_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_144__i4_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__38556),
            .in2(_gnd_net_),
            .in3(N__38542),
            .lcout(\tok.uart.rxclkcounter_4 ),
            .ltout(),
            .carryin(\tok.uart.n4827 ),
            .carryout(\tok.uart.n4828 ),
            .clk(N__38508),
            .ce(),
            .sr(N__38251));
    defparam \tok.uart.rxclkcounter_144__i5_LC_13_11_5 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_144__i5_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_144__i5_LC_13_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_144__i5_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__38539),
            .in2(_gnd_net_),
            .in3(N__38527),
            .lcout(\tok.uart.rxclkcounter_5 ),
            .ltout(),
            .carryin(\tok.uart.n4828 ),
            .carryout(\tok.uart.n4829 ),
            .clk(N__38508),
            .ce(),
            .sr(N__38251));
    defparam \tok.uart.rxclkcounter_144__i6_LC_13_11_6 .C_ON=1'b0;
    defparam \tok.uart.rxclkcounter_144__i6_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_144__i6_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_144__i6_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__38521),
            .in2(_gnd_net_),
            .in3(N__38524),
            .lcout(\tok.uart.rxclkcounter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38508),
            .ce(),
            .sr(N__38251));
endmodule // top
