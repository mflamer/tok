-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Dec 29 2020 20:58:24

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    tx : out std_logic;
    rx : in std_logic;
    reset : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__30069\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \VCCG0\ : std_logic;
signal \tok.C_stk.n5447_cascade_\ : std_logic;
signal \tok.C_stk.tail_3\ : std_logic;
signal \tok.tail_11\ : std_logic;
signal \tok.C_stk.tail_19\ : std_logic;
signal \tok.tail_27\ : std_logic;
signal \tok.C_stk.tail_35\ : std_logic;
signal \tok.C_stk.n5456_cascade_\ : std_logic;
signal \tok.C_stk.tail_0\ : std_logic;
signal \tok.tail_8\ : std_logic;
signal \tok.C_stk.tail_16\ : std_logic;
signal \tok.tail_24\ : std_logic;
signal \tok.C_stk.tail_32\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \tok.uart.n4827\ : std_logic;
signal \tok.uart.n4828\ : std_logic;
signal \tok.uart.n4829\ : std_logic;
signal \tok.uart.n4830\ : std_logic;
signal \tok.uart.n4831\ : std_logic;
signal \tok.uart.n4832\ : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal \tok.uart.n4814\ : std_logic;
signal \tok.uart.n4815\ : std_logic;
signal \tok.uart.n4816\ : std_logic;
signal \tok.uart.n4817\ : std_logic;
signal \tok.uart.n4818\ : std_logic;
signal \tok.uart.n4819\ : std_logic;
signal \tok.uart.n4820\ : std_logic;
signal \tok.uart.n4821\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \tok.C_stk.n5453_cascade_\ : std_logic;
signal \tok.C_stk.tail_1\ : std_logic;
signal \tok.tail_9\ : std_logic;
signal \tok.C_stk.tail_17\ : std_logic;
signal \tok.tail_25\ : std_logic;
signal \tok.C_stk.tail_33\ : std_logic;
signal \tok.C_stk.n5450_cascade_\ : std_logic;
signal \tok.C_stk.tail_2\ : std_logic;
signal \tok.tail_10\ : std_logic;
signal \tok.C_stk.tail_18\ : std_logic;
signal \tok.tail_26\ : std_logic;
signal \tok.C_stk.tail_34\ : std_logic;
signal \tok.tail_43\ : std_logic;
signal \tok.tail_42\ : std_logic;
signal \tok.tail_41\ : std_logic;
signal \tok.tail_40\ : std_logic;
signal \tok.tail_60\ : std_logic;
signal \tok.tail_51\ : std_logic;
signal \tok.tail_59\ : std_logic;
signal \tok.tail_50\ : std_logic;
signal \tok.tail_58\ : std_logic;
signal \tok.tail_49\ : std_logic;
signal \tok.tail_57\ : std_logic;
signal \tok.tail_48\ : std_logic;
signal \tok.tail_56\ : std_logic;
signal \tok.tail_63\ : std_logic;
signal \tok.C_stk.n5435_cascade_\ : std_logic;
signal \tok.C_stk.tail_7\ : std_logic;
signal \tok.tail_15\ : std_logic;
signal \tok.C_stk.tail_23\ : std_logic;
signal \tok.tail_31\ : std_logic;
signal \tok.C_stk.tail_39\ : std_logic;
signal \tok.tail_55\ : std_logic;
signal \tok.tail_47\ : std_logic;
signal \tok.tail_12\ : std_logic;
signal \tok.C_stk.tail_20\ : std_logic;
signal \tok.tail_28\ : std_logic;
signal \tok.C_stk.tail_36\ : std_logic;
signal \tok.tail_52\ : std_logic;
signal \tok.tail_44\ : std_logic;
signal \bfn_2_2_0_\ : std_logic;
signal \tok.uart.n4822\ : std_logic;
signal \tok.uart.n4823\ : std_logic;
signal \tok.uart.n4824\ : std_logic;
signal \tok.uart.n4825\ : std_logic;
signal \tok.uart.n4826\ : std_logic;
signal \tok.uart.rxclkcounter_5\ : std_logic;
signal \tok.uart.rxclkcounter_3\ : std_logic;
signal \tok.uart.rxclkcounter_2\ : std_logic;
signal \n813_cascade_\ : std_logic;
signal n971 : std_logic;
signal \tok.uart.rxclkcounter_6\ : std_logic;
signal \tok.uart.rxclkcounter_0\ : std_logic;
signal \tok.uart.rxclkcounter_4\ : std_logic;
signal \tok.uart.rxclkcounter_1\ : std_logic;
signal \tok.uart.n12_adj_640\ : std_logic;
signal \tok.uart.sentbits_3\ : std_logic;
signal \tok.uart.txclkcounter_5\ : std_logic;
signal \tok.uart.txclkcounter_2\ : std_logic;
signal \tok.uart.txclkcounter_8\ : std_logic;
signal \tok.uart.txclkcounter_3\ : std_logic;
signal \tok.uart.sentbits_2\ : std_logic;
signal \tok.uart.txclkcounter_4\ : std_logic;
signal \tok.uart.txclkcounter_7\ : std_logic;
signal \tok.uart.txclkcounter_6\ : std_logic;
signal \tok.uart.txclkcounter_0\ : std_logic;
signal \tok.uart.txclkcounter_1\ : std_logic;
signal \tok.uart.n5418_cascade_\ : std_logic;
signal \tok.uart.n12\ : std_logic;
signal \txtick_cascade_\ : std_logic;
signal \tok.tail_61\ : std_logic;
signal \tok.uart.n2_cascade_\ : std_logic;
signal \tok.uart.rxclkcounter_6__N_477\ : std_logic;
signal \tok.uart.bytephase_2\ : std_logic;
signal \tok.uart.n13_cascade_\ : std_logic;
signal \tok.uart.bytephase_4\ : std_logic;
signal \bytephase_5__N_510\ : std_logic;
signal \tok.uart.bytephase_0\ : std_logic;
signal n813 : std_logic;
signal \tok.uart.bytephase_1\ : std_logic;
signal \tok.c_stk_r_2\ : std_logic;
signal \tok.ram.n5585\ : std_logic;
signal \tok.n3_adj_645_cascade_\ : std_logic;
signal \tok.n83\ : std_logic;
signal \tok.n5603\ : std_logic;
signal \tok.n31_adj_795_cascade_\ : std_logic;
signal \tok.n5473\ : std_logic;
signal \tok.C_stk.n5441_cascade_\ : std_logic;
signal \tok.C_stk.tail_5\ : std_logic;
signal \tok.tail_13\ : std_logic;
signal \tok.C_stk.tail_21\ : std_logic;
signal \tok.tail_29\ : std_logic;
signal \tok.C_stk.tail_37\ : std_logic;
signal \tok.tail_53\ : std_logic;
signal \tok.tail_45\ : std_logic;
signal \tok.tc_0\ : std_logic;
signal n92 : std_logic;
signal \n92_cascade_\ : std_logic;
signal \tok.tc_3\ : std_logic;
signal \tok.n13_adj_646\ : std_logic;
signal \n10_cascade_\ : std_logic;
signal \tok.tc_2\ : std_logic;
signal n10 : std_logic;
signal \tok.n36_cascade_\ : std_logic;
signal \tok.n83_adj_842_cascade_\ : std_logic;
signal \tok.ram.n5597_cascade_\ : std_logic;
signal \tok.c_stk_r_0\ : std_logic;
signal \tok.n5583\ : std_logic;
signal \tok.n3_adj_863_cascade_\ : std_logic;
signal \tok.n5_adj_864\ : std_logic;
signal \tok.n83_adj_714_cascade_\ : std_logic;
signal \tok.tc_7\ : std_logic;
signal \tok.ram.n5600_cascade_\ : std_logic;
signal \tok.c_stk_r_7\ : std_logic;
signal \tok.n5511\ : std_logic;
signal \tok.n3_adj_719_cascade_\ : std_logic;
signal \tok.n5_adj_720_cascade_\ : std_logic;
signal n92_adj_869 : std_logic;
signal \n92_adj_869_cascade_\ : std_logic;
signal \tok.n5507\ : std_logic;
signal \tok.C_stk.tail_4\ : std_logic;
signal \tok.tail_62\ : std_logic;
signal \tok.C_stk.n5444\ : std_logic;
signal \tok.tail_54\ : std_logic;
signal \tok.C_stk.tail_38\ : std_logic;
signal \tok.tail_46\ : std_logic;
signal sender_1 : std_logic;
signal tx_c : std_logic;
signal \tok.A_stk.tail_17\ : std_logic;
signal \tok.A_stk.tail_33\ : std_logic;
signal \tok.A_stk.tail_49\ : std_logic;
signal \tok.A_stk.tail_65\ : std_logic;
signal \tok.A_stk.tail_81\ : std_logic;
signal \tok.A_stk.tail_1\ : std_logic;
signal \tok.A_stk_delta_1__N_4_cascade_\ : std_logic;
signal \tok.depth_1_cascade_\ : std_logic;
signal \tok.n37\ : std_logic;
signal \tok.n2585_cascade_\ : std_logic;
signal \tok.n59\ : std_logic;
signal \tok.depth_3\ : std_logic;
signal \tok.n60\ : std_logic;
signal \tok.depth_2\ : std_logic;
signal \tok.n807\ : std_logic;
signal \n23_cascade_\ : std_logic;
signal txtick : std_logic;
signal \tok.uart.sentbits_0\ : std_logic;
signal \tok.uart.sentbits_1\ : std_logic;
signal \tok.uart.n1023\ : std_logic;
signal \tok.uart.n1093\ : std_logic;
signal \tok.n4_adj_707\ : std_logic;
signal \tok.n42\ : std_logic;
signal \tok.n5287\ : std_logic;
signal \tok.n5287_cascade_\ : std_logic;
signal \tok.n7\ : std_logic;
signal \tok.n5312_cascade_\ : std_logic;
signal \tok.n15_adj_817_cascade_\ : std_logic;
signal \tok.n898\ : std_logic;
signal \tok.n898_cascade_\ : std_logic;
signal \tok.uart.n6\ : std_logic;
signal \tok.ram.n5608_cascade_\ : std_logic;
signal \tok.c_stk_r_5\ : std_logic;
signal \tok.n83_adj_678_cascade_\ : std_logic;
signal \tok.n3_adj_683\ : std_logic;
signal \tok.n5483_cascade_\ : std_logic;
signal \tok.n5_adj_684_cascade_\ : std_logic;
signal \n92_adj_868_cascade_\ : std_logic;
signal \tok.tc_5\ : std_logic;
signal n92_adj_868 : std_logic;
signal \tok.table_wr_data_4\ : std_logic;
signal \tok.table_wr_data_15\ : std_logic;
signal \tok.table_wr_data_14\ : std_logic;
signal \tok.table_wr_data_3\ : std_logic;
signal \tok.table_wr_data_2\ : std_logic;
signal \tok.table_wr_data_1\ : std_logic;
signal \tok.table_wr_data_5\ : std_logic;
signal \tok.table_wr_data_7\ : std_logic;
signal \tok.table_wr_data_13\ : std_logic;
signal \tok.table_wr_data_12\ : std_logic;
signal \tok.table_wr_data_11\ : std_logic;
signal \tok.table_wr_data_10\ : std_logic;
signal \tok.table_wr_data_9\ : std_logic;
signal \tok.table_wr_data_8\ : std_logic;
signal \tok.table_wr_data_0\ : std_logic;
signal \tok.n8_adj_790\ : std_logic;
signal \tok.n14_adj_644_cascade_\ : std_logic;
signal \tok.n7_adj_785\ : std_logic;
signal tail_97 : std_logic;
signal tail_113 : std_logic;
signal \tok.n27_adj_828_cascade_\ : std_logic;
signal \tok.n27_adj_831_cascade_\ : std_logic;
signal \tok.n27_adj_833_cascade_\ : std_logic;
signal \tok.n27_adj_825\ : std_logic;
signal \tok.n5285_cascade_\ : std_logic;
signal \tok.n1_adj_715_cascade_\ : std_logic;
signal \tok.n190\ : std_logic;
signal \tok.n890\ : std_logic;
signal \tok.n10_adj_763_cascade_\ : std_logic;
signal \tok.n5338\ : std_logic;
signal \tok.n5340\ : std_logic;
signal \tok.A_stk_delta_1__N_4\ : std_logic;
signal \tok.n61\ : std_logic;
signal \tok.n4_adj_813\ : std_logic;
signal \tok.n13_adj_691_cascade_\ : std_logic;
signal \n10_adj_871_cascade_\ : std_logic;
signal \tok.tc_6\ : std_logic;
signal \tok.ram.n5605_cascade_\ : std_logic;
signal \tok.n3_adj_690\ : std_logic;
signal \tok.n83_adj_687_cascade_\ : std_logic;
signal \tok.n5505\ : std_logic;
signal n10_adj_871 : std_logic;
signal \tok.n83_adj_848_cascade_\ : std_logic;
signal \tok.c_stk_r_1\ : std_logic;
signal \tok.ram.n5594_cascade_\ : std_logic;
signal \tok.n5610\ : std_logic;
signal \tok.n3_cascade_\ : std_logic;
signal \tok.n13_cascade_\ : std_logic;
signal \tok.uart.n5\ : std_logic;
signal \tok.key_rd_10\ : std_logic;
signal \tok.key_rd_12\ : std_logic;
signal \tok.n21_adj_733_cascade_\ : std_logic;
signal \tok.key_rd_7\ : std_logic;
signal \tok.key_rd_2\ : std_logic;
signal \tok.n22_adj_721\ : std_logic;
signal \tok.n23_adj_731\ : std_logic;
signal \tok.n24_adj_651\ : std_logic;
signal \tok.key_rd_14\ : std_logic;
signal \tok.key_rd_15\ : std_logic;
signal \tok.key_rd_9\ : std_logic;
signal \tok.key_rd_11\ : std_logic;
signal tc_0 : std_logic;
signal \tok.tc_plus_1_0\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \tok.tc_plus_1_1\ : std_logic;
signal \tok.n4754\ : std_logic;
signal tc_2 : std_logic;
signal \tok.tc_plus_1_2\ : std_logic;
signal \tok.n4755\ : std_logic;
signal tc_3 : std_logic;
signal \tok.n4756\ : std_logic;
signal \tok.n4757\ : std_logic;
signal tc_5 : std_logic;
signal \tok.tc_plus_1_5\ : std_logic;
signal \tok.n4758\ : std_logic;
signal \tok.n4759\ : std_logic;
signal tc_7 : std_logic;
signal \tok.n4760\ : std_logic;
signal \tok.tc_plus_1_7\ : std_logic;
signal \tok.n9_adj_798\ : std_logic;
signal \tok.n5293\ : std_logic;
signal \tok.n5391\ : std_logic;
signal \tok.n14_adj_688_cascade_\ : std_logic;
signal \tok.n2735_cascade_\ : std_logic;
signal \tok.n1_adj_850_cascade_\ : std_logic;
signal \tok.n26_adj_750\ : std_logic;
signal \tok.n5380\ : std_logic;
signal \tok.n8_adj_805\ : std_logic;
signal \tok.n11_adj_793\ : std_logic;
signal \tok.n5271_cascade_\ : std_logic;
signal \tok.n5318\ : std_logic;
signal \tok.n11_adj_694\ : std_logic;
signal \tok.n15_adj_695\ : std_logic;
signal uart_rx_data_4 : std_logic;
signal \tok.n12_adj_826\ : std_logic;
signal \tok.n11_adj_788\ : std_logic;
signal sender_2 : std_logic;
signal \tok.uart.sender_3\ : std_logic;
signal \tok.uart.sender_4\ : std_logic;
signal \tok.uart.sender_5\ : std_logic;
signal \tok.uart.sender_6\ : std_logic;
signal \tok.uart.sender_7\ : std_logic;
signal sender_9 : std_logic;
signal n23 : std_logic;
signal \tok.uart.sender_8\ : std_logic;
signal \tok.uart.n1017\ : std_logic;
signal \tok.C_stk.n602\ : std_logic;
signal \tok.n241\ : std_logic;
signal \tok.C_stk.n5438_cascade_\ : std_logic;
signal tc_6 : std_logic;
signal \tok.c_stk_r_6\ : std_logic;
signal \tok.C_stk.tail_6\ : std_logic;
signal \tok.n2515\ : std_logic;
signal \tok.tail_14\ : std_logic;
signal \tok.tail_30\ : std_logic;
signal \tok.n29_adj_787\ : std_logic;
signal \tok.C_stk.tail_22\ : std_logic;
signal \tok.C_stk_delta_0\ : std_logic;
signal reset_c : std_logic;
signal \tok.A_stk.tail_16\ : std_logic;
signal \tok.A_stk.tail_32\ : std_logic;
signal \tok.A_stk.tail_48\ : std_logic;
signal \tok.A_stk.tail_64\ : std_logic;
signal tail_112 : std_logic;
signal \tok.A_stk.tail_80\ : std_logic;
signal tail_96 : std_logic;
signal \tok.A_stk.tail_0\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \tok.n4747\ : std_logic;
signal \tok.n4748\ : std_logic;
signal \tok.n4749\ : std_logic;
signal \tok.idx_4\ : std_logic;
signal \tok.n33_adj_819\ : std_logic;
signal \tok.n4750\ : std_logic;
signal \tok.idx_5\ : std_logic;
signal \tok.n33_adj_811\ : std_logic;
signal \tok.n4751\ : std_logic;
signal \tok.idx_6\ : std_logic;
signal \tok.n33_adj_804\ : std_logic;
signal \tok.n4752\ : std_logic;
signal \tok.idx_7\ : std_logic;
signal \tok.n4753\ : std_logic;
signal \tok.n33_adj_801\ : std_logic;
signal \tok.n5_cascade_\ : std_logic;
signal \tok.n5\ : std_logic;
signal \tok.n33\ : std_logic;
signal \tok.n27_cascade_\ : std_logic;
signal \tok.idx_0\ : std_logic;
signal \tok.n83_adj_652_cascade_\ : std_logic;
signal \tok.c_stk_r_3\ : std_logic;
signal \tok.ram.n5580_cascade_\ : std_logic;
signal \tok.n5460\ : std_logic;
signal \tok.n3_adj_659_cascade_\ : std_logic;
signal \tok.tc_plus_1_3\ : std_logic;
signal \tok.n13_adj_660_cascade_\ : std_logic;
signal n92_adj_867 : std_logic;
signal \tok.n17_adj_777\ : std_logic;
signal \tok.n4_adj_778_cascade_\ : std_logic;
signal \tok.n26_adj_760_cascade_\ : std_logic;
signal \tok.n30_adj_761\ : std_logic;
signal \tok.n5587_cascade_\ : std_logic;
signal \tok.key_rd_8\ : std_logic;
signal \tok.n28_adj_755\ : std_logic;
signal \tok.n26_adj_756_cascade_\ : std_logic;
signal \tok.n27_adj_757\ : std_logic;
signal \tok.found_slot_N_145\ : std_logic;
signal \tok.found_slot\ : std_logic;
signal \tok.write_slot\ : std_logic;
signal \tok.key_rd_3\ : std_logic;
signal \tok.key_rd_5\ : std_logic;
signal \tok.n20\ : std_logic;
signal \tok.n18_adj_759\ : std_logic;
signal \tok.key_rd_1\ : std_logic;
signal \tok.key_rd_4\ : std_logic;
signal \tok.n25_adj_758\ : std_logic;
signal \tok.key_rd_0\ : std_logic;
signal \tok.key_rd_6\ : std_logic;
signal \tok.n5590\ : std_logic;
signal uart_rx_data_6 : std_logic;
signal \tok.n6_adj_843\ : std_logic;
signal \tok.n31_adj_844_cascade_\ : std_logic;
signal uart_rx_data_3 : std_logic;
signal capture_4 : std_logic;
signal \tok.tc_plus_1_6\ : std_logic;
signal \tok.table_wr_data_6\ : std_logic;
signal \tok.n10_adj_747\ : std_logic;
signal \tok.n2635\ : std_logic;
signal \tok.n11\ : std_logic;
signal \tok.n2697\ : std_logic;
signal \tok.n15_adj_789\ : std_logic;
signal \tok.n2520\ : std_logic;
signal \tok.n10_adj_803\ : std_logic;
signal \tok.n2520_cascade_\ : std_logic;
signal \tok.n9_adj_802\ : std_logic;
signal \tok.table_rd_3\ : std_logic;
signal \tok.n2661_cascade_\ : std_logic;
signal \tok.n10_adj_845\ : std_logic;
signal \tok.n9_adj_847_cascade_\ : std_logic;
signal \tok.n14_adj_701\ : std_logic;
signal \tok.n5429\ : std_logic;
signal \tok.n5406\ : std_logic;
signal \tok.n5433_cascade_\ : std_logic;
signal \tok.n5272\ : std_logic;
signal \tok.n10_adj_796\ : std_logic;
signal \tok.n14_adj_807\ : std_logic;
signal \tok.n5175\ : std_logic;
signal n10_adj_866 : std_logic;
signal tc_1 : std_logic;
signal \tok.tc_1\ : std_logic;
signal \tok.n2_adj_808\ : std_logic;
signal \tok.n5423\ : std_logic;
signal \tok.n42_adj_751\ : std_logic;
signal capture_9 : std_logic;
signal \tok.n2609\ : std_logic;
signal \tok.n4_adj_712\ : std_logic;
signal \tok.ram.n5577_cascade_\ : std_logic;
signal \tok.n101\ : std_logic;
signal \tok.n3_adj_672\ : std_logic;
signal \tok.n820\ : std_logic;
signal \tok.n5298\ : std_logic;
signal \tok.n13_adj_673_cascade_\ : std_logic;
signal \tok.tc_plus_1_4\ : std_logic;
signal \n10_adj_870_cascade_\ : std_logic;
signal \tok.tc_4\ : std_logic;
signal \stall_\ : std_logic;
signal n10_adj_870 : std_logic;
signal tc_4 : std_logic;
signal \tok.c_stk_r_4\ : std_logic;
signal \tok.n83_adj_665_cascade_\ : std_logic;
signal \tok.n5487\ : std_logic;
signal \tok.A_stk.tail_94\ : std_logic;
signal \tok.A_stk.tail_78\ : std_logic;
signal \tok.A_stk.tail_62\ : std_logic;
signal \tok.A_stk.tail_46\ : std_logic;
signal \tok.A_stk.tail_30\ : std_logic;
signal tail_127 : std_logic;
signal \tok.n33_adj_814\ : std_logic;
signal \tok.n62\ : std_logic;
signal \tok.n1_adj_715\ : std_logic;
signal \tok.depth_0_cascade_\ : std_logic;
signal \tok.n5408\ : std_logic;
signal \tok.n33_adj_816\ : std_logic;
signal \tok.n27_adj_818_cascade_\ : std_logic;
signal \tok.idx_2\ : std_logic;
signal \tok.stall\ : std_logic;
signal \tok.n33_adj_821\ : std_logic;
signal \tok.search_clk\ : std_logic;
signal \tok.n27_adj_822_cascade_\ : std_logic;
signal \tok.idx_3\ : std_logic;
signal \tok.n2699\ : std_logic;
signal \tok.n5282\ : std_logic;
signal \tok.n27_adj_815\ : std_logic;
signal \tok.idx_1\ : std_logic;
signal \rd_15__N_301_cascade_\ : std_logic;
signal \tok.n797\ : std_logic;
signal \tok.n2585\ : std_logic;
signal \A_stk_delta_1_cascade_\ : std_logic;
signal tail_110 : std_logic;
signal tail_126 : std_logic;
signal tail_111 : std_logic;
signal rx_c : std_logic;
signal \tok.uart.n5235\ : std_logic;
signal \tok.uart.bytephase_5\ : std_logic;
signal \tok.uart.bytephase_3\ : std_logic;
signal \tok.uart.n5374\ : std_logic;
signal \tok.key_rd_13\ : std_logic;
signal \tok.n14_adj_647\ : std_logic;
signal capture_0 : std_logic;
signal capture_1 : std_logic;
signal uart_rx_data_0 : std_logic;
signal \tok.n6_adj_794_cascade_\ : std_logic;
signal \tok.table_rd_6\ : std_logic;
signal \tok.n5553_cascade_\ : std_logic;
signal \tok.table_rd_14\ : std_logic;
signal \tok.table_rd_12\ : std_logic;
signal \tok.n14_adj_735_cascade_\ : std_logic;
signal \tok.n6_adj_754\ : std_logic;
signal \tok.table_rd_4\ : std_logic;
signal \tok.n16_adj_851_cascade_\ : std_logic;
signal \tok.n17_adj_853\ : std_logic;
signal \tok.n5562_cascade_\ : std_logic;
signal \tok.n13_adj_852\ : std_logic;
signal \tok.n14_adj_854\ : std_logic;
signal capture_3 : std_logic;
signal \tok.table_rd_0\ : std_logic;
signal \tok.n31\ : std_logic;
signal \tok.n5463_cascade_\ : std_logic;
signal \tok.n2607\ : std_logic;
signal \tok.n14_adj_765\ : std_logic;
signal \tok.table_rd_1\ : std_logic;
signal \tok.n5334_cascade_\ : std_logic;
signal \tok.n5462\ : std_logic;
signal \tok.n5566\ : std_logic;
signal \tok.n5561\ : std_logic;
signal \tok.n9_adj_766\ : std_logic;
signal \tok.n10_adj_643\ : std_logic;
signal \tok.uart_tx_busy\ : std_logic;
signal \tok.n15_adj_655_cascade_\ : std_logic;
signal \tok.uart_stall\ : std_logic;
signal \tok.uart_rx_valid\ : std_logic;
signal \tok.uart.n953\ : std_logic;
signal \tok.n15_adj_667_cascade_\ : std_logic;
signal \tok.table_rd_2\ : std_logic;
signal \tok.n28_adj_771_cascade_\ : std_logic;
signal \tok.n5470\ : std_logic;
signal \tok.n5467_cascade_\ : std_logic;
signal \tok.n34\ : std_logic;
signal \tok.n82_cascade_\ : std_logic;
signal \tok.n878\ : std_logic;
signal \tok.n8_adj_846\ : std_logic;
signal \tok.n41\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \tok.T_1\ : std_logic;
signal \tok.n4761\ : std_logic;
signal \tok.n15_adj_664\ : std_logic;
signal \tok.n4762\ : std_logic;
signal \tok.n82\ : std_logic;
signal \tok.T_3\ : std_logic;
signal \tok.n11_adj_830\ : std_logic;
signal \tok.n4763\ : std_logic;
signal \tok.n212\ : std_logic;
signal \tok.n4764\ : std_logic;
signal \tok.n4765\ : std_logic;
signal \tok.n210\ : std_logic;
signal \tok.n4766\ : std_logic;
signal \tok.n4767\ : std_logic;
signal \tok.n4768\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal tail_121 : std_logic;
signal tail_105 : std_logic;
signal \tok.A_stk.tail_89\ : std_logic;
signal \tok.A_stk.tail_73\ : std_logic;
signal \tok.A_stk.tail_57\ : std_logic;
signal \tok.A_stk.tail_41\ : std_logic;
signal \tok.A_stk.tail_25\ : std_logic;
signal \tok.A_stk.tail_9\ : std_logic;
signal tail_115 : std_logic;
signal tail_99 : std_logic;
signal \tok.A_stk.tail_84\ : std_logic;
signal \tok.A_stk.tail_68\ : std_logic;
signal \tok.A_stk.tail_52\ : std_logic;
signal \tok.A_stk.tail_36\ : std_logic;
signal tail_119 : std_logic;
signal \tok.A_stk.tail_20\ : std_logic;
signal tail_103 : std_logic;
signal \tok.A_stk.tail_71\ : std_logic;
signal \tok.A_stk.tail_87\ : std_logic;
signal tail_120 : std_logic;
signal \tok.A_stk.tail_88\ : std_logic;
signal tail_104 : std_logic;
signal \tok.n9_adj_786\ : std_logic;
signal \tok.table_rd_7\ : std_logic;
signal \tok.n5548_cascade_\ : std_logic;
signal \tok.n285_cascade_\ : std_logic;
signal \tok.n12_adj_824\ : std_logic;
signal \tok.n1_adj_862_cascade_\ : std_logic;
signal \tok.T_6\ : std_logic;
signal \tok.T_4\ : std_logic;
signal \tok.T_5\ : std_logic;
signal \tok.n6_adj_650_cascade_\ : std_logic;
signal \tok.n13_adj_654_cascade_\ : std_logic;
signal \tok.n5547\ : std_logic;
signal \tok.n5546_cascade_\ : std_logic;
signal \tok.n14\ : std_logic;
signal \tok.n17\ : std_logic;
signal \tok.n13_adj_641_cascade_\ : std_logic;
signal \tok.n5552\ : std_logic;
signal \tok.n5551_cascade_\ : std_logic;
signal \tok.n5465\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \tok.n4784\ : std_logic;
signal \tok.n4785\ : std_logic;
signal \tok.n4_adj_806\ : std_logic;
signal \tok.n4786\ : std_logic;
signal \tok.n5564\ : std_logic;
signal \tok.n4787\ : std_logic;
signal \tok.n4788\ : std_logic;
signal \tok.n5554\ : std_logic;
signal \tok.n4789\ : std_logic;
signal \tok.n5549\ : std_logic;
signal \tok.n4790\ : std_logic;
signal \tok.n4791\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \tok.n4792\ : std_logic;
signal \tok.n4793\ : std_logic;
signal \tok.n4794\ : std_logic;
signal \tok.n5_adj_734\ : std_logic;
signal \tok.n4795\ : std_logic;
signal \tok.n4796\ : std_logic;
signal \tok.n5_adj_716\ : std_logic;
signal \tok.n4797\ : std_logic;
signal \tok.n399\ : std_logic;
signal \tok.n4798\ : std_logic;
signal \tok.n8_adj_837\ : std_logic;
signal \tok.n5574\ : std_logic;
signal \tok.n5334\ : std_logic;
signal \tok.n5254\ : std_logic;
signal \tok.n5414_cascade_\ : std_logic;
signal \tok.n8_adj_767\ : std_logic;
signal \tok.n904_cascade_\ : std_logic;
signal \tok.n11_adj_840\ : std_logic;
signal \tok.n5346_cascade_\ : std_logic;
signal \tok.n16_adj_810\ : std_logic;
signal \tok.n14_adj_841_cascade_\ : std_logic;
signal \tok.n5571\ : std_logic;
signal \tok.n5569\ : std_logic;
signal \tok.n45_adj_849\ : std_logic;
signal \tok.n4848\ : std_logic;
signal \tok.table_rd_9\ : std_logic;
signal \tok.n45_cascade_\ : std_logic;
signal \tok.n39\ : std_logic;
signal \tok.n11_adj_680\ : std_logic;
signal \tok.table_rd_10\ : std_logic;
signal \tok.n14_adj_679\ : std_logic;
signal \tok.n45_adj_696\ : std_logic;
signal \tok.n39_adj_697_cascade_\ : std_logic;
signal \tok.n10_adj_700_cascade_\ : std_logic;
signal \tok.n5536\ : std_logic;
signal \tok.n11_adj_730\ : std_logic;
signal \tok.n26_cascade_\ : std_logic;
signal \tok.tc__7__N_134\ : std_logic;
signal \tok.n25_adj_710\ : std_logic;
signal \tok.n28_adj_708\ : std_logic;
signal \tok.n27_adj_709\ : std_logic;
signal \tok.n14_adj_764\ : std_logic;
signal \tok.T_0\ : std_logic;
signal \tok.n10_adj_858\ : std_logic;
signal \tok.table_rd_13\ : std_logic;
signal \tok.n5_adj_732\ : std_logic;
signal \tok.n12_adj_779\ : std_logic;
signal \tok.n14_adj_776_cascade_\ : std_logic;
signal \tok.n13_adj_780\ : std_logic;
signal \tok.n20_adj_784_cascade_\ : std_logic;
signal \tok.n9_adj_781\ : std_logic;
signal \tok.n5_adj_713\ : std_logic;
signal \tok.table_rd_15\ : std_logic;
signal \tok.n16_adj_782\ : std_logic;
signal \tok.n209\ : std_logic;
signal \tok.n14_adj_658\ : std_logic;
signal \tok.n2_adj_775\ : std_logic;
signal tail_118 : std_logic;
signal tail_100 : std_logic;
signal tail_116 : std_logic;
signal tail_114 : std_logic;
signal tail_98 : std_logic;
signal \tok.A_stk.tail_82\ : std_logic;
signal \tok.A_stk.tail_72\ : std_logic;
signal tail_102 : std_logic;
signal \tok.A_stk.tail_70\ : std_logic;
signal \tok.A_stk.tail_86\ : std_logic;
signal \tok.A_stk.tail_55\ : std_logic;
signal \tok.A_stk.tail_39\ : std_logic;
signal \tok.A_stk.tail_83\ : std_logic;
signal \tok.A_stk.tail_4\ : std_logic;
signal \tok.A_stk.tail_6\ : std_logic;
signal \tok.A_stk.tail_54\ : std_logic;
signal \tok.A_stk.tail_22\ : std_logic;
signal \tok.A_stk.tail_38\ : std_logic;
signal \tok.A_stk.tail_23\ : std_logic;
signal \tok.n3_adj_692\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \tok.n4799\ : std_logic;
signal \tok.n4800\ : std_logic;
signal \tok.n22_adj_829\ : std_logic;
signal \tok.n4801\ : std_logic;
signal \tok.n10_adj_827\ : std_logic;
signal \tok.n4802\ : std_logic;
signal \tok.n4803\ : std_logic;
signal \tok.n10_adj_820\ : std_logic;
signal \tok.n4804\ : std_logic;
signal \tok.n10_adj_653\ : std_logic;
signal \tok.n4805\ : std_logic;
signal \tok.n4806\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \tok.n4807\ : std_logic;
signal \tok.n20_adj_663\ : std_logic;
signal \tok.n4808\ : std_logic;
signal \tok.n4809\ : std_logic;
signal \tok.n10_adj_738\ : std_logic;
signal \tok.n4810\ : std_logic;
signal \tok.n4811\ : std_logic;
signal \tok.n10_adj_768\ : std_logic;
signal \tok.n4812\ : std_logic;
signal \tok.write_flag\ : std_logic;
signal \tok.n4813\ : std_logic;
signal \tok.n5516\ : std_logic;
signal \tok.n18_adj_739\ : std_logic;
signal \tok.n12_adj_737_cascade_\ : std_logic;
signal \tok.n1_cascade_\ : std_logic;
signal \tok.n17_adj_656\ : std_logic;
signal \tok.n12\ : std_logic;
signal uart_rx_data_7 : std_logic;
signal \tok.n177\ : std_logic;
signal \tok.n17_adj_812\ : std_logic;
signal \tok.n9_adj_838\ : std_logic;
signal \tok.n23_adj_682\ : std_logic;
signal \tok.n25\ : std_logic;
signal \tok.n4_cascade_\ : std_logic;
signal \tok.n5350\ : std_logic;
signal capture_2 : std_logic;
signal \tok.n9\ : std_logic;
signal \tok.n5342_cascade_\ : std_logic;
signal \tok.n10_adj_686\ : std_logic;
signal \tok.A_low_1\ : std_logic;
signal \tok.n5336\ : std_logic;
signal \tok.table_rd_11\ : std_logic;
signal \tok.n5_adj_726\ : std_logic;
signal \tok.n13_adj_724_cascade_\ : std_logic;
signal \tok.n12_adj_723\ : std_logic;
signal \tok.n5534\ : std_logic;
signal \tok.n16\ : std_logic;
signal \tok.n20_adj_729_cascade_\ : std_logic;
signal \tok.n9_adj_725\ : std_logic;
signal \tok.n5531\ : std_logic;
signal \tok.n2\ : std_logic;
signal \tok.n14_adj_722\ : std_logic;
signal \tok.n20_adj_740\ : std_logic;
signal \tok.n5527_cascade_\ : std_logic;
signal \tok.n5513\ : std_logic;
signal \tok.n5539\ : std_logic;
signal \tok.n5348\ : std_logic;
signal \tok.n13_adj_746_cascade_\ : std_logic;
signal \tok.n12_adj_745\ : std_logic;
signal \tok.n5525\ : std_logic;
signal \tok.n16_adj_749\ : std_logic;
signal \tok.n20_adj_753_cascade_\ : std_logic;
signal \tok.n5522\ : std_logic;
signal \tok.n8\ : std_logic;
signal \tok.n14_adj_744\ : std_logic;
signal \tok.n9_adj_748\ : std_logic;
signal \tok.n2_adj_743\ : std_logic;
signal \tok.n204_cascade_\ : std_logic;
signal \tok.n16_adj_741\ : std_logic;
signal tail_125 : std_logic;
signal tail_109 : std_logic;
signal \tok.A_stk.tail_93\ : std_logic;
signal \tok.A_stk.tail_77\ : std_logic;
signal \tok.A_stk.tail_61\ : std_logic;
signal \tok.A_stk.tail_45\ : std_logic;
signal \tok.A_stk.tail_29\ : std_logic;
signal \tok.A_stk.tail_13\ : std_logic;
signal tail_123 : std_logic;
signal tail_107 : std_logic;
signal \tok.A_stk.tail_91\ : std_logic;
signal tail_124 : std_logic;
signal tail_108 : std_logic;
signal \tok.A_stk.tail_92\ : std_logic;
signal \tok.A_stk.tail_76\ : std_logic;
signal \tok.A_stk.tail_60\ : std_logic;
signal \tok.A_stk.tail_7\ : std_logic;
signal \tok.A_stk.tail_2\ : std_logic;
signal \tok.A_stk.tail_18\ : std_logic;
signal \tok.A_stk.tail_34\ : std_logic;
signal \tok.A_stk.tail_66\ : std_logic;
signal \tok.A_stk.tail_50\ : std_logic;
signal \tok.A_stk.tail_44\ : std_logic;
signal \tok.A_stk.tail_28\ : std_logic;
signal \tok.A_stk.tail_12\ : std_logic;
signal \tok.A_12\ : std_logic;
signal \tok.A_stk.tail_8\ : std_logic;
signal \tok.A_stk.tail_24\ : std_logic;
signal \tok.A_stk.tail_56\ : std_logic;
signal \tok.A_stk.tail_40\ : std_logic;
signal \tok.n22\ : std_logic;
signal \tok.n24\ : std_logic;
signal \tok.n21\ : std_logic;
signal \tok.n30_cascade_\ : std_logic;
signal \tok.n15_adj_671\ : std_logic;
signal \tok.A_low_6\ : std_logic;
signal \tok.n18\ : std_logic;
signal \tok.n17_adj_661_cascade_\ : std_logic;
signal \tok.n19\ : std_logic;
signal \tok.n29\ : std_logic;
signal \tok.A_low_2\ : std_logic;
signal \tok.n22_adj_698\ : std_logic;
signal \tok.n24_adj_703\ : std_logic;
signal \tok.n4_adj_699_cascade_\ : std_logic;
signal \tok.n9_adj_705\ : std_logic;
signal uart_rx_data_1 : std_logic;
signal \tok.n14_adj_662\ : std_logic;
signal \tok.n6_adj_834\ : std_logic;
signal \tok.n23_adj_718\ : std_logic;
signal \tok.n5_adj_835_cascade_\ : std_logic;
signal \tok.n14_adj_644\ : std_logic;
signal \tok.n10_adj_836\ : std_logic;
signal \A_low_7\ : std_logic;
signal \tok.n6_adj_650\ : std_logic;
signal \tok.T_7\ : std_logic;
signal \tok.n11_adj_706\ : std_logic;
signal uart_rx_data_2 : std_logic;
signal \tok.n12_adj_832\ : std_logic;
signal \tok.n6_adj_839_cascade_\ : std_logic;
signal \tok.n11_adj_681\ : std_logic;
signal \tok.n32\ : std_logic;
signal \tok.n15_adj_655\ : std_logic;
signal \tok.A_13\ : std_logic;
signal \tok.n211\ : std_logic;
signal \tok.n184\ : std_logic;
signal capture_5 : std_logic;
signal capture_8 : std_logic;
signal n4858 : std_logic;
signal capture_7 : std_logic;
signal \tok.n17_adj_711\ : std_logic;
signal \tok.S_0\ : std_logic;
signal \tok.n11_adj_809\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \tok.n301\ : std_logic;
signal \tok.S_1\ : std_logic;
signal \tok.n20_adj_799\ : std_logic;
signal \tok.n4769\ : std_logic;
signal \tok.S_2\ : std_logic;
signal \tok.n300\ : std_logic;
signal \tok.n22_adj_797\ : std_logic;
signal \tok.n4770\ : std_logic;
signal \tok.n10_adj_791\ : std_logic;
signal \tok.n4771\ : std_logic;
signal \tok.S_4\ : std_logic;
signal \tok.n6_adj_762\ : std_logic;
signal \tok.n4772\ : std_logic;
signal \tok.n4773\ : std_logic;
signal \tok.S_6\ : std_logic;
signal \tok.n296\ : std_logic;
signal \tok.n6\ : std_logic;
signal \tok.n4774\ : std_logic;
signal \tok.S_7\ : std_logic;
signal \tok.n295\ : std_logic;
signal \tok.n6_adj_657\ : std_logic;
signal \tok.n4775\ : std_logic;
signal \tok.n4776\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \tok.n293\ : std_logic;
signal \tok.n28\ : std_logic;
signal \tok.n4777\ : std_logic;
signal \tok.n8_adj_792\ : std_logic;
signal \tok.n292\ : std_logic;
signal \tok.n27_adj_704\ : std_logic;
signal \tok.n4778\ : std_logic;
signal \tok.n291\ : std_logic;
signal \tok.n6_adj_728\ : std_logic;
signal \tok.n4779\ : std_logic;
signal \tok.n290\ : std_logic;
signal \tok.S_12\ : std_logic;
signal \tok.n6_adj_742\ : std_logic;
signal \tok.n4780\ : std_logic;
signal \tok.n289\ : std_logic;
signal \tok.S_13\ : std_logic;
signal \tok.n6_adj_752\ : std_logic;
signal \tok.n4781\ : std_logic;
signal \tok.n4782\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \tok.n4783\ : std_logic;
signal \tok.n4783_THRU_CRY_0_THRU_CO\ : std_logic;
signal \tok.n400\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \tok.n6_adj_783\ : std_logic;
signal \tok.n287\ : std_logic;
signal \tok.A_15\ : std_logic;
signal \tok.S_15\ : std_logic;
signal \tok.A_stk.tail_15\ : std_logic;
signal \tok.A_stk.tail_31\ : std_logic;
signal \tok.A_stk.tail_47\ : std_logic;
signal \tok.A_stk.tail_95\ : std_logic;
signal \tok.A_stk.tail_63\ : std_logic;
signal \tok.A_stk.tail_79\ : std_logic;
signal \tok.A_stk.tail_74\ : std_logic;
signal \tok.A_stk.tail_58\ : std_logic;
signal \tok.A_stk.tail_42\ : std_logic;
signal \tok.A_stk.tail_26\ : std_logic;
signal \tok.A_stk.tail_10\ : std_logic;
signal tail_117 : std_logic;
signal tail_101 : std_logic;
signal \tok.A_stk.tail_85\ : std_logic;
signal \tok.A_stk.tail_69\ : std_logic;
signal \tok.A_stk.tail_53\ : std_logic;
signal \tok.A_stk.tail_37\ : std_logic;
signal \tok.A_stk.tail_21\ : std_logic;
signal \tok.A_stk.tail_90\ : std_logic;
signal tail_122 : std_logic;
signal tail_106 : std_logic;
signal \tok.n23_adj_642\ : std_logic;
signal \tok.n288\ : std_logic;
signal \tok.A_11\ : std_logic;
signal \tok.A_stk.tail_14\ : std_logic;
signal \tok.S_11\ : std_logic;
signal \tok.A_stk.tail_11\ : std_logic;
signal \tok.A_stk.tail_27\ : std_logic;
signal \tok.A_stk.tail_43\ : std_logic;
signal \tok.A_stk.tail_75\ : std_logic;
signal \tok.A_stk.tail_59\ : std_logic;
signal \tok.n20_adj_648\ : std_logic;
signal \tok.n299\ : std_logic;
signal \tok.n238\ : std_logic;
signal \tok.A_stk.tail_5\ : std_logic;
signal \tok.S_3\ : std_logic;
signal \tok.A_stk.tail_3\ : std_logic;
signal \tok.A_stk.tail_19\ : std_logic;
signal \tok.A_stk.tail_35\ : std_logic;
signal \tok.A_stk.tail_67\ : std_logic;
signal \A_stk_delta_1\ : std_logic;
signal \tok.A_stk.tail_51\ : std_logic;
signal \rd_15__N_301\ : std_logic;
signal \tok.n175\ : std_logic;
signal \tok.n15_adj_770\ : std_logic;
signal \tok.n14_adj_769\ : std_logic;
signal \tok.n13_adj_772_cascade_\ : std_logic;
signal \tok.n5412\ : std_logic;
signal \tok.n22_adj_773_cascade_\ : std_logic;
signal \tok.A_14\ : std_logic;
signal \rx_data_7__N_511\ : std_logic;
signal capture_6 : std_logic;
signal \tok.S_5\ : std_logic;
signal uart_rx_data_5 : std_logic;
signal \tok.n6_adj_717\ : std_logic;
signal \tok.table_rd_5\ : std_logic;
signal \tok.n16_adj_855\ : std_logic;
signal \tok.n5_adj_800\ : std_logic;
signal \tok.n10_adj_823\ : std_logic;
signal \tok.n20_adj_857_cascade_\ : std_logic;
signal \tok.n14_adj_856\ : std_logic;
signal \tok.n5559\ : std_logic;
signal \tok.n3_adj_859\ : std_logic;
signal \tok.n22_adj_861_cascade_\ : std_logic;
signal \tok.n18_adj_860\ : std_logic;
signal \tok.n5556\ : std_logic;
signal \tok.n15\ : std_logic;
signal \tok.n5_adj_669\ : std_logic;
signal \tok.table_rd_8\ : std_logic;
signal \tok.n4908\ : std_logic;
signal \tok.n181\ : std_logic;
signal \tok.n2735\ : std_logic;
signal \tok.n15_adj_670\ : std_logic;
signal \tok.n13_adj_674_cascade_\ : std_logic;
signal \tok.n5416\ : std_logic;
signal \tok.n23\ : std_logic;
signal \tok.n22_adj_676_cascade_\ : std_logic;
signal clk : std_logic;
signal \tok.n995\ : std_logic;
signal \tok.reset_N_2\ : std_logic;
signal \tok.S_8\ : std_logic;
signal \tok.n5544\ : std_logic;
signal \tok.n5542\ : std_logic;
signal \tok.n10_adj_666\ : std_logic;
signal \tok.n15_adj_667\ : std_logic;
signal \tok.n14_adj_668\ : std_logic;
signal \tok.n880\ : std_logic;
signal \tok.A_low_0\ : std_logic;
signal \tok.n904\ : std_logic;
signal \tok.n5372\ : std_logic;
signal \tok.S_9\ : std_logic;
signal \tok.n8_adj_689\ : std_logic;
signal \tok.S_10\ : std_logic;
signal \tok.n8_adj_702\ : std_logic;
signal \tok.n298\ : std_logic;
signal \tok.A_low_5\ : std_logic;
signal \tok.n297\ : std_logic;
signal \tok.T_2\ : std_logic;
signal \tok.n5366\ : std_logic;
signal \tok.A_low_3\ : std_logic;
signal \tok.A_low_4\ : std_logic;
signal \tok.n5396_cascade_\ : std_logic;
signal \tok.n18_adj_677\ : std_logic;
signal \tok.A_8\ : std_logic;
signal \tok.n294\ : std_logic;
signal \tok.n191\ : std_logic;
signal \tok.A_10\ : std_logic;
signal \tok.n2703\ : std_logic;
signal \tok.A_9\ : std_logic;
signal \tok.n202_cascade_\ : std_logic;
signal \tok.n2743\ : std_logic;
signal \tok.n5520\ : std_logic;
signal \tok.S_14\ : std_logic;
signal \tok.n18_adj_774_cascade_\ : std_logic;
signal \tok.n2661\ : std_logic;
signal \tok.n5518\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal rx_wire : std_logic;
signal tx_wire : std_logic;
signal reset_wire : std_logic;
signal \tok.vals.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.vals.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.vals.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.vals.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \tok.vals.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.keys.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.keys.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.keys.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.keys.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \tok.keys.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.ram.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \tok.ram.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.ram.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \tok.ram.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \tok.ram.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    rx_wire <= rx;
    tx <= tx_wire;
    reset_wire <= reset;
    \tok.table_rd_15\ <= \tok.vals.mem1_physical_RDATA_wire\(15);
    \tok.table_rd_14\ <= \tok.vals.mem1_physical_RDATA_wire\(14);
    \tok.table_rd_13\ <= \tok.vals.mem1_physical_RDATA_wire\(13);
    \tok.table_rd_12\ <= \tok.vals.mem1_physical_RDATA_wire\(12);
    \tok.table_rd_11\ <= \tok.vals.mem1_physical_RDATA_wire\(11);
    \tok.table_rd_10\ <= \tok.vals.mem1_physical_RDATA_wire\(10);
    \tok.table_rd_9\ <= \tok.vals.mem1_physical_RDATA_wire\(9);
    \tok.table_rd_8\ <= \tok.vals.mem1_physical_RDATA_wire\(8);
    \tok.table_rd_7\ <= \tok.vals.mem1_physical_RDATA_wire\(7);
    \tok.table_rd_6\ <= \tok.vals.mem1_physical_RDATA_wire\(6);
    \tok.table_rd_5\ <= \tok.vals.mem1_physical_RDATA_wire\(5);
    \tok.table_rd_4\ <= \tok.vals.mem1_physical_RDATA_wire\(4);
    \tok.table_rd_3\ <= \tok.vals.mem1_physical_RDATA_wire\(3);
    \tok.table_rd_2\ <= \tok.vals.mem1_physical_RDATA_wire\(2);
    \tok.table_rd_1\ <= \tok.vals.mem1_physical_RDATA_wire\(1);
    \tok.table_rd_0\ <= \tok.vals.mem1_physical_RDATA_wire\(0);
    \tok.vals.mem1_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__14563\&\N__14638\&\N__14719\&\N__14794\&\N__16786\&\N__16996\&\N__16654\&\N__14872\;
    \tok.vals.mem1_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__14560\&\N__14635\&\N__14710\&\N__14785\&\N__16795\&\N__16993\&\N__16645\&\N__14863\;
    \tok.vals.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \tok.vals.mem1_physical_WDATA_wire\ <= \N__12224\&\N__12212\&\N__12152\&\N__12143\&\N__12266\&\N__12257\&\N__12251\&\N__12245\&\N__12161\&\N__15290\&\N__12170\&\N__12065\&\N__12206\&\N__12194\&\N__12179\&\N__12239\;
    \tok.key_rd_15\ <= \tok.keys.mem0_physical_RDATA_wire\(15);
    \tok.key_rd_14\ <= \tok.keys.mem0_physical_RDATA_wire\(14);
    \tok.key_rd_13\ <= \tok.keys.mem0_physical_RDATA_wire\(13);
    \tok.key_rd_12\ <= \tok.keys.mem0_physical_RDATA_wire\(12);
    \tok.key_rd_11\ <= \tok.keys.mem0_physical_RDATA_wire\(11);
    \tok.key_rd_10\ <= \tok.keys.mem0_physical_RDATA_wire\(10);
    \tok.key_rd_9\ <= \tok.keys.mem0_physical_RDATA_wire\(9);
    \tok.key_rd_8\ <= \tok.keys.mem0_physical_RDATA_wire\(8);
    \tok.key_rd_7\ <= \tok.keys.mem0_physical_RDATA_wire\(7);
    \tok.key_rd_6\ <= \tok.keys.mem0_physical_RDATA_wire\(6);
    \tok.key_rd_5\ <= \tok.keys.mem0_physical_RDATA_wire\(5);
    \tok.key_rd_4\ <= \tok.keys.mem0_physical_RDATA_wire\(4);
    \tok.key_rd_3\ <= \tok.keys.mem0_physical_RDATA_wire\(3);
    \tok.key_rd_2\ <= \tok.keys.mem0_physical_RDATA_wire\(2);
    \tok.key_rd_1\ <= \tok.keys.mem0_physical_RDATA_wire\(1);
    \tok.key_rd_0\ <= \tok.keys.mem0_physical_RDATA_wire\(0);
    \tok.keys.mem0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__14573\&\N__14648\&\N__14726\&\N__14801\&\N__16798\&\N__17006\&\N__16661\&\N__14879\;
    \tok.keys.mem0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__14572\&\N__14647\&\N__14722\&\N__14797\&\N__16802\&\N__17005\&\N__16657\&\N__14875\;
    \tok.keys.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \tok.keys.mem0_physical_WDATA_wire\ <= \N__24863\&\N__25766\&\N__23156\&\N__21633\&\N__25160\&\N__29268\&\N__29080\&\N__29471\&\N__22327\&\N__21895\&\N__27326\&\N__29609\&\N__29730\&\N__22766\&\N__21141\&\N__27780\;
    \tok.T_7\ <= \tok.ram.mem2_physical_RDATA_wire\(14);
    \tok.T_6\ <= \tok.ram.mem2_physical_RDATA_wire\(12);
    \tok.T_5\ <= \tok.ram.mem2_physical_RDATA_wire\(10);
    \tok.T_4\ <= \tok.ram.mem2_physical_RDATA_wire\(8);
    \tok.T_3\ <= \tok.ram.mem2_physical_RDATA_wire\(6);
    \tok.T_2\ <= \tok.ram.mem2_physical_RDATA_wire\(4);
    \tok.T_1\ <= \tok.ram.mem2_physical_RDATA_wire\(2);
    \tok.T_0\ <= \tok.ram.mem2_physical_RDATA_wire\(0);
    \tok.ram.mem2_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__11597\&\N__12524\&\N__12086\&\N__16220\&\N__11366\&\N__11342\&\N__15695\&\N__11390\;
    \tok.ram.mem2_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__23558\&\N__23678\&\N__27221\&\N__23795\&\N__25379\&\N__23939\&\N__24050\&\N__22879\;
    \tok.ram.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \tok.ram.mem2_physical_WDATA_wire\ <= '0'&\N__22328\&'0'&\N__21896\&'0'&\N__27352\&'0'&\N__29600\&'0'&\N__29729\&'0'&\N__22765\&'0'&\N__21140\&'0'&\N__27781\;

    \tok.vals.mem1_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \tok.vals.mem1_physical_RDATA_wire\,
            RADDR => \tok.vals.mem1_physical_RADDR_wire\,
            WADDR => \tok.vals.mem1_physical_WADDR_wire\,
            MASK => \tok.vals.mem1_physical_MASK_wire\,
            WDATA => \tok.vals.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__28504\,
            RE => \N__24254\,
            WCLKE => 'H',
            WCLK => \N__28503\,
            WE => \N__15164\
        );

    \tok.keys.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \tok.keys.mem0_physical_RDATA_wire\,
            RADDR => \tok.keys.mem0_physical_RADDR_wire\,
            WADDR => \tok.keys.mem0_physical_WADDR_wire\,
            MASK => \tok.keys.mem0_physical_MASK_wire\,
            WDATA => \tok.keys.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__28490\,
            RE => \N__24260\,
            WCLKE => 'H',
            WCLK => \N__28491\,
            WE => \N__15163\
        );

    \tok.ram.mem2_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101000100000100000001000001010101000101",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \tok.ram.mem2_physical_RDATA_wire\,
            RADDR => \tok.ram.mem2_physical_RADDR_wire\,
            WADDR => \tok.ram.mem2_physical_WADDR_wire\,
            MASK => \tok.ram.mem2_physical_MASK_wire\,
            WDATA => \tok.ram.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__28515\,
            RE => \N__24247\,
            WCLKE => 'H',
            WCLK => \N__28516\,
            WE => \N__20764\
        );

    \rx_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30069\,
            DIN => \N__30068\,
            DOUT => \N__30067\,
            PACKAGEPIN => rx_wire
        );

    \rx_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30069\,
            PADOUT => \N__30068\,
            PADIN => \N__30067\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => rx_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \tx_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30060\,
            DIN => \N__30059\,
            DOUT => \N__30058\,
            PACKAGEPIN => tx_wire
        );

    \tx_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30060\,
            PADOUT => \N__30059\,
            PADIN => \N__30058\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11621\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \reset_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30051\,
            DIN => \N__30050\,
            DOUT => \N__30049\,
            PACKAGEPIN => reset_wire
        );

    \reset_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30051\,
            PADOUT => \N__30050\,
            PADIN => \N__30049\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => reset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__7478\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30022\
        );

    \I__7477\ : InMux
    port map (
            O => \N__30031\,
            I => \N__30008\
        );

    \I__7476\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30008\
        );

    \I__7475\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30003\
        );

    \I__7474\ : InMux
    port map (
            O => \N__30028\,
            I => \N__30003\
        );

    \I__7473\ : InMux
    port map (
            O => \N__30027\,
            I => \N__29998\
        );

    \I__7472\ : InMux
    port map (
            O => \N__30026\,
            I => \N__29998\
        );

    \I__7471\ : InMux
    port map (
            O => \N__30025\,
            I => \N__29990\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__30022\,
            I => \N__29987\
        );

    \I__7469\ : InMux
    port map (
            O => \N__30021\,
            I => \N__29981\
        );

    \I__7468\ : InMux
    port map (
            O => \N__30020\,
            I => \N__29978\
        );

    \I__7467\ : InMux
    port map (
            O => \N__30019\,
            I => \N__29973\
        );

    \I__7466\ : InMux
    port map (
            O => \N__30018\,
            I => \N__29973\
        );

    \I__7465\ : InMux
    port map (
            O => \N__30017\,
            I => \N__29970\
        );

    \I__7464\ : CascadeMux
    port map (
            O => \N__30016\,
            I => \N__29966\
        );

    \I__7463\ : CascadeMux
    port map (
            O => \N__30015\,
            I => \N__29963\
        );

    \I__7462\ : CascadeMux
    port map (
            O => \N__30014\,
            I => \N__29959\
        );

    \I__7461\ : InMux
    port map (
            O => \N__30013\,
            I => \N__29955\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__30008\,
            I => \N__29948\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__30003\,
            I => \N__29948\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__29998\,
            I => \N__29948\
        );

    \I__7457\ : InMux
    port map (
            O => \N__29997\,
            I => \N__29931\
        );

    \I__7456\ : InMux
    port map (
            O => \N__29996\,
            I => \N__29931\
        );

    \I__7455\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29931\
        );

    \I__7454\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29931\
        );

    \I__7453\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29931\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__29990\,
            I => \N__29928\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__29987\,
            I => \N__29924\
        );

    \I__7450\ : InMux
    port map (
            O => \N__29986\,
            I => \N__29919\
        );

    \I__7449\ : InMux
    port map (
            O => \N__29985\,
            I => \N__29919\
        );

    \I__7448\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29916\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__29981\,
            I => \N__29901\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__29978\,
            I => \N__29901\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__29973\,
            I => \N__29901\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__29970\,
            I => \N__29901\
        );

    \I__7443\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29890\
        );

    \I__7442\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29890\
        );

    \I__7441\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29890\
        );

    \I__7440\ : InMux
    port map (
            O => \N__29962\,
            I => \N__29890\
        );

    \I__7439\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29890\
        );

    \I__7438\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29887\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__29955\,
            I => \N__29882\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__29948\,
            I => \N__29882\
        );

    \I__7435\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29879\
        );

    \I__7434\ : InMux
    port map (
            O => \N__29946\,
            I => \N__29873\
        );

    \I__7433\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29873\
        );

    \I__7432\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29866\
        );

    \I__7431\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29866\
        );

    \I__7430\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29866\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__29931\,
            I => \N__29861\
        );

    \I__7428\ : Span4Mux_h
    port map (
            O => \N__29928\,
            I => \N__29861\
        );

    \I__7427\ : CascadeMux
    port map (
            O => \N__29927\,
            I => \N__29847\
        );

    \I__7426\ : Span4Mux_h
    port map (
            O => \N__29924\,
            I => \N__29844\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__29919\,
            I => \N__29839\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__29916\,
            I => \N__29839\
        );

    \I__7423\ : InMux
    port map (
            O => \N__29915\,
            I => \N__29826\
        );

    \I__7422\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29826\
        );

    \I__7421\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29826\
        );

    \I__7420\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29826\
        );

    \I__7419\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29826\
        );

    \I__7418\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29826\
        );

    \I__7417\ : Span4Mux_s3_v
    port map (
            O => \N__29901\,
            I => \N__29819\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__29890\,
            I => \N__29819\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__29887\,
            I => \N__29819\
        );

    \I__7414\ : Span4Mux_v
    port map (
            O => \N__29882\,
            I => \N__29816\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__29879\,
            I => \N__29813\
        );

    \I__7412\ : InMux
    port map (
            O => \N__29878\,
            I => \N__29810\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__29873\,
            I => \N__29803\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29803\
        );

    \I__7409\ : Span4Mux_v
    port map (
            O => \N__29861\,
            I => \N__29803\
        );

    \I__7408\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29790\
        );

    \I__7407\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29790\
        );

    \I__7406\ : InMux
    port map (
            O => \N__29858\,
            I => \N__29790\
        );

    \I__7405\ : InMux
    port map (
            O => \N__29857\,
            I => \N__29790\
        );

    \I__7404\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29790\
        );

    \I__7403\ : InMux
    port map (
            O => \N__29855\,
            I => \N__29790\
        );

    \I__7402\ : InMux
    port map (
            O => \N__29854\,
            I => \N__29777\
        );

    \I__7401\ : InMux
    port map (
            O => \N__29853\,
            I => \N__29777\
        );

    \I__7400\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29777\
        );

    \I__7399\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29777\
        );

    \I__7398\ : InMux
    port map (
            O => \N__29850\,
            I => \N__29777\
        );

    \I__7397\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29777\
        );

    \I__7396\ : Span4Mux_h
    port map (
            O => \N__29844\,
            I => \N__29770\
        );

    \I__7395\ : Span4Mux_v
    port map (
            O => \N__29839\,
            I => \N__29770\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__29826\,
            I => \N__29770\
        );

    \I__7393\ : Span4Mux_h
    port map (
            O => \N__29819\,
            I => \N__29767\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__29816\,
            I => \tok.T_2\
        );

    \I__7391\ : Odrv4
    port map (
            O => \N__29813\,
            I => \tok.T_2\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__29810\,
            I => \tok.T_2\
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__29803\,
            I => \tok.T_2\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__29790\,
            I => \tok.T_2\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__29777\,
            I => \tok.T_2\
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__29770\,
            I => \tok.T_2\
        );

    \I__7385\ : Odrv4
    port map (
            O => \N__29767\,
            I => \tok.T_2\
        );

    \I__7384\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29747\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__29747\,
            I => \N__29744\
        );

    \I__7382\ : Span4Mux_v
    port map (
            O => \N__29744\,
            I => \N__29741\
        );

    \I__7381\ : Odrv4
    port map (
            O => \N__29741\,
            I => \tok.n5366\
        );

    \I__7380\ : CascadeMux
    port map (
            O => \N__29738\,
            I => \N__29735\
        );

    \I__7379\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29725\
        );

    \I__7378\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29717\
        );

    \I__7377\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29717\
        );

    \I__7376\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29717\
        );

    \I__7375\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29714\
        );

    \I__7374\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29711\
        );

    \I__7373\ : InMux
    port map (
            O => \N__29729\,
            I => \N__29708\
        );

    \I__7372\ : InMux
    port map (
            O => \N__29728\,
            I => \N__29705\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__29725\,
            I => \N__29697\
        );

    \I__7370\ : InMux
    port map (
            O => \N__29724\,
            I => \N__29694\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__29717\,
            I => \N__29691\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__29714\,
            I => \N__29688\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__29711\,
            I => \N__29684\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__29708\,
            I => \N__29681\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29678\
        );

    \I__7364\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29675\
        );

    \I__7363\ : InMux
    port map (
            O => \N__29703\,
            I => \N__29672\
        );

    \I__7362\ : InMux
    port map (
            O => \N__29702\,
            I => \N__29669\
        );

    \I__7361\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29666\
        );

    \I__7360\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29663\
        );

    \I__7359\ : Span4Mux_v
    port map (
            O => \N__29697\,
            I => \N__29658\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__29694\,
            I => \N__29658\
        );

    \I__7357\ : Span4Mux_s2_h
    port map (
            O => \N__29691\,
            I => \N__29655\
        );

    \I__7356\ : Span4Mux_v
    port map (
            O => \N__29688\,
            I => \N__29652\
        );

    \I__7355\ : InMux
    port map (
            O => \N__29687\,
            I => \N__29649\
        );

    \I__7354\ : Span4Mux_h
    port map (
            O => \N__29684\,
            I => \N__29642\
        );

    \I__7353\ : Span4Mux_h
    port map (
            O => \N__29681\,
            I => \N__29642\
        );

    \I__7352\ : Span4Mux_h
    port map (
            O => \N__29678\,
            I => \N__29642\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__29675\,
            I => \N__29637\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__29672\,
            I => \N__29637\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__29669\,
            I => \N__29632\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__29666\,
            I => \N__29632\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__29663\,
            I => \N__29629\
        );

    \I__7346\ : Span4Mux_h
    port map (
            O => \N__29658\,
            I => \N__29624\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__29655\,
            I => \N__29624\
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__29652\,
            I => \tok.A_low_3\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__29649\,
            I => \tok.A_low_3\
        );

    \I__7342\ : Odrv4
    port map (
            O => \N__29642\,
            I => \tok.A_low_3\
        );

    \I__7341\ : Odrv12
    port map (
            O => \N__29637\,
            I => \tok.A_low_3\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__29632\,
            I => \tok.A_low_3\
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__29629\,
            I => \tok.A_low_3\
        );

    \I__7338\ : Odrv4
    port map (
            O => \N__29624\,
            I => \tok.A_low_3\
        );

    \I__7337\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29604\
        );

    \I__7336\ : CascadeMux
    port map (
            O => \N__29608\,
            I => \N__29601\
        );

    \I__7335\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29593\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__29604\,
            I => \N__29590\
        );

    \I__7333\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29587\
        );

    \I__7332\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29582\
        );

    \I__7331\ : InMux
    port map (
            O => \N__29599\,
            I => \N__29579\
        );

    \I__7330\ : InMux
    port map (
            O => \N__29598\,
            I => \N__29576\
        );

    \I__7329\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29573\
        );

    \I__7328\ : InMux
    port map (
            O => \N__29596\,
            I => \N__29570\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__29593\,
            I => \N__29567\
        );

    \I__7326\ : Span4Mux_h
    port map (
            O => \N__29590\,
            I => \N__29559\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__29587\,
            I => \N__29559\
        );

    \I__7324\ : InMux
    port map (
            O => \N__29586\,
            I => \N__29556\
        );

    \I__7323\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29553\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__29582\,
            I => \N__29549\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__29579\,
            I => \N__29546\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__29576\,
            I => \N__29540\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__29573\,
            I => \N__29540\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__29570\,
            I => \N__29537\
        );

    \I__7317\ : Sp12to4
    port map (
            O => \N__29567\,
            I => \N__29534\
        );

    \I__7316\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29527\
        );

    \I__7315\ : InMux
    port map (
            O => \N__29565\,
            I => \N__29527\
        );

    \I__7314\ : InMux
    port map (
            O => \N__29564\,
            I => \N__29527\
        );

    \I__7313\ : Span4Mux_h
    port map (
            O => \N__29559\,
            I => \N__29520\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__29556\,
            I => \N__29520\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__29553\,
            I => \N__29520\
        );

    \I__7310\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29517\
        );

    \I__7309\ : Span4Mux_h
    port map (
            O => \N__29549\,
            I => \N__29514\
        );

    \I__7308\ : Span12Mux_s9_v
    port map (
            O => \N__29546\,
            I => \N__29511\
        );

    \I__7307\ : InMux
    port map (
            O => \N__29545\,
            I => \N__29508\
        );

    \I__7306\ : Span4Mux_h
    port map (
            O => \N__29540\,
            I => \N__29505\
        );

    \I__7305\ : Span12Mux_s4_v
    port map (
            O => \N__29537\,
            I => \N__29498\
        );

    \I__7304\ : Span12Mux_s9_v
    port map (
            O => \N__29534\,
            I => \N__29498\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__29527\,
            I => \N__29498\
        );

    \I__7302\ : Span4Mux_v
    port map (
            O => \N__29520\,
            I => \N__29493\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__29517\,
            I => \N__29493\
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__29514\,
            I => \tok.A_low_4\
        );

    \I__7299\ : Odrv12
    port map (
            O => \N__29511\,
            I => \tok.A_low_4\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__29508\,
            I => \tok.A_low_4\
        );

    \I__7297\ : Odrv4
    port map (
            O => \N__29505\,
            I => \tok.A_low_4\
        );

    \I__7296\ : Odrv12
    port map (
            O => \N__29498\,
            I => \tok.A_low_4\
        );

    \I__7295\ : Odrv4
    port map (
            O => \N__29493\,
            I => \tok.A_low_4\
        );

    \I__7294\ : CascadeMux
    port map (
            O => \N__29480\,
            I => \tok.n5396_cascade_\
        );

    \I__7293\ : InMux
    port map (
            O => \N__29477\,
            I => \N__29474\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__29474\,
            I => \tok.n18_adj_677\
        );

    \I__7291\ : InMux
    port map (
            O => \N__29471\,
            I => \N__29465\
        );

    \I__7290\ : CascadeMux
    port map (
            O => \N__29470\,
            I => \N__29461\
        );

    \I__7289\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29456\
        );

    \I__7288\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29453\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__29465\,
            I => \N__29449\
        );

    \I__7286\ : InMux
    port map (
            O => \N__29464\,
            I => \N__29442\
        );

    \I__7285\ : InMux
    port map (
            O => \N__29461\,
            I => \N__29442\
        );

    \I__7284\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29438\
        );

    \I__7283\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29435\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__29456\,
            I => \N__29430\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__29453\,
            I => \N__29430\
        );

    \I__7280\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29427\
        );

    \I__7279\ : Span4Mux_v
    port map (
            O => \N__29449\,
            I => \N__29424\
        );

    \I__7278\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29421\
        );

    \I__7277\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29418\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29415\
        );

    \I__7275\ : CascadeMux
    port map (
            O => \N__29441\,
            I => \N__29412\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__29438\,
            I => \N__29408\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__29435\,
            I => \N__29402\
        );

    \I__7272\ : Span4Mux_h
    port map (
            O => \N__29430\,
            I => \N__29402\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__29427\,
            I => \N__29399\
        );

    \I__7270\ : Span4Mux_h
    port map (
            O => \N__29424\,
            I => \N__29390\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__29421\,
            I => \N__29390\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__29418\,
            I => \N__29390\
        );

    \I__7267\ : Span4Mux_v
    port map (
            O => \N__29415\,
            I => \N__29390\
        );

    \I__7266\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29385\
        );

    \I__7265\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29385\
        );

    \I__7264\ : Span4Mux_v
    port map (
            O => \N__29408\,
            I => \N__29382\
        );

    \I__7263\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29379\
        );

    \I__7262\ : Span4Mux_h
    port map (
            O => \N__29402\,
            I => \N__29376\
        );

    \I__7261\ : Span4Mux_v
    port map (
            O => \N__29399\,
            I => \N__29371\
        );

    \I__7260\ : Span4Mux_h
    port map (
            O => \N__29390\,
            I => \N__29371\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__29385\,
            I => \tok.A_8\
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__29382\,
            I => \tok.A_8\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__29379\,
            I => \tok.A_8\
        );

    \I__7256\ : Odrv4
    port map (
            O => \N__29376\,
            I => \tok.A_8\
        );

    \I__7255\ : Odrv4
    port map (
            O => \N__29371\,
            I => \tok.A_8\
        );

    \I__7254\ : InMux
    port map (
            O => \N__29360\,
            I => \N__29357\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__29357\,
            I => \tok.n294\
        );

    \I__7252\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29350\
        );

    \I__7251\ : InMux
    port map (
            O => \N__29353\,
            I => \N__29346\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__29350\,
            I => \N__29340\
        );

    \I__7249\ : InMux
    port map (
            O => \N__29349\,
            I => \N__29337\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__29346\,
            I => \N__29334\
        );

    \I__7247\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29329\
        );

    \I__7246\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29329\
        );

    \I__7245\ : InMux
    port map (
            O => \N__29343\,
            I => \N__29326\
        );

    \I__7244\ : Span4Mux_v
    port map (
            O => \N__29340\,
            I => \N__29323\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__29337\,
            I => \N__29320\
        );

    \I__7242\ : Span4Mux_s2_h
    port map (
            O => \N__29334\,
            I => \N__29314\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__29329\,
            I => \N__29314\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__29326\,
            I => \N__29311\
        );

    \I__7239\ : Span4Mux_h
    port map (
            O => \N__29323\,
            I => \N__29305\
        );

    \I__7238\ : Span4Mux_v
    port map (
            O => \N__29320\,
            I => \N__29305\
        );

    \I__7237\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29302\
        );

    \I__7236\ : Span4Mux_h
    port map (
            O => \N__29314\,
            I => \N__29299\
        );

    \I__7235\ : Span4Mux_h
    port map (
            O => \N__29311\,
            I => \N__29296\
        );

    \I__7234\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29293\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__29305\,
            I => \tok.n191\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__29302\,
            I => \tok.n191\
        );

    \I__7231\ : Odrv4
    port map (
            O => \N__29299\,
            I => \tok.n191\
        );

    \I__7230\ : Odrv4
    port map (
            O => \N__29296\,
            I => \tok.n191\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__29293\,
            I => \tok.n191\
        );

    \I__7228\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29279\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29275\
        );

    \I__7226\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29272\
        );

    \I__7225\ : Span4Mux_s3_v
    port map (
            O => \N__29275\,
            I => \N__29263\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__29272\,
            I => \N__29260\
        );

    \I__7223\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29257\
        );

    \I__7222\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29254\
        );

    \I__7221\ : InMux
    port map (
            O => \N__29269\,
            I => \N__29250\
        );

    \I__7220\ : InMux
    port map (
            O => \N__29268\,
            I => \N__29246\
        );

    \I__7219\ : InMux
    port map (
            O => \N__29267\,
            I => \N__29241\
        );

    \I__7218\ : InMux
    port map (
            O => \N__29266\,
            I => \N__29241\
        );

    \I__7217\ : Span4Mux_v
    port map (
            O => \N__29263\,
            I => \N__29233\
        );

    \I__7216\ : Span4Mux_v
    port map (
            O => \N__29260\,
            I => \N__29233\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__29257\,
            I => \N__29233\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__29254\,
            I => \N__29230\
        );

    \I__7213\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29227\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__29250\,
            I => \N__29224\
        );

    \I__7211\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29221\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__29246\,
            I => \N__29216\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__29241\,
            I => \N__29216\
        );

    \I__7208\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29212\
        );

    \I__7207\ : Span4Mux_h
    port map (
            O => \N__29233\,
            I => \N__29209\
        );

    \I__7206\ : Span4Mux_v
    port map (
            O => \N__29230\,
            I => \N__29204\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__29227\,
            I => \N__29204\
        );

    \I__7204\ : Span4Mux_h
    port map (
            O => \N__29224\,
            I => \N__29199\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__29221\,
            I => \N__29199\
        );

    \I__7202\ : Span4Mux_h
    port map (
            O => \N__29216\,
            I => \N__29196\
        );

    \I__7201\ : InMux
    port map (
            O => \N__29215\,
            I => \N__29193\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__29212\,
            I => \tok.A_10\
        );

    \I__7199\ : Odrv4
    port map (
            O => \N__29209\,
            I => \tok.A_10\
        );

    \I__7198\ : Odrv4
    port map (
            O => \N__29204\,
            I => \tok.A_10\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__29199\,
            I => \tok.A_10\
        );

    \I__7196\ : Odrv4
    port map (
            O => \N__29196\,
            I => \tok.A_10\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__29193\,
            I => \tok.A_10\
        );

    \I__7194\ : InMux
    port map (
            O => \N__29180\,
            I => \N__29175\
        );

    \I__7193\ : InMux
    port map (
            O => \N__29179\,
            I => \N__29172\
        );

    \I__7192\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29168\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__29175\,
            I => \N__29164\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__29172\,
            I => \N__29161\
        );

    \I__7189\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29157\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__29168\,
            I => \N__29154\
        );

    \I__7187\ : InMux
    port map (
            O => \N__29167\,
            I => \N__29150\
        );

    \I__7186\ : Span4Mux_s1_h
    port map (
            O => \N__29164\,
            I => \N__29143\
        );

    \I__7185\ : Span4Mux_v
    port map (
            O => \N__29161\,
            I => \N__29143\
        );

    \I__7184\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29140\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__29157\,
            I => \N__29135\
        );

    \I__7182\ : Span4Mux_s3_h
    port map (
            O => \N__29154\,
            I => \N__29132\
        );

    \I__7181\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29129\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__29150\,
            I => \N__29126\
        );

    \I__7179\ : InMux
    port map (
            O => \N__29149\,
            I => \N__29123\
        );

    \I__7178\ : InMux
    port map (
            O => \N__29148\,
            I => \N__29120\
        );

    \I__7177\ : Span4Mux_h
    port map (
            O => \N__29143\,
            I => \N__29114\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__29140\,
            I => \N__29114\
        );

    \I__7175\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29109\
        );

    \I__7174\ : InMux
    port map (
            O => \N__29138\,
            I => \N__29109\
        );

    \I__7173\ : Span4Mux_s2_v
    port map (
            O => \N__29135\,
            I => \N__29102\
        );

    \I__7172\ : Span4Mux_v
    port map (
            O => \N__29132\,
            I => \N__29102\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__29129\,
            I => \N__29102\
        );

    \I__7170\ : Sp12to4
    port map (
            O => \N__29126\,
            I => \N__29095\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__29123\,
            I => \N__29095\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__29120\,
            I => \N__29095\
        );

    \I__7167\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29092\
        );

    \I__7166\ : Odrv4
    port map (
            O => \N__29114\,
            I => \tok.n2703\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__29109\,
            I => \tok.n2703\
        );

    \I__7164\ : Odrv4
    port map (
            O => \N__29102\,
            I => \tok.n2703\
        );

    \I__7163\ : Odrv12
    port map (
            O => \N__29095\,
            I => \tok.n2703\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__29092\,
            I => \tok.n2703\
        );

    \I__7161\ : InMux
    port map (
            O => \N__29081\,
            I => \N__29076\
        );

    \I__7160\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29071\
        );

    \I__7159\ : InMux
    port map (
            O => \N__29079\,
            I => \N__29067\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__29076\,
            I => \N__29062\
        );

    \I__7157\ : InMux
    port map (
            O => \N__29075\,
            I => \N__29056\
        );

    \I__7156\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29056\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__29071\,
            I => \N__29053\
        );

    \I__7154\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29050\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__29067\,
            I => \N__29047\
        );

    \I__7152\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29044\
        );

    \I__7151\ : CascadeMux
    port map (
            O => \N__29065\,
            I => \N__29041\
        );

    \I__7150\ : Span4Mux_s2_v
    port map (
            O => \N__29062\,
            I => \N__29035\
        );

    \I__7149\ : InMux
    port map (
            O => \N__29061\,
            I => \N__29032\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__29056\,
            I => \N__29029\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__29053\,
            I => \N__29024\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__29050\,
            I => \N__29024\
        );

    \I__7145\ : Sp12to4
    port map (
            O => \N__29047\,
            I => \N__29021\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__29044\,
            I => \N__29018\
        );

    \I__7143\ : InMux
    port map (
            O => \N__29041\,
            I => \N__29015\
        );

    \I__7142\ : InMux
    port map (
            O => \N__29040\,
            I => \N__29012\
        );

    \I__7141\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29009\
        );

    \I__7140\ : InMux
    port map (
            O => \N__29038\,
            I => \N__29006\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__29035\,
            I => \N__28997\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__29032\,
            I => \N__28997\
        );

    \I__7137\ : Span4Mux_h
    port map (
            O => \N__29029\,
            I => \N__28997\
        );

    \I__7136\ : Span4Mux_h
    port map (
            O => \N__29024\,
            I => \N__28997\
        );

    \I__7135\ : Odrv12
    port map (
            O => \N__29021\,
            I => \tok.A_9\
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__29018\,
            I => \tok.A_9\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__29015\,
            I => \tok.A_9\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__29012\,
            I => \tok.A_9\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__29009\,
            I => \tok.A_9\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__29006\,
            I => \tok.A_9\
        );

    \I__7129\ : Odrv4
    port map (
            O => \N__28997\,
            I => \tok.A_9\
        );

    \I__7128\ : CascadeMux
    port map (
            O => \N__28982\,
            I => \tok.n202_cascade_\
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__28979\,
            I => \N__28974\
        );

    \I__7126\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28967\
        );

    \I__7125\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28964\
        );

    \I__7124\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28957\
        );

    \I__7123\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28957\
        );

    \I__7122\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28957\
        );

    \I__7121\ : InMux
    port map (
            O => \N__28971\,
            I => \N__28954\
        );

    \I__7120\ : InMux
    port map (
            O => \N__28970\,
            I => \N__28951\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__28967\,
            I => \N__28946\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__28964\,
            I => \N__28943\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__28957\,
            I => \N__28940\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__28954\,
            I => \N__28930\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28930\
        );

    \I__7114\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28925\
        );

    \I__7113\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28925\
        );

    \I__7112\ : Span4Mux_v
    port map (
            O => \N__28946\,
            I => \N__28922\
        );

    \I__7111\ : Span4Mux_v
    port map (
            O => \N__28943\,
            I => \N__28917\
        );

    \I__7110\ : Span4Mux_v
    port map (
            O => \N__28940\,
            I => \N__28917\
        );

    \I__7109\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28914\
        );

    \I__7108\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28905\
        );

    \I__7107\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28905\
        );

    \I__7106\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28905\
        );

    \I__7105\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28905\
        );

    \I__7104\ : Span4Mux_h
    port map (
            O => \N__28930\,
            I => \N__28901\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__28925\,
            I => \N__28898\
        );

    \I__7102\ : Span4Mux_v
    port map (
            O => \N__28922\,
            I => \N__28893\
        );

    \I__7101\ : Span4Mux_h
    port map (
            O => \N__28917\,
            I => \N__28893\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__28914\,
            I => \N__28888\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__28905\,
            I => \N__28888\
        );

    \I__7098\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28885\
        );

    \I__7097\ : Odrv4
    port map (
            O => \N__28901\,
            I => \tok.n2743\
        );

    \I__7096\ : Odrv4
    port map (
            O => \N__28898\,
            I => \tok.n2743\
        );

    \I__7095\ : Odrv4
    port map (
            O => \N__28893\,
            I => \tok.n2743\
        );

    \I__7094\ : Odrv12
    port map (
            O => \N__28888\,
            I => \tok.n2743\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__28885\,
            I => \tok.n2743\
        );

    \I__7092\ : InMux
    port map (
            O => \N__28874\,
            I => \N__28871\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__28871\,
            I => \tok.n5520\
        );

    \I__7090\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28863\
        );

    \I__7089\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28860\
        );

    \I__7088\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28854\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__28863\,
            I => \N__28851\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__28860\,
            I => \N__28847\
        );

    \I__7085\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28844\
        );

    \I__7084\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28841\
        );

    \I__7083\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28838\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__28854\,
            I => \N__28834\
        );

    \I__7081\ : Span4Mux_s3_v
    port map (
            O => \N__28851\,
            I => \N__28831\
        );

    \I__7080\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28828\
        );

    \I__7079\ : Span4Mux_h
    port map (
            O => \N__28847\,
            I => \N__28823\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__28844\,
            I => \N__28823\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__28841\,
            I => \N__28818\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__28838\,
            I => \N__28818\
        );

    \I__7075\ : CascadeMux
    port map (
            O => \N__28837\,
            I => \N__28815\
        );

    \I__7074\ : Span4Mux_v
    port map (
            O => \N__28834\,
            I => \N__28812\
        );

    \I__7073\ : Span4Mux_h
    port map (
            O => \N__28831\,
            I => \N__28803\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__28828\,
            I => \N__28803\
        );

    \I__7071\ : Span4Mux_h
    port map (
            O => \N__28823\,
            I => \N__28803\
        );

    \I__7070\ : Span4Mux_v
    port map (
            O => \N__28818\,
            I => \N__28803\
        );

    \I__7069\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28800\
        );

    \I__7068\ : Odrv4
    port map (
            O => \N__28812\,
            I => \tok.S_14\
        );

    \I__7067\ : Odrv4
    port map (
            O => \N__28803\,
            I => \tok.S_14\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__28800\,
            I => \tok.S_14\
        );

    \I__7065\ : CascadeMux
    port map (
            O => \N__28793\,
            I => \tok.n18_adj_774_cascade_\
        );

    \I__7064\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28778\
        );

    \I__7063\ : CascadeMux
    port map (
            O => \N__28789\,
            I => \N__28774\
        );

    \I__7062\ : InMux
    port map (
            O => \N__28788\,
            I => \N__28771\
        );

    \I__7061\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28768\
        );

    \I__7060\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28763\
        );

    \I__7059\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28763\
        );

    \I__7058\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28759\
        );

    \I__7057\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28755\
        );

    \I__7056\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28752\
        );

    \I__7055\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28748\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__28778\,
            I => \N__28745\
        );

    \I__7053\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28742\
        );

    \I__7052\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28739\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__28771\,
            I => \N__28736\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__28768\,
            I => \N__28731\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__28763\,
            I => \N__28731\
        );

    \I__7048\ : CascadeMux
    port map (
            O => \N__28762\,
            I => \N__28727\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__28759\,
            I => \N__28724\
        );

    \I__7046\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28721\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__28755\,
            I => \N__28716\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28716\
        );

    \I__7043\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28713\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__28748\,
            I => \N__28704\
        );

    \I__7041\ : Span4Mux_h
    port map (
            O => \N__28745\,
            I => \N__28704\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__28742\,
            I => \N__28704\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__28739\,
            I => \N__28704\
        );

    \I__7038\ : Span4Mux_v
    port map (
            O => \N__28736\,
            I => \N__28699\
        );

    \I__7037\ : Span4Mux_v
    port map (
            O => \N__28731\,
            I => \N__28699\
        );

    \I__7036\ : InMux
    port map (
            O => \N__28730\,
            I => \N__28696\
        );

    \I__7035\ : InMux
    port map (
            O => \N__28727\,
            I => \N__28693\
        );

    \I__7034\ : Span4Mux_s3_h
    port map (
            O => \N__28724\,
            I => \N__28686\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__28721\,
            I => \N__28686\
        );

    \I__7032\ : Span4Mux_v
    port map (
            O => \N__28716\,
            I => \N__28686\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__28713\,
            I => \N__28683\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__28704\,
            I => \N__28678\
        );

    \I__7029\ : Span4Mux_h
    port map (
            O => \N__28699\,
            I => \N__28678\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__28696\,
            I => \tok.n2661\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__28693\,
            I => \tok.n2661\
        );

    \I__7026\ : Odrv4
    port map (
            O => \N__28686\,
            I => \tok.n2661\
        );

    \I__7025\ : Odrv12
    port map (
            O => \N__28683\,
            I => \tok.n2661\
        );

    \I__7024\ : Odrv4
    port map (
            O => \N__28678\,
            I => \tok.n2661\
        );

    \I__7023\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28664\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__28664\,
            I => \N__28661\
        );

    \I__7021\ : Odrv12
    port map (
            O => \N__28661\,
            I => \tok.n5518\
        );

    \I__7020\ : CascadeMux
    port map (
            O => \N__28658\,
            I => \N__28654\
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__28657\,
            I => \N__28649\
        );

    \I__7018\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28639\
        );

    \I__7017\ : InMux
    port map (
            O => \N__28653\,
            I => \N__28639\
        );

    \I__7016\ : InMux
    port map (
            O => \N__28652\,
            I => \N__28639\
        );

    \I__7015\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28639\
        );

    \I__7014\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28633\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__28639\,
            I => \N__28630\
        );

    \I__7012\ : CascadeMux
    port map (
            O => \N__28638\,
            I => \N__28627\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__28637\,
            I => \N__28621\
        );

    \I__7010\ : CascadeMux
    port map (
            O => \N__28636\,
            I => \N__28615\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__28633\,
            I => \N__28610\
        );

    \I__7008\ : Span4Mux_h
    port map (
            O => \N__28630\,
            I => \N__28610\
        );

    \I__7007\ : InMux
    port map (
            O => \N__28627\,
            I => \N__28605\
        );

    \I__7006\ : InMux
    port map (
            O => \N__28626\,
            I => \N__28605\
        );

    \I__7005\ : InMux
    port map (
            O => \N__28625\,
            I => \N__28590\
        );

    \I__7004\ : InMux
    port map (
            O => \N__28624\,
            I => \N__28590\
        );

    \I__7003\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28590\
        );

    \I__7002\ : InMux
    port map (
            O => \N__28620\,
            I => \N__28590\
        );

    \I__7001\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28590\
        );

    \I__7000\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28590\
        );

    \I__6999\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28590\
        );

    \I__6998\ : Span4Mux_v
    port map (
            O => \N__28610\,
            I => \N__28583\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__28605\,
            I => \N__28583\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__28590\,
            I => \N__28579\
        );

    \I__6995\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28574\
        );

    \I__6994\ : InMux
    port map (
            O => \N__28588\,
            I => \N__28574\
        );

    \I__6993\ : Span4Mux_v
    port map (
            O => \N__28583\,
            I => \N__28571\
        );

    \I__6992\ : InMux
    port map (
            O => \N__28582\,
            I => \N__28568\
        );

    \I__6991\ : Span4Mux_v
    port map (
            O => \N__28579\,
            I => \N__28563\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__28574\,
            I => \N__28563\
        );

    \I__6989\ : Span4Mux_h
    port map (
            O => \N__28571\,
            I => \N__28558\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__28568\,
            I => \N__28558\
        );

    \I__6987\ : Span4Mux_v
    port map (
            O => \N__28563\,
            I => \N__28555\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__28558\,
            I => \N__28552\
        );

    \I__6985\ : Odrv4
    port map (
            O => \N__28555\,
            I => \tok.n23\
        );

    \I__6984\ : Odrv4
    port map (
            O => \N__28552\,
            I => \tok.n23\
        );

    \I__6983\ : CascadeMux
    port map (
            O => \N__28547\,
            I => \tok.n22_adj_676_cascade_\
        );

    \I__6982\ : ClkMux
    port map (
            O => \N__28544\,
            I => \N__28307\
        );

    \I__6981\ : ClkMux
    port map (
            O => \N__28543\,
            I => \N__28307\
        );

    \I__6980\ : ClkMux
    port map (
            O => \N__28542\,
            I => \N__28307\
        );

    \I__6979\ : ClkMux
    port map (
            O => \N__28541\,
            I => \N__28307\
        );

    \I__6978\ : ClkMux
    port map (
            O => \N__28540\,
            I => \N__28307\
        );

    \I__6977\ : ClkMux
    port map (
            O => \N__28539\,
            I => \N__28307\
        );

    \I__6976\ : ClkMux
    port map (
            O => \N__28538\,
            I => \N__28307\
        );

    \I__6975\ : ClkMux
    port map (
            O => \N__28537\,
            I => \N__28307\
        );

    \I__6974\ : ClkMux
    port map (
            O => \N__28536\,
            I => \N__28307\
        );

    \I__6973\ : ClkMux
    port map (
            O => \N__28535\,
            I => \N__28307\
        );

    \I__6972\ : ClkMux
    port map (
            O => \N__28534\,
            I => \N__28307\
        );

    \I__6971\ : ClkMux
    port map (
            O => \N__28533\,
            I => \N__28307\
        );

    \I__6970\ : ClkMux
    port map (
            O => \N__28532\,
            I => \N__28307\
        );

    \I__6969\ : ClkMux
    port map (
            O => \N__28531\,
            I => \N__28307\
        );

    \I__6968\ : ClkMux
    port map (
            O => \N__28530\,
            I => \N__28307\
        );

    \I__6967\ : ClkMux
    port map (
            O => \N__28529\,
            I => \N__28307\
        );

    \I__6966\ : ClkMux
    port map (
            O => \N__28528\,
            I => \N__28307\
        );

    \I__6965\ : ClkMux
    port map (
            O => \N__28527\,
            I => \N__28307\
        );

    \I__6964\ : ClkMux
    port map (
            O => \N__28526\,
            I => \N__28307\
        );

    \I__6963\ : ClkMux
    port map (
            O => \N__28525\,
            I => \N__28307\
        );

    \I__6962\ : ClkMux
    port map (
            O => \N__28524\,
            I => \N__28307\
        );

    \I__6961\ : ClkMux
    port map (
            O => \N__28523\,
            I => \N__28307\
        );

    \I__6960\ : ClkMux
    port map (
            O => \N__28522\,
            I => \N__28307\
        );

    \I__6959\ : ClkMux
    port map (
            O => \N__28521\,
            I => \N__28307\
        );

    \I__6958\ : ClkMux
    port map (
            O => \N__28520\,
            I => \N__28307\
        );

    \I__6957\ : ClkMux
    port map (
            O => \N__28519\,
            I => \N__28307\
        );

    \I__6956\ : ClkMux
    port map (
            O => \N__28518\,
            I => \N__28307\
        );

    \I__6955\ : ClkMux
    port map (
            O => \N__28517\,
            I => \N__28307\
        );

    \I__6954\ : ClkMux
    port map (
            O => \N__28516\,
            I => \N__28307\
        );

    \I__6953\ : ClkMux
    port map (
            O => \N__28515\,
            I => \N__28307\
        );

    \I__6952\ : ClkMux
    port map (
            O => \N__28514\,
            I => \N__28307\
        );

    \I__6951\ : ClkMux
    port map (
            O => \N__28513\,
            I => \N__28307\
        );

    \I__6950\ : ClkMux
    port map (
            O => \N__28512\,
            I => \N__28307\
        );

    \I__6949\ : ClkMux
    port map (
            O => \N__28511\,
            I => \N__28307\
        );

    \I__6948\ : ClkMux
    port map (
            O => \N__28510\,
            I => \N__28307\
        );

    \I__6947\ : ClkMux
    port map (
            O => \N__28509\,
            I => \N__28307\
        );

    \I__6946\ : ClkMux
    port map (
            O => \N__28508\,
            I => \N__28307\
        );

    \I__6945\ : ClkMux
    port map (
            O => \N__28507\,
            I => \N__28307\
        );

    \I__6944\ : ClkMux
    port map (
            O => \N__28506\,
            I => \N__28307\
        );

    \I__6943\ : ClkMux
    port map (
            O => \N__28505\,
            I => \N__28307\
        );

    \I__6942\ : ClkMux
    port map (
            O => \N__28504\,
            I => \N__28307\
        );

    \I__6941\ : ClkMux
    port map (
            O => \N__28503\,
            I => \N__28307\
        );

    \I__6940\ : ClkMux
    port map (
            O => \N__28502\,
            I => \N__28307\
        );

    \I__6939\ : ClkMux
    port map (
            O => \N__28501\,
            I => \N__28307\
        );

    \I__6938\ : ClkMux
    port map (
            O => \N__28500\,
            I => \N__28307\
        );

    \I__6937\ : ClkMux
    port map (
            O => \N__28499\,
            I => \N__28307\
        );

    \I__6936\ : ClkMux
    port map (
            O => \N__28498\,
            I => \N__28307\
        );

    \I__6935\ : ClkMux
    port map (
            O => \N__28497\,
            I => \N__28307\
        );

    \I__6934\ : ClkMux
    port map (
            O => \N__28496\,
            I => \N__28307\
        );

    \I__6933\ : ClkMux
    port map (
            O => \N__28495\,
            I => \N__28307\
        );

    \I__6932\ : ClkMux
    port map (
            O => \N__28494\,
            I => \N__28307\
        );

    \I__6931\ : ClkMux
    port map (
            O => \N__28493\,
            I => \N__28307\
        );

    \I__6930\ : ClkMux
    port map (
            O => \N__28492\,
            I => \N__28307\
        );

    \I__6929\ : ClkMux
    port map (
            O => \N__28491\,
            I => \N__28307\
        );

    \I__6928\ : ClkMux
    port map (
            O => \N__28490\,
            I => \N__28307\
        );

    \I__6927\ : ClkMux
    port map (
            O => \N__28489\,
            I => \N__28307\
        );

    \I__6926\ : ClkMux
    port map (
            O => \N__28488\,
            I => \N__28307\
        );

    \I__6925\ : ClkMux
    port map (
            O => \N__28487\,
            I => \N__28307\
        );

    \I__6924\ : ClkMux
    port map (
            O => \N__28486\,
            I => \N__28307\
        );

    \I__6923\ : ClkMux
    port map (
            O => \N__28485\,
            I => \N__28307\
        );

    \I__6922\ : ClkMux
    port map (
            O => \N__28484\,
            I => \N__28307\
        );

    \I__6921\ : ClkMux
    port map (
            O => \N__28483\,
            I => \N__28307\
        );

    \I__6920\ : ClkMux
    port map (
            O => \N__28482\,
            I => \N__28307\
        );

    \I__6919\ : ClkMux
    port map (
            O => \N__28481\,
            I => \N__28307\
        );

    \I__6918\ : ClkMux
    port map (
            O => \N__28480\,
            I => \N__28307\
        );

    \I__6917\ : ClkMux
    port map (
            O => \N__28479\,
            I => \N__28307\
        );

    \I__6916\ : ClkMux
    port map (
            O => \N__28478\,
            I => \N__28307\
        );

    \I__6915\ : ClkMux
    port map (
            O => \N__28477\,
            I => \N__28307\
        );

    \I__6914\ : ClkMux
    port map (
            O => \N__28476\,
            I => \N__28307\
        );

    \I__6913\ : ClkMux
    port map (
            O => \N__28475\,
            I => \N__28307\
        );

    \I__6912\ : ClkMux
    port map (
            O => \N__28474\,
            I => \N__28307\
        );

    \I__6911\ : ClkMux
    port map (
            O => \N__28473\,
            I => \N__28307\
        );

    \I__6910\ : ClkMux
    port map (
            O => \N__28472\,
            I => \N__28307\
        );

    \I__6909\ : ClkMux
    port map (
            O => \N__28471\,
            I => \N__28307\
        );

    \I__6908\ : ClkMux
    port map (
            O => \N__28470\,
            I => \N__28307\
        );

    \I__6907\ : ClkMux
    port map (
            O => \N__28469\,
            I => \N__28307\
        );

    \I__6906\ : ClkMux
    port map (
            O => \N__28468\,
            I => \N__28307\
        );

    \I__6905\ : ClkMux
    port map (
            O => \N__28467\,
            I => \N__28307\
        );

    \I__6904\ : ClkMux
    port map (
            O => \N__28466\,
            I => \N__28307\
        );

    \I__6903\ : GlobalMux
    port map (
            O => \N__28307\,
            I => \N__28304\
        );

    \I__6902\ : DummyBuf
    port map (
            O => \N__28304\,
            I => clk
        );

    \I__6901\ : CEMux
    port map (
            O => \N__28301\,
            I => \N__28297\
        );

    \I__6900\ : CEMux
    port map (
            O => \N__28300\,
            I => \N__28293\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28289\
        );

    \I__6898\ : CEMux
    port map (
            O => \N__28296\,
            I => \N__28286\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__28293\,
            I => \N__28282\
        );

    \I__6896\ : CEMux
    port map (
            O => \N__28292\,
            I => \N__28279\
        );

    \I__6895\ : Span4Mux_s3_h
    port map (
            O => \N__28289\,
            I => \N__28274\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__28286\,
            I => \N__28274\
        );

    \I__6893\ : CEMux
    port map (
            O => \N__28285\,
            I => \N__28271\
        );

    \I__6892\ : Span4Mux_h
    port map (
            O => \N__28282\,
            I => \N__28268\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__28279\,
            I => \N__28265\
        );

    \I__6890\ : Span4Mux_v
    port map (
            O => \N__28274\,
            I => \N__28262\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__28271\,
            I => \N__28259\
        );

    \I__6888\ : Span4Mux_s1_h
    port map (
            O => \N__28268\,
            I => \N__28254\
        );

    \I__6887\ : Span4Mux_v
    port map (
            O => \N__28265\,
            I => \N__28254\
        );

    \I__6886\ : Span4Mux_v
    port map (
            O => \N__28262\,
            I => \N__28251\
        );

    \I__6885\ : Span4Mux_v
    port map (
            O => \N__28259\,
            I => \N__28246\
        );

    \I__6884\ : Span4Mux_h
    port map (
            O => \N__28254\,
            I => \N__28246\
        );

    \I__6883\ : Sp12to4
    port map (
            O => \N__28251\,
            I => \N__28243\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__28246\,
            I => \tok.n995\
        );

    \I__6881\ : Odrv12
    port map (
            O => \N__28243\,
            I => \tok.n995\
        );

    \I__6880\ : SRMux
    port map (
            O => \N__28238\,
            I => \N__28227\
        );

    \I__6879\ : SRMux
    port map (
            O => \N__28237\,
            I => \N__28223\
        );

    \I__6878\ : SRMux
    port map (
            O => \N__28236\,
            I => \N__28220\
        );

    \I__6877\ : SRMux
    port map (
            O => \N__28235\,
            I => \N__28217\
        );

    \I__6876\ : SRMux
    port map (
            O => \N__28234\,
            I => \N__28214\
        );

    \I__6875\ : SRMux
    port map (
            O => \N__28233\,
            I => \N__28209\
        );

    \I__6874\ : SRMux
    port map (
            O => \N__28232\,
            I => \N__28206\
        );

    \I__6873\ : SRMux
    port map (
            O => \N__28231\,
            I => \N__28202\
        );

    \I__6872\ : SRMux
    port map (
            O => \N__28230\,
            I => \N__28199\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__28227\,
            I => \N__28196\
        );

    \I__6870\ : SRMux
    port map (
            O => \N__28226\,
            I => \N__28193\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__28223\,
            I => \N__28189\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__28220\,
            I => \N__28186\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__28217\,
            I => \N__28181\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__28214\,
            I => \N__28181\
        );

    \I__6865\ : SRMux
    port map (
            O => \N__28213\,
            I => \N__28178\
        );

    \I__6864\ : SRMux
    port map (
            O => \N__28212\,
            I => \N__28175\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__28209\,
            I => \N__28171\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__28206\,
            I => \N__28168\
        );

    \I__6861\ : SRMux
    port map (
            O => \N__28205\,
            I => \N__28165\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__28202\,
            I => \N__28162\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__28199\,
            I => \N__28159\
        );

    \I__6858\ : Span4Mux_v
    port map (
            O => \N__28196\,
            I => \N__28154\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__28193\,
            I => \N__28154\
        );

    \I__6856\ : SRMux
    port map (
            O => \N__28192\,
            I => \N__28151\
        );

    \I__6855\ : Span4Mux_h
    port map (
            O => \N__28189\,
            I => \N__28140\
        );

    \I__6854\ : Span4Mux_h
    port map (
            O => \N__28186\,
            I => \N__28140\
        );

    \I__6853\ : Span4Mux_s3_v
    port map (
            O => \N__28181\,
            I => \N__28140\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__28178\,
            I => \N__28140\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__28175\,
            I => \N__28140\
        );

    \I__6850\ : SRMux
    port map (
            O => \N__28174\,
            I => \N__28137\
        );

    \I__6849\ : Span4Mux_v
    port map (
            O => \N__28171\,
            I => \N__28134\
        );

    \I__6848\ : Span4Mux_v
    port map (
            O => \N__28168\,
            I => \N__28129\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__28165\,
            I => \N__28129\
        );

    \I__6846\ : Span4Mux_s3_h
    port map (
            O => \N__28162\,
            I => \N__28125\
        );

    \I__6845\ : Span4Mux_v
    port map (
            O => \N__28159\,
            I => \N__28122\
        );

    \I__6844\ : Span4Mux_h
    port map (
            O => \N__28154\,
            I => \N__28117\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28117\
        );

    \I__6842\ : Span4Mux_v
    port map (
            O => \N__28140\,
            I => \N__28114\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__28137\,
            I => \N__28111\
        );

    \I__6840\ : Span4Mux_v
    port map (
            O => \N__28134\,
            I => \N__28108\
        );

    \I__6839\ : Span4Mux_v
    port map (
            O => \N__28129\,
            I => \N__28105\
        );

    \I__6838\ : SRMux
    port map (
            O => \N__28128\,
            I => \N__28102\
        );

    \I__6837\ : Span4Mux_h
    port map (
            O => \N__28125\,
            I => \N__28099\
        );

    \I__6836\ : Span4Mux_h
    port map (
            O => \N__28122\,
            I => \N__28094\
        );

    \I__6835\ : Span4Mux_h
    port map (
            O => \N__28117\,
            I => \N__28094\
        );

    \I__6834\ : Span4Mux_v
    port map (
            O => \N__28114\,
            I => \N__28089\
        );

    \I__6833\ : Span4Mux_h
    port map (
            O => \N__28111\,
            I => \N__28089\
        );

    \I__6832\ : Span4Mux_h
    port map (
            O => \N__28108\,
            I => \N__28082\
        );

    \I__6831\ : Span4Mux_v
    port map (
            O => \N__28105\,
            I => \N__28082\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__28102\,
            I => \N__28082\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__28099\,
            I => \tok.reset_N_2\
        );

    \I__6828\ : Odrv4
    port map (
            O => \N__28094\,
            I => \tok.reset_N_2\
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__28089\,
            I => \tok.reset_N_2\
        );

    \I__6826\ : Odrv4
    port map (
            O => \N__28082\,
            I => \tok.reset_N_2\
        );

    \I__6825\ : CascadeMux
    port map (
            O => \N__28073\,
            I => \N__28068\
        );

    \I__6824\ : InMux
    port map (
            O => \N__28072\,
            I => \N__28061\
        );

    \I__6823\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28061\
        );

    \I__6822\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28058\
        );

    \I__6821\ : CascadeMux
    port map (
            O => \N__28067\,
            I => \N__28054\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__28066\,
            I => \N__28051\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__28061\,
            I => \N__28048\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__28058\,
            I => \N__28045\
        );

    \I__6817\ : InMux
    port map (
            O => \N__28057\,
            I => \N__28042\
        );

    \I__6816\ : InMux
    port map (
            O => \N__28054\,
            I => \N__28039\
        );

    \I__6815\ : InMux
    port map (
            O => \N__28051\,
            I => \N__28036\
        );

    \I__6814\ : Span4Mux_v
    port map (
            O => \N__28048\,
            I => \N__28032\
        );

    \I__6813\ : Span4Mux_v
    port map (
            O => \N__28045\,
            I => \N__28029\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__28042\,
            I => \N__28025\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__28039\,
            I => \N__28022\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__28036\,
            I => \N__28019\
        );

    \I__6809\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28016\
        );

    \I__6808\ : Span4Mux_s1_h
    port map (
            O => \N__28032\,
            I => \N__28013\
        );

    \I__6807\ : Span4Mux_h
    port map (
            O => \N__28029\,
            I => \N__28010\
        );

    \I__6806\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28007\
        );

    \I__6805\ : Span4Mux_h
    port map (
            O => \N__28025\,
            I => \N__28004\
        );

    \I__6804\ : Span4Mux_v
    port map (
            O => \N__28022\,
            I => \N__27999\
        );

    \I__6803\ : Span4Mux_h
    port map (
            O => \N__28019\,
            I => \N__27999\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__28016\,
            I => \tok.S_8\
        );

    \I__6801\ : Odrv4
    port map (
            O => \N__28013\,
            I => \tok.S_8\
        );

    \I__6800\ : Odrv4
    port map (
            O => \N__28010\,
            I => \tok.S_8\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__28007\,
            I => \tok.S_8\
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__28004\,
            I => \tok.S_8\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__27999\,
            I => \tok.S_8\
        );

    \I__6796\ : CascadeMux
    port map (
            O => \N__27986\,
            I => \N__27983\
        );

    \I__6795\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27980\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__27980\,
            I => \tok.n5544\
        );

    \I__6793\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27974\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__27974\,
            I => \tok.n5542\
        );

    \I__6791\ : InMux
    port map (
            O => \N__27971\,
            I => \N__27968\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__6789\ : Span4Mux_v
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__6788\ : Odrv4
    port map (
            O => \N__27962\,
            I => \tok.n10_adj_666\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__27959\,
            I => \N__27954\
        );

    \I__6786\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27950\
        );

    \I__6785\ : InMux
    port map (
            O => \N__27957\,
            I => \N__27947\
        );

    \I__6784\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27944\
        );

    \I__6783\ : CascadeMux
    port map (
            O => \N__27953\,
            I => \N__27941\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__27950\,
            I => \N__27935\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__27947\,
            I => \N__27935\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__27944\,
            I => \N__27932\
        );

    \I__6779\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27929\
        );

    \I__6778\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27926\
        );

    \I__6777\ : Span4Mux_v
    port map (
            O => \N__27935\,
            I => \N__27923\
        );

    \I__6776\ : Span4Mux_s3_v
    port map (
            O => \N__27932\,
            I => \N__27918\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27918\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27915\
        );

    \I__6773\ : Span4Mux_h
    port map (
            O => \N__27923\,
            I => \N__27908\
        );

    \I__6772\ : Span4Mux_v
    port map (
            O => \N__27918\,
            I => \N__27908\
        );

    \I__6771\ : Span4Mux_v
    port map (
            O => \N__27915\,
            I => \N__27905\
        );

    \I__6770\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27900\
        );

    \I__6769\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27900\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__27908\,
            I => \tok.n15_adj_667\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__27905\,
            I => \tok.n15_adj_667\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__27900\,
            I => \tok.n15_adj_667\
        );

    \I__6765\ : InMux
    port map (
            O => \N__27893\,
            I => \N__27890\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__27890\,
            I => \tok.n14_adj_668\
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__27887\,
            I => \N__27879\
        );

    \I__6762\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27869\
        );

    \I__6761\ : InMux
    port map (
            O => \N__27885\,
            I => \N__27869\
        );

    \I__6760\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27864\
        );

    \I__6759\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27864\
        );

    \I__6758\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27859\
        );

    \I__6757\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27859\
        );

    \I__6756\ : CascadeMux
    port map (
            O => \N__27878\,
            I => \N__27851\
        );

    \I__6755\ : InMux
    port map (
            O => \N__27877\,
            I => \N__27847\
        );

    \I__6754\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27840\
        );

    \I__6753\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27840\
        );

    \I__6752\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27840\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__27869\,
            I => \N__27835\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__27864\,
            I => \N__27835\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__27859\,
            I => \N__27832\
        );

    \I__6748\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27825\
        );

    \I__6747\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27825\
        );

    \I__6746\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27825\
        );

    \I__6745\ : InMux
    port map (
            O => \N__27855\,
            I => \N__27818\
        );

    \I__6744\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27818\
        );

    \I__6743\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27818\
        );

    \I__6742\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27815\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__27847\,
            I => \N__27810\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__27840\,
            I => \N__27810\
        );

    \I__6739\ : Span4Mux_v
    port map (
            O => \N__27835\,
            I => \N__27807\
        );

    \I__6738\ : Span4Mux_h
    port map (
            O => \N__27832\,
            I => \N__27800\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__27825\,
            I => \N__27800\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__27818\,
            I => \N__27800\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__27815\,
            I => \N__27797\
        );

    \I__6734\ : Span4Mux_v
    port map (
            O => \N__27810\,
            I => \N__27790\
        );

    \I__6733\ : Span4Mux_h
    port map (
            O => \N__27807\,
            I => \N__27790\
        );

    \I__6732\ : Span4Mux_v
    port map (
            O => \N__27800\,
            I => \N__27790\
        );

    \I__6731\ : Odrv4
    port map (
            O => \N__27797\,
            I => \tok.n880\
        );

    \I__6730\ : Odrv4
    port map (
            O => \N__27790\,
            I => \tok.n880\
        );

    \I__6729\ : InMux
    port map (
            O => \N__27785\,
            I => \N__27775\
        );

    \I__6728\ : InMux
    port map (
            O => \N__27784\,
            I => \N__27775\
        );

    \I__6727\ : InMux
    port map (
            O => \N__27783\,
            I => \N__27771\
        );

    \I__6726\ : CascadeMux
    port map (
            O => \N__27782\,
            I => \N__27767\
        );

    \I__6725\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27763\
        );

    \I__6724\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27760\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__27775\,
            I => \N__27757\
        );

    \I__6722\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27751\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__27771\,
            I => \N__27748\
        );

    \I__6720\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27745\
        );

    \I__6719\ : InMux
    port map (
            O => \N__27767\,
            I => \N__27742\
        );

    \I__6718\ : InMux
    port map (
            O => \N__27766\,
            I => \N__27739\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__27763\,
            I => \N__27735\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__27760\,
            I => \N__27732\
        );

    \I__6715\ : Span4Mux_s2_h
    port map (
            O => \N__27757\,
            I => \N__27729\
        );

    \I__6714\ : InMux
    port map (
            O => \N__27756\,
            I => \N__27726\
        );

    \I__6713\ : InMux
    port map (
            O => \N__27755\,
            I => \N__27722\
        );

    \I__6712\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27719\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__27751\,
            I => \N__27716\
        );

    \I__6710\ : Span4Mux_s2_v
    port map (
            O => \N__27748\,
            I => \N__27709\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__27745\,
            I => \N__27709\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__27742\,
            I => \N__27709\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__27739\,
            I => \N__27706\
        );

    \I__6706\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27703\
        );

    \I__6705\ : Span4Mux_v
    port map (
            O => \N__27735\,
            I => \N__27694\
        );

    \I__6704\ : Span4Mux_v
    port map (
            O => \N__27732\,
            I => \N__27694\
        );

    \I__6703\ : Span4Mux_h
    port map (
            O => \N__27729\,
            I => \N__27694\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__27726\,
            I => \N__27694\
        );

    \I__6701\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27691\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__27722\,
            I => \N__27687\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__27719\,
            I => \N__27676\
        );

    \I__6698\ : Span4Mux_v
    port map (
            O => \N__27716\,
            I => \N__27676\
        );

    \I__6697\ : Span4Mux_v
    port map (
            O => \N__27709\,
            I => \N__27676\
        );

    \I__6696\ : Span4Mux_v
    port map (
            O => \N__27706\,
            I => \N__27676\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__27703\,
            I => \N__27676\
        );

    \I__6694\ : Span4Mux_h
    port map (
            O => \N__27694\,
            I => \N__27671\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__27691\,
            I => \N__27671\
        );

    \I__6692\ : InMux
    port map (
            O => \N__27690\,
            I => \N__27668\
        );

    \I__6691\ : Span4Mux_h
    port map (
            O => \N__27687\,
            I => \N__27663\
        );

    \I__6690\ : Span4Mux_h
    port map (
            O => \N__27676\,
            I => \N__27663\
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__27671\,
            I => \tok.A_low_0\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__27668\,
            I => \tok.A_low_0\
        );

    \I__6687\ : Odrv4
    port map (
            O => \N__27663\,
            I => \tok.A_low_0\
        );

    \I__6686\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27644\
        );

    \I__6685\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27644\
        );

    \I__6684\ : InMux
    port map (
            O => \N__27654\,
            I => \N__27639\
        );

    \I__6683\ : InMux
    port map (
            O => \N__27653\,
            I => \N__27639\
        );

    \I__6682\ : InMux
    port map (
            O => \N__27652\,
            I => \N__27634\
        );

    \I__6681\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27634\
        );

    \I__6680\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27626\
        );

    \I__6679\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27621\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__27644\,
            I => \N__27618\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__27639\,
            I => \N__27615\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__27634\,
            I => \N__27612\
        );

    \I__6675\ : InMux
    port map (
            O => \N__27633\,
            I => \N__27609\
        );

    \I__6674\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27602\
        );

    \I__6673\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27602\
        );

    \I__6672\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27602\
        );

    \I__6671\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27599\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__27626\,
            I => \N__27596\
        );

    \I__6669\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27593\
        );

    \I__6668\ : InMux
    port map (
            O => \N__27624\,
            I => \N__27590\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__27621\,
            I => \N__27587\
        );

    \I__6666\ : Span4Mux_s1_h
    port map (
            O => \N__27618\,
            I => \N__27582\
        );

    \I__6665\ : Span4Mux_v
    port map (
            O => \N__27615\,
            I => \N__27582\
        );

    \I__6664\ : Odrv4
    port map (
            O => \N__27612\,
            I => \tok.n904\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__27609\,
            I => \tok.n904\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__27602\,
            I => \tok.n904\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__27599\,
            I => \tok.n904\
        );

    \I__6660\ : Odrv4
    port map (
            O => \N__27596\,
            I => \tok.n904\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__27593\,
            I => \tok.n904\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__27590\,
            I => \tok.n904\
        );

    \I__6657\ : Odrv4
    port map (
            O => \N__27587\,
            I => \tok.n904\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__27582\,
            I => \tok.n904\
        );

    \I__6655\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27560\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__27560\,
            I => \N__27557\
        );

    \I__6653\ : Odrv12
    port map (
            O => \N__27557\,
            I => \tok.n5372\
        );

    \I__6652\ : CascadeMux
    port map (
            O => \N__27554\,
            I => \N__27551\
        );

    \I__6651\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27546\
        );

    \I__6650\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27540\
        );

    \I__6649\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27540\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__27546\,
            I => \N__27535\
        );

    \I__6647\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27532\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__27540\,
            I => \N__27528\
        );

    \I__6645\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27525\
        );

    \I__6644\ : InMux
    port map (
            O => \N__27538\,
            I => \N__27522\
        );

    \I__6643\ : Span4Mux_s1_h
    port map (
            O => \N__27535\,
            I => \N__27517\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__27532\,
            I => \N__27517\
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__27531\,
            I => \N__27514\
        );

    \I__6640\ : Span4Mux_v
    port map (
            O => \N__27528\,
            I => \N__27510\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__27525\,
            I => \N__27507\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__27522\,
            I => \N__27504\
        );

    \I__6637\ : Span4Mux_h
    port map (
            O => \N__27517\,
            I => \N__27501\
        );

    \I__6636\ : InMux
    port map (
            O => \N__27514\,
            I => \N__27498\
        );

    \I__6635\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27495\
        );

    \I__6634\ : Span4Mux_v
    port map (
            O => \N__27510\,
            I => \N__27490\
        );

    \I__6633\ : Span4Mux_v
    port map (
            O => \N__27507\,
            I => \N__27490\
        );

    \I__6632\ : Span12Mux_s8_h
    port map (
            O => \N__27504\,
            I => \N__27483\
        );

    \I__6631\ : Sp12to4
    port map (
            O => \N__27501\,
            I => \N__27483\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__27498\,
            I => \N__27483\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__27495\,
            I => \tok.S_9\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__27490\,
            I => \tok.S_9\
        );

    \I__6627\ : Odrv12
    port map (
            O => \N__27483\,
            I => \tok.S_9\
        );

    \I__6626\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27473\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__27473\,
            I => \N__27470\
        );

    \I__6624\ : Span4Mux_v
    port map (
            O => \N__27470\,
            I => \N__27467\
        );

    \I__6623\ : Odrv4
    port map (
            O => \N__27467\,
            I => \tok.n8_adj_689\
        );

    \I__6622\ : CascadeMux
    port map (
            O => \N__27464\,
            I => \N__27461\
        );

    \I__6621\ : InMux
    port map (
            O => \N__27461\,
            I => \N__27456\
        );

    \I__6620\ : CascadeMux
    port map (
            O => \N__27460\,
            I => \N__27453\
        );

    \I__6619\ : CascadeMux
    port map (
            O => \N__27459\,
            I => \N__27449\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__27456\,
            I => \N__27445\
        );

    \I__6617\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27442\
        );

    \I__6616\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27437\
        );

    \I__6615\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27434\
        );

    \I__6614\ : CascadeMux
    port map (
            O => \N__27448\,
            I => \N__27431\
        );

    \I__6613\ : Span4Mux_v
    port map (
            O => \N__27445\,
            I => \N__27426\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27426\
        );

    \I__6611\ : InMux
    port map (
            O => \N__27441\,
            I => \N__27423\
        );

    \I__6610\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27420\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__27437\,
            I => \N__27415\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__27434\,
            I => \N__27415\
        );

    \I__6607\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27411\
        );

    \I__6606\ : Span4Mux_v
    port map (
            O => \N__27426\,
            I => \N__27408\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__27423\,
            I => \N__27405\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__27420\,
            I => \N__27402\
        );

    \I__6603\ : Span4Mux_v
    port map (
            O => \N__27415\,
            I => \N__27399\
        );

    \I__6602\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27396\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__27411\,
            I => \N__27393\
        );

    \I__6600\ : Span4Mux_h
    port map (
            O => \N__27408\,
            I => \N__27390\
        );

    \I__6599\ : Span4Mux_v
    port map (
            O => \N__27405\,
            I => \N__27387\
        );

    \I__6598\ : Span4Mux_v
    port map (
            O => \N__27402\,
            I => \N__27382\
        );

    \I__6597\ : Span4Mux_h
    port map (
            O => \N__27399\,
            I => \N__27382\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__27396\,
            I => \tok.S_10\
        );

    \I__6595\ : Odrv12
    port map (
            O => \N__27393\,
            I => \tok.S_10\
        );

    \I__6594\ : Odrv4
    port map (
            O => \N__27390\,
            I => \tok.S_10\
        );

    \I__6593\ : Odrv4
    port map (
            O => \N__27387\,
            I => \tok.S_10\
        );

    \I__6592\ : Odrv4
    port map (
            O => \N__27382\,
            I => \tok.S_10\
        );

    \I__6591\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27368\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__27368\,
            I => \N__27365\
        );

    \I__6589\ : Odrv12
    port map (
            O => \N__27365\,
            I => \tok.n8_adj_702\
        );

    \I__6588\ : CascadeMux
    port map (
            O => \N__27362\,
            I => \N__27359\
        );

    \I__6587\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27356\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__27356\,
            I => \tok.n298\
        );

    \I__6585\ : CascadeMux
    port map (
            O => \N__27353\,
            I => \N__27348\
        );

    \I__6584\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27344\
        );

    \I__6583\ : CascadeMux
    port map (
            O => \N__27351\,
            I => \N__27340\
        );

    \I__6582\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27337\
        );

    \I__6581\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27334\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__27344\,
            I => \N__27331\
        );

    \I__6579\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27328\
        );

    \I__6578\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27321\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__27337\,
            I => \N__27318\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__27334\,
            I => \N__27313\
        );

    \I__6575\ : Span4Mux_h
    port map (
            O => \N__27331\,
            I => \N__27313\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__27328\,
            I => \N__27310\
        );

    \I__6573\ : InMux
    port map (
            O => \N__27327\,
            I => \N__27307\
        );

    \I__6572\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27304\
        );

    \I__6571\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27298\
        );

    \I__6570\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27298\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__27321\,
            I => \N__27293\
        );

    \I__6568\ : Span4Mux_h
    port map (
            O => \N__27318\,
            I => \N__27287\
        );

    \I__6567\ : Span4Mux_h
    port map (
            O => \N__27313\,
            I => \N__27280\
        );

    \I__6566\ : Span4Mux_s3_v
    port map (
            O => \N__27310\,
            I => \N__27280\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__27307\,
            I => \N__27280\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__27304\,
            I => \N__27277\
        );

    \I__6563\ : InMux
    port map (
            O => \N__27303\,
            I => \N__27274\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__27298\,
            I => \N__27271\
        );

    \I__6561\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27266\
        );

    \I__6560\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27266\
        );

    \I__6559\ : Span4Mux_h
    port map (
            O => \N__27293\,
            I => \N__27263\
        );

    \I__6558\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27260\
        );

    \I__6557\ : InMux
    port map (
            O => \N__27291\,
            I => \N__27255\
        );

    \I__6556\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27255\
        );

    \I__6555\ : Span4Mux_v
    port map (
            O => \N__27287\,
            I => \N__27250\
        );

    \I__6554\ : Span4Mux_v
    port map (
            O => \N__27280\,
            I => \N__27250\
        );

    \I__6553\ : Span12Mux_s7_v
    port map (
            O => \N__27277\,
            I => \N__27245\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__27274\,
            I => \N__27245\
        );

    \I__6551\ : Span4Mux_h
    port map (
            O => \N__27271\,
            I => \N__27238\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27238\
        );

    \I__6549\ : Span4Mux_h
    port map (
            O => \N__27263\,
            I => \N__27238\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__27260\,
            I => \tok.A_low_5\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__27255\,
            I => \tok.A_low_5\
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__27250\,
            I => \tok.A_low_5\
        );

    \I__6545\ : Odrv12
    port map (
            O => \N__27245\,
            I => \tok.A_low_5\
        );

    \I__6544\ : Odrv4
    port map (
            O => \N__27238\,
            I => \tok.A_low_5\
        );

    \I__6543\ : InMux
    port map (
            O => \N__27227\,
            I => \N__27224\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__27224\,
            I => \tok.n297\
        );

    \I__6541\ : CascadeMux
    port map (
            O => \N__27221\,
            I => \N__27218\
        );

    \I__6540\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27215\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__27215\,
            I => \N__27210\
        );

    \I__6538\ : CascadeMux
    port map (
            O => \N__27214\,
            I => \N__27206\
        );

    \I__6537\ : InMux
    port map (
            O => \N__27213\,
            I => \N__27203\
        );

    \I__6536\ : Span4Mux_s3_v
    port map (
            O => \N__27210\,
            I => \N__27200\
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__27209\,
            I => \N__27197\
        );

    \I__6534\ : InMux
    port map (
            O => \N__27206\,
            I => \N__27192\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__27203\,
            I => \N__27189\
        );

    \I__6532\ : Span4Mux_v
    port map (
            O => \N__27200\,
            I => \N__27184\
        );

    \I__6531\ : InMux
    port map (
            O => \N__27197\,
            I => \N__27181\
        );

    \I__6530\ : CascadeMux
    port map (
            O => \N__27196\,
            I => \N__27177\
        );

    \I__6529\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27174\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__27192\,
            I => \N__27171\
        );

    \I__6527\ : Span4Mux_v
    port map (
            O => \N__27189\,
            I => \N__27168\
        );

    \I__6526\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27165\
        );

    \I__6525\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27162\
        );

    \I__6524\ : Span4Mux_h
    port map (
            O => \N__27184\,
            I => \N__27157\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__27181\,
            I => \N__27157\
        );

    \I__6522\ : InMux
    port map (
            O => \N__27180\,
            I => \N__27154\
        );

    \I__6521\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27151\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__27174\,
            I => \N__27146\
        );

    \I__6519\ : Span4Mux_h
    port map (
            O => \N__27171\,
            I => \N__27146\
        );

    \I__6518\ : Span4Mux_h
    port map (
            O => \N__27168\,
            I => \N__27141\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__27165\,
            I => \N__27141\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__27162\,
            I => \N__27136\
        );

    \I__6515\ : Span4Mux_h
    port map (
            O => \N__27157\,
            I => \N__27136\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__27154\,
            I => \tok.S_5\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__27151\,
            I => \tok.S_5\
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__27146\,
            I => \tok.S_5\
        );

    \I__6511\ : Odrv4
    port map (
            O => \N__27141\,
            I => \tok.S_5\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__27136\,
            I => \tok.S_5\
        );

    \I__6509\ : CascadeMux
    port map (
            O => \N__27125\,
            I => \N__27121\
        );

    \I__6508\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27116\
        );

    \I__6507\ : InMux
    port map (
            O => \N__27121\,
            I => \N__27116\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__27116\,
            I => uart_rx_data_5
        );

    \I__6505\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27110\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__27110\,
            I => \tok.n6_adj_717\
        );

    \I__6503\ : CascadeMux
    port map (
            O => \N__27107\,
            I => \N__27103\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__27106\,
            I => \N__27100\
        );

    \I__6501\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27097\
        );

    \I__6500\ : InMux
    port map (
            O => \N__27100\,
            I => \N__27094\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__27097\,
            I => \N__27091\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__27094\,
            I => \N__27088\
        );

    \I__6497\ : Span12Mux_s10_h
    port map (
            O => \N__27091\,
            I => \N__27085\
        );

    \I__6496\ : Span4Mux_v
    port map (
            O => \N__27088\,
            I => \N__27082\
        );

    \I__6495\ : Odrv12
    port map (
            O => \N__27085\,
            I => \tok.table_rd_5\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__27082\,
            I => \tok.table_rd_5\
        );

    \I__6493\ : InMux
    port map (
            O => \N__27077\,
            I => \N__27074\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__27074\,
            I => \tok.n16_adj_855\
        );

    \I__6491\ : InMux
    port map (
            O => \N__27071\,
            I => \N__27068\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__27068\,
            I => \N__27065\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__27065\,
            I => \N__27062\
        );

    \I__6488\ : Span4Mux_h
    port map (
            O => \N__27062\,
            I => \N__27059\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__27059\,
            I => \tok.n5_adj_800\
        );

    \I__6486\ : InMux
    port map (
            O => \N__27056\,
            I => \N__27053\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__27053\,
            I => \N__27050\
        );

    \I__6484\ : Span4Mux_h
    port map (
            O => \N__27050\,
            I => \N__27047\
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__27047\,
            I => \tok.n10_adj_823\
        );

    \I__6482\ : CascadeMux
    port map (
            O => \N__27044\,
            I => \tok.n20_adj_857_cascade_\
        );

    \I__6481\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27038\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__27038\,
            I => \tok.n14_adj_856\
        );

    \I__6479\ : InMux
    port map (
            O => \N__27035\,
            I => \N__27032\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__6477\ : Odrv4
    port map (
            O => \N__27029\,
            I => \tok.n5559\
        );

    \I__6476\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27023\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__27023\,
            I => \N__27020\
        );

    \I__6474\ : Span4Mux_s1_h
    port map (
            O => \N__27020\,
            I => \N__27017\
        );

    \I__6473\ : Span4Mux_h
    port map (
            O => \N__27017\,
            I => \N__27014\
        );

    \I__6472\ : Odrv4
    port map (
            O => \N__27014\,
            I => \tok.n3_adj_859\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__27011\,
            I => \tok.n22_adj_861_cascade_\
        );

    \I__6470\ : InMux
    port map (
            O => \N__27008\,
            I => \N__27005\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__27005\,
            I => \tok.n18_adj_860\
        );

    \I__6468\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26999\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__26999\,
            I => \tok.n5556\
        );

    \I__6466\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26988\
        );

    \I__6465\ : InMux
    port map (
            O => \N__26995\,
            I => \N__26988\
        );

    \I__6464\ : InMux
    port map (
            O => \N__26994\,
            I => \N__26985\
        );

    \I__6463\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26980\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__26988\,
            I => \N__26976\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__26985\,
            I => \N__26969\
        );

    \I__6460\ : InMux
    port map (
            O => \N__26984\,
            I => \N__26964\
        );

    \I__6459\ : InMux
    port map (
            O => \N__26983\,
            I => \N__26964\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__26980\,
            I => \N__26961\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__26979\,
            I => \N__26955\
        );

    \I__6456\ : Span4Mux_s2_h
    port map (
            O => \N__26976\,
            I => \N__26951\
        );

    \I__6455\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26948\
        );

    \I__6454\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26941\
        );

    \I__6453\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26941\
        );

    \I__6452\ : InMux
    port map (
            O => \N__26972\,
            I => \N__26941\
        );

    \I__6451\ : Span4Mux_v
    port map (
            O => \N__26969\,
            I => \N__26935\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__26964\,
            I => \N__26935\
        );

    \I__6449\ : Span4Mux_h
    port map (
            O => \N__26961\,
            I => \N__26932\
        );

    \I__6448\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26927\
        );

    \I__6447\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26927\
        );

    \I__6446\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26922\
        );

    \I__6445\ : InMux
    port map (
            O => \N__26955\,
            I => \N__26922\
        );

    \I__6444\ : InMux
    port map (
            O => \N__26954\,
            I => \N__26919\
        );

    \I__6443\ : Span4Mux_h
    port map (
            O => \N__26951\,
            I => \N__26914\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__26948\,
            I => \N__26914\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__26941\,
            I => \N__26911\
        );

    \I__6440\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26908\
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__26935\,
            I => \tok.n15\
        );

    \I__6438\ : Odrv4
    port map (
            O => \N__26932\,
            I => \tok.n15\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__26927\,
            I => \tok.n15\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__26922\,
            I => \tok.n15\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__26919\,
            I => \tok.n15\
        );

    \I__6434\ : Odrv4
    port map (
            O => \N__26914\,
            I => \tok.n15\
        );

    \I__6433\ : Odrv4
    port map (
            O => \N__26911\,
            I => \tok.n15\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__26908\,
            I => \tok.n15\
        );

    \I__6431\ : InMux
    port map (
            O => \N__26891\,
            I => \N__26888\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__26888\,
            I => \N__26885\
        );

    \I__6429\ : Odrv12
    port map (
            O => \N__26885\,
            I => \tok.n5_adj_669\
        );

    \I__6428\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26879\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__26879\,
            I => \N__26876\
        );

    \I__6426\ : Span12Mux_s8_v
    port map (
            O => \N__26876\,
            I => \N__26873\
        );

    \I__6425\ : Odrv12
    port map (
            O => \N__26873\,
            I => \tok.table_rd_8\
        );

    \I__6424\ : CascadeMux
    port map (
            O => \N__26870\,
            I => \N__26865\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__26869\,
            I => \N__26861\
        );

    \I__6422\ : InMux
    port map (
            O => \N__26868\,
            I => \N__26839\
        );

    \I__6421\ : InMux
    port map (
            O => \N__26865\,
            I => \N__26839\
        );

    \I__6420\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26839\
        );

    \I__6419\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26839\
        );

    \I__6418\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26839\
        );

    \I__6417\ : InMux
    port map (
            O => \N__26859\,
            I => \N__26839\
        );

    \I__6416\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26839\
        );

    \I__6415\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26830\
        );

    \I__6414\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26830\
        );

    \I__6413\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26830\
        );

    \I__6412\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26830\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__26839\,
            I => \N__26824\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__26830\,
            I => \N__26821\
        );

    \I__6409\ : CascadeMux
    port map (
            O => \N__26829\,
            I => \N__26818\
        );

    \I__6408\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26813\
        );

    \I__6407\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26813\
        );

    \I__6406\ : Span4Mux_h
    port map (
            O => \N__26824\,
            I => \N__26808\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__26821\,
            I => \N__26808\
        );

    \I__6404\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26805\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__26813\,
            I => \N__26802\
        );

    \I__6402\ : Span4Mux_h
    port map (
            O => \N__26808\,
            I => \N__26797\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__26805\,
            I => \N__26797\
        );

    \I__6400\ : Span4Mux_h
    port map (
            O => \N__26802\,
            I => \N__26790\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__26797\,
            I => \N__26790\
        );

    \I__6398\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26785\
        );

    \I__6397\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26785\
        );

    \I__6396\ : Odrv4
    port map (
            O => \N__26790\,
            I => \tok.n4908\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__26785\,
            I => \tok.n4908\
        );

    \I__6394\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26777\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__6392\ : Span4Mux_s2_h
    port map (
            O => \N__26774\,
            I => \N__26771\
        );

    \I__6391\ : Span4Mux_v
    port map (
            O => \N__26771\,
            I => \N__26768\
        );

    \I__6390\ : Odrv4
    port map (
            O => \N__26768\,
            I => \tok.n181\
        );

    \I__6389\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26757\
        );

    \I__6388\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26754\
        );

    \I__6387\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26744\
        );

    \I__6386\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26741\
        );

    \I__6385\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26736\
        );

    \I__6384\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26736\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__26757\,
            I => \N__26733\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26730\
        );

    \I__6381\ : InMux
    port map (
            O => \N__26753\,
            I => \N__26727\
        );

    \I__6380\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26722\
        );

    \I__6379\ : InMux
    port map (
            O => \N__26751\,
            I => \N__26722\
        );

    \I__6378\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26719\
        );

    \I__6377\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26716\
        );

    \I__6376\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26711\
        );

    \I__6375\ : InMux
    port map (
            O => \N__26747\,
            I => \N__26711\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__26744\,
            I => \N__26707\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__26741\,
            I => \N__26704\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__26736\,
            I => \N__26699\
        );

    \I__6371\ : Span4Mux_s3_h
    port map (
            O => \N__26733\,
            I => \N__26699\
        );

    \I__6370\ : Span4Mux_v
    port map (
            O => \N__26730\,
            I => \N__26694\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__26727\,
            I => \N__26694\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__26722\,
            I => \N__26685\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26685\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__26716\,
            I => \N__26685\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__26711\,
            I => \N__26685\
        );

    \I__6364\ : InMux
    port map (
            O => \N__26710\,
            I => \N__26682\
        );

    \I__6363\ : Span4Mux_h
    port map (
            O => \N__26707\,
            I => \N__26679\
        );

    \I__6362\ : Span4Mux_h
    port map (
            O => \N__26704\,
            I => \N__26674\
        );

    \I__6361\ : Span4Mux_h
    port map (
            O => \N__26699\,
            I => \N__26674\
        );

    \I__6360\ : Span4Mux_h
    port map (
            O => \N__26694\,
            I => \N__26667\
        );

    \I__6359\ : Span4Mux_v
    port map (
            O => \N__26685\,
            I => \N__26667\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__26682\,
            I => \N__26667\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__26679\,
            I => \tok.n2735\
        );

    \I__6356\ : Odrv4
    port map (
            O => \N__26674\,
            I => \tok.n2735\
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__26667\,
            I => \tok.n2735\
        );

    \I__6354\ : InMux
    port map (
            O => \N__26660\,
            I => \N__26657\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__26657\,
            I => \tok.n15_adj_670\
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__26654\,
            I => \tok.n13_adj_674_cascade_\
        );

    \I__6351\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26648\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__26648\,
            I => \tok.n5416\
        );

    \I__6349\ : InMux
    port map (
            O => \N__26645\,
            I => \N__26639\
        );

    \I__6348\ : InMux
    port map (
            O => \N__26644\,
            I => \N__26639\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__26639\,
            I => \tok.A_stk.tail_19\
        );

    \I__6346\ : InMux
    port map (
            O => \N__26636\,
            I => \N__26630\
        );

    \I__6345\ : InMux
    port map (
            O => \N__26635\,
            I => \N__26630\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__26630\,
            I => \tok.A_stk.tail_35\
        );

    \I__6343\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26624\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__26624\,
            I => \N__26620\
        );

    \I__6341\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26617\
        );

    \I__6340\ : Span4Mux_s3_h
    port map (
            O => \N__26620\,
            I => \N__26614\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__26617\,
            I => \N__26611\
        );

    \I__6338\ : Odrv4
    port map (
            O => \N__26614\,
            I => \tok.A_stk.tail_67\
        );

    \I__6337\ : Odrv4
    port map (
            O => \N__26611\,
            I => \tok.A_stk.tail_67\
        );

    \I__6336\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26591\
        );

    \I__6335\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26591\
        );

    \I__6334\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26591\
        );

    \I__6333\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26591\
        );

    \I__6332\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26591\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26550\
        );

    \I__6330\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26541\
        );

    \I__6329\ : InMux
    port map (
            O => \N__26589\,
            I => \N__26541\
        );

    \I__6328\ : InMux
    port map (
            O => \N__26588\,
            I => \N__26541\
        );

    \I__6327\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26541\
        );

    \I__6326\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26532\
        );

    \I__6325\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26532\
        );

    \I__6324\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26532\
        );

    \I__6323\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26532\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__26582\,
            I => \N__26513\
        );

    \I__6321\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26503\
        );

    \I__6320\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26486\
        );

    \I__6319\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26486\
        );

    \I__6318\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26486\
        );

    \I__6317\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26486\
        );

    \I__6316\ : InMux
    port map (
            O => \N__26576\,
            I => \N__26486\
        );

    \I__6315\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26486\
        );

    \I__6314\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26486\
        );

    \I__6313\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26473\
        );

    \I__6312\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26473\
        );

    \I__6311\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26473\
        );

    \I__6310\ : InMux
    port map (
            O => \N__26570\,
            I => \N__26473\
        );

    \I__6309\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26473\
        );

    \I__6308\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26473\
        );

    \I__6307\ : InMux
    port map (
            O => \N__26567\,
            I => \N__26456\
        );

    \I__6306\ : InMux
    port map (
            O => \N__26566\,
            I => \N__26456\
        );

    \I__6305\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26456\
        );

    \I__6304\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26456\
        );

    \I__6303\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26456\
        );

    \I__6302\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26456\
        );

    \I__6301\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26456\
        );

    \I__6300\ : InMux
    port map (
            O => \N__26560\,
            I => \N__26456\
        );

    \I__6299\ : InMux
    port map (
            O => \N__26559\,
            I => \N__26434\
        );

    \I__6298\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26434\
        );

    \I__6297\ : InMux
    port map (
            O => \N__26557\,
            I => \N__26434\
        );

    \I__6296\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26434\
        );

    \I__6295\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26434\
        );

    \I__6294\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26434\
        );

    \I__6293\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26434\
        );

    \I__6292\ : Span4Mux_v
    port map (
            O => \N__26550\,
            I => \N__26429\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__26541\,
            I => \N__26429\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__26532\,
            I => \N__26426\
        );

    \I__6289\ : InMux
    port map (
            O => \N__26531\,
            I => \N__26415\
        );

    \I__6288\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26415\
        );

    \I__6287\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26415\
        );

    \I__6286\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26415\
        );

    \I__6285\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26415\
        );

    \I__6284\ : InMux
    port map (
            O => \N__26526\,
            I => \N__26390\
        );

    \I__6283\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26373\
        );

    \I__6282\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26373\
        );

    \I__6281\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26373\
        );

    \I__6280\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26373\
        );

    \I__6279\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26373\
        );

    \I__6278\ : InMux
    port map (
            O => \N__26520\,
            I => \N__26373\
        );

    \I__6277\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26373\
        );

    \I__6276\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26373\
        );

    \I__6275\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26364\
        );

    \I__6274\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26364\
        );

    \I__6273\ : InMux
    port map (
            O => \N__26513\,
            I => \N__26364\
        );

    \I__6272\ : InMux
    port map (
            O => \N__26512\,
            I => \N__26364\
        );

    \I__6271\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26351\
        );

    \I__6270\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26351\
        );

    \I__6269\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26351\
        );

    \I__6268\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26351\
        );

    \I__6267\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26351\
        );

    \I__6266\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26351\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26340\
        );

    \I__6264\ : InMux
    port map (
            O => \N__26502\,
            I => \N__26335\
        );

    \I__6263\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26335\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26332\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__26473\,
            I => \N__26327\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__26456\,
            I => \N__26327\
        );

    \I__6259\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26312\
        );

    \I__6258\ : InMux
    port map (
            O => \N__26454\,
            I => \N__26312\
        );

    \I__6257\ : InMux
    port map (
            O => \N__26453\,
            I => \N__26312\
        );

    \I__6256\ : InMux
    port map (
            O => \N__26452\,
            I => \N__26312\
        );

    \I__6255\ : InMux
    port map (
            O => \N__26451\,
            I => \N__26312\
        );

    \I__6254\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26312\
        );

    \I__6253\ : InMux
    port map (
            O => \N__26449\,
            I => \N__26312\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__26434\,
            I => \N__26309\
        );

    \I__6251\ : Span4Mux_v
    port map (
            O => \N__26429\,
            I => \N__26302\
        );

    \I__6250\ : Span4Mux_s1_h
    port map (
            O => \N__26426\,
            I => \N__26302\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__26415\,
            I => \N__26302\
        );

    \I__6248\ : InMux
    port map (
            O => \N__26414\,
            I => \N__26287\
        );

    \I__6247\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26287\
        );

    \I__6246\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26287\
        );

    \I__6245\ : InMux
    port map (
            O => \N__26411\,
            I => \N__26287\
        );

    \I__6244\ : InMux
    port map (
            O => \N__26410\,
            I => \N__26287\
        );

    \I__6243\ : InMux
    port map (
            O => \N__26409\,
            I => \N__26287\
        );

    \I__6242\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26287\
        );

    \I__6241\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26264\
        );

    \I__6240\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26264\
        );

    \I__6239\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26264\
        );

    \I__6238\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26264\
        );

    \I__6237\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26264\
        );

    \I__6236\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26264\
        );

    \I__6235\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26264\
        );

    \I__6234\ : InMux
    port map (
            O => \N__26400\,
            I => \N__26247\
        );

    \I__6233\ : InMux
    port map (
            O => \N__26399\,
            I => \N__26247\
        );

    \I__6232\ : InMux
    port map (
            O => \N__26398\,
            I => \N__26247\
        );

    \I__6231\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26247\
        );

    \I__6230\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26247\
        );

    \I__6229\ : InMux
    port map (
            O => \N__26395\,
            I => \N__26247\
        );

    \I__6228\ : InMux
    port map (
            O => \N__26394\,
            I => \N__26247\
        );

    \I__6227\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26247\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26235\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__26373\,
            I => \N__26230\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__26364\,
            I => \N__26230\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__26351\,
            I => \N__26227\
        );

    \I__6222\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26210\
        );

    \I__6221\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26210\
        );

    \I__6220\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26210\
        );

    \I__6219\ : InMux
    port map (
            O => \N__26347\,
            I => \N__26210\
        );

    \I__6218\ : InMux
    port map (
            O => \N__26346\,
            I => \N__26210\
        );

    \I__6217\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26210\
        );

    \I__6216\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26210\
        );

    \I__6215\ : InMux
    port map (
            O => \N__26343\,
            I => \N__26210\
        );

    \I__6214\ : Span4Mux_s3_v
    port map (
            O => \N__26340\,
            I => \N__26207\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__26335\,
            I => \N__26204\
        );

    \I__6212\ : Span4Mux_s2_v
    port map (
            O => \N__26332\,
            I => \N__26197\
        );

    \I__6211\ : Span4Mux_s2_h
    port map (
            O => \N__26327\,
            I => \N__26197\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__26312\,
            I => \N__26197\
        );

    \I__6209\ : Span4Mux_s3_v
    port map (
            O => \N__26309\,
            I => \N__26189\
        );

    \I__6208\ : Span4Mux_h
    port map (
            O => \N__26302\,
            I => \N__26184\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26184\
        );

    \I__6206\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26167\
        );

    \I__6205\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26167\
        );

    \I__6204\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26167\
        );

    \I__6203\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26167\
        );

    \I__6202\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26167\
        );

    \I__6201\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26167\
        );

    \I__6200\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26167\
        );

    \I__6199\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26167\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__26264\,
            I => \N__26162\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__26247\,
            I => \N__26162\
        );

    \I__6196\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26159\
        );

    \I__6195\ : InMux
    port map (
            O => \N__26245\,
            I => \N__26142\
        );

    \I__6194\ : InMux
    port map (
            O => \N__26244\,
            I => \N__26142\
        );

    \I__6193\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26142\
        );

    \I__6192\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26142\
        );

    \I__6191\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26142\
        );

    \I__6190\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26142\
        );

    \I__6189\ : InMux
    port map (
            O => \N__26239\,
            I => \N__26142\
        );

    \I__6188\ : InMux
    port map (
            O => \N__26238\,
            I => \N__26142\
        );

    \I__6187\ : Span4Mux_s3_v
    port map (
            O => \N__26235\,
            I => \N__26129\
        );

    \I__6186\ : Span4Mux_s3_h
    port map (
            O => \N__26230\,
            I => \N__26129\
        );

    \I__6185\ : Span4Mux_v
    port map (
            O => \N__26227\,
            I => \N__26129\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__26210\,
            I => \N__26129\
        );

    \I__6183\ : Span4Mux_h
    port map (
            O => \N__26207\,
            I => \N__26129\
        );

    \I__6182\ : Span4Mux_s3_v
    port map (
            O => \N__26204\,
            I => \N__26129\
        );

    \I__6181\ : Span4Mux_h
    port map (
            O => \N__26197\,
            I => \N__26126\
        );

    \I__6180\ : InMux
    port map (
            O => \N__26196\,
            I => \N__26115\
        );

    \I__6179\ : InMux
    port map (
            O => \N__26195\,
            I => \N__26115\
        );

    \I__6178\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26115\
        );

    \I__6177\ : InMux
    port map (
            O => \N__26193\,
            I => \N__26115\
        );

    \I__6176\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26115\
        );

    \I__6175\ : Odrv4
    port map (
            O => \N__26189\,
            I => \A_stk_delta_1\
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__26184\,
            I => \A_stk_delta_1\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__26167\,
            I => \A_stk_delta_1\
        );

    \I__6172\ : Odrv4
    port map (
            O => \N__26162\,
            I => \A_stk_delta_1\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__26159\,
            I => \A_stk_delta_1\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__26142\,
            I => \A_stk_delta_1\
        );

    \I__6169\ : Odrv4
    port map (
            O => \N__26129\,
            I => \A_stk_delta_1\
        );

    \I__6168\ : Odrv4
    port map (
            O => \N__26126\,
            I => \A_stk_delta_1\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__26115\,
            I => \A_stk_delta_1\
        );

    \I__6166\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26093\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26089\
        );

    \I__6164\ : InMux
    port map (
            O => \N__26092\,
            I => \N__26086\
        );

    \I__6163\ : Span12Mux_s5_v
    port map (
            O => \N__26089\,
            I => \N__26083\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__26086\,
            I => \tok.A_stk.tail_51\
        );

    \I__6161\ : Odrv12
    port map (
            O => \N__26083\,
            I => \tok.A_stk.tail_51\
        );

    \I__6160\ : CEMux
    port map (
            O => \N__26078\,
            I => \N__26075\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__26075\,
            I => \N__26068\
        );

    \I__6158\ : CEMux
    port map (
            O => \N__26074\,
            I => \N__26065\
        );

    \I__6157\ : CEMux
    port map (
            O => \N__26073\,
            I => \N__26062\
        );

    \I__6156\ : CEMux
    port map (
            O => \N__26072\,
            I => \N__26050\
        );

    \I__6155\ : CEMux
    port map (
            O => \N__26071\,
            I => \N__26044\
        );

    \I__6154\ : Span4Mux_v
    port map (
            O => \N__26068\,
            I => \N__26039\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__26065\,
            I => \N__26039\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__26062\,
            I => \N__26036\
        );

    \I__6151\ : CEMux
    port map (
            O => \N__26061\,
            I => \N__26032\
        );

    \I__6150\ : CEMux
    port map (
            O => \N__26060\,
            I => \N__26028\
        );

    \I__6149\ : CEMux
    port map (
            O => \N__26059\,
            I => \N__26025\
        );

    \I__6148\ : CEMux
    port map (
            O => \N__26058\,
            I => \N__26022\
        );

    \I__6147\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26016\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__26056\,
            I => \N__26013\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__26055\,
            I => \N__26007\
        );

    \I__6144\ : CascadeMux
    port map (
            O => \N__26054\,
            I => \N__26003\
        );

    \I__6143\ : CascadeMux
    port map (
            O => \N__26053\,
            I => \N__26000\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__26050\,
            I => \N__25996\
        );

    \I__6141\ : CEMux
    port map (
            O => \N__26049\,
            I => \N__25993\
        );

    \I__6140\ : CEMux
    port map (
            O => \N__26048\,
            I => \N__25990\
        );

    \I__6139\ : CEMux
    port map (
            O => \N__26047\,
            I => \N__25987\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__26044\,
            I => \N__25983\
        );

    \I__6137\ : Span4Mux_v
    port map (
            O => \N__26039\,
            I => \N__25978\
        );

    \I__6136\ : Span4Mux_s3_v
    port map (
            O => \N__26036\,
            I => \N__25978\
        );

    \I__6135\ : CEMux
    port map (
            O => \N__26035\,
            I => \N__25975\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__26032\,
            I => \N__25972\
        );

    \I__6133\ : CEMux
    port map (
            O => \N__26031\,
            I => \N__25969\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__26028\,
            I => \N__25965\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__26025\,
            I => \N__25960\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__26022\,
            I => \N__25960\
        );

    \I__6129\ : CEMux
    port map (
            O => \N__26021\,
            I => \N__25957\
        );

    \I__6128\ : CEMux
    port map (
            O => \N__26020\,
            I => \N__25954\
        );

    \I__6127\ : CEMux
    port map (
            O => \N__26019\,
            I => \N__25951\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__26016\,
            I => \N__25948\
        );

    \I__6125\ : InMux
    port map (
            O => \N__26013\,
            I => \N__25943\
        );

    \I__6124\ : InMux
    port map (
            O => \N__26012\,
            I => \N__25943\
        );

    \I__6123\ : InMux
    port map (
            O => \N__26011\,
            I => \N__25928\
        );

    \I__6122\ : InMux
    port map (
            O => \N__26010\,
            I => \N__25928\
        );

    \I__6121\ : InMux
    port map (
            O => \N__26007\,
            I => \N__25928\
        );

    \I__6120\ : InMux
    port map (
            O => \N__26006\,
            I => \N__25928\
        );

    \I__6119\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25928\
        );

    \I__6118\ : InMux
    port map (
            O => \N__26000\,
            I => \N__25928\
        );

    \I__6117\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25928\
        );

    \I__6116\ : Span4Mux_s3_v
    port map (
            O => \N__25996\,
            I => \N__25923\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__25993\,
            I => \N__25918\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__25990\,
            I => \N__25918\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__25987\,
            I => \N__25915\
        );

    \I__6112\ : CEMux
    port map (
            O => \N__25986\,
            I => \N__25912\
        );

    \I__6111\ : Span4Mux_s3_v
    port map (
            O => \N__25983\,
            I => \N__25901\
        );

    \I__6110\ : Span4Mux_s1_h
    port map (
            O => \N__25978\,
            I => \N__25901\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__25975\,
            I => \N__25901\
        );

    \I__6108\ : Span4Mux_s3_v
    port map (
            O => \N__25972\,
            I => \N__25901\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__25969\,
            I => \N__25901\
        );

    \I__6106\ : CEMux
    port map (
            O => \N__25968\,
            I => \N__25898\
        );

    \I__6105\ : Span4Mux_s2_h
    port map (
            O => \N__25965\,
            I => \N__25889\
        );

    \I__6104\ : Span4Mux_v
    port map (
            O => \N__25960\,
            I => \N__25889\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__25957\,
            I => \N__25889\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__25954\,
            I => \N__25889\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__25951\,
            I => \N__25886\
        );

    \I__6100\ : Span4Mux_s3_v
    port map (
            O => \N__25948\,
            I => \N__25883\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__25943\,
            I => \N__25880\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__25928\,
            I => \N__25877\
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__25927\,
            I => \N__25874\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__25926\,
            I => \N__25871\
        );

    \I__6095\ : Span4Mux_h
    port map (
            O => \N__25923\,
            I => \N__25863\
        );

    \I__6094\ : Span4Mux_s3_v
    port map (
            O => \N__25918\,
            I => \N__25863\
        );

    \I__6093\ : Span4Mux_s1_v
    port map (
            O => \N__25915\,
            I => \N__25860\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__25912\,
            I => \N__25853\
        );

    \I__6091\ : Sp12to4
    port map (
            O => \N__25901\,
            I => \N__25853\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__25898\,
            I => \N__25853\
        );

    \I__6089\ : Span4Mux_h
    port map (
            O => \N__25889\,
            I => \N__25850\
        );

    \I__6088\ : Span4Mux_s3_v
    port map (
            O => \N__25886\,
            I => \N__25841\
        );

    \I__6087\ : Span4Mux_h
    port map (
            O => \N__25883\,
            I => \N__25841\
        );

    \I__6086\ : Span4Mux_s3_v
    port map (
            O => \N__25880\,
            I => \N__25841\
        );

    \I__6085\ : Span4Mux_s3_v
    port map (
            O => \N__25877\,
            I => \N__25841\
        );

    \I__6084\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25830\
        );

    \I__6083\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25830\
        );

    \I__6082\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25830\
        );

    \I__6081\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25830\
        );

    \I__6080\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25830\
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__25863\,
            I => \rd_15__N_301\
        );

    \I__6078\ : Odrv4
    port map (
            O => \N__25860\,
            I => \rd_15__N_301\
        );

    \I__6077\ : Odrv12
    port map (
            O => \N__25853\,
            I => \rd_15__N_301\
        );

    \I__6076\ : Odrv4
    port map (
            O => \N__25850\,
            I => \rd_15__N_301\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__25841\,
            I => \rd_15__N_301\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__25830\,
            I => \rd_15__N_301\
        );

    \I__6073\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25814\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__25814\,
            I => \tok.n175\
        );

    \I__6071\ : InMux
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__25808\,
            I => \N__25805\
        );

    \I__6069\ : Span4Mux_s3_h
    port map (
            O => \N__25805\,
            I => \N__25802\
        );

    \I__6068\ : Odrv4
    port map (
            O => \N__25802\,
            I => \tok.n15_adj_770\
        );

    \I__6067\ : InMux
    port map (
            O => \N__25799\,
            I => \N__25796\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__6065\ : Span4Mux_s3_h
    port map (
            O => \N__25793\,
            I => \N__25790\
        );

    \I__6064\ : Span4Mux_v
    port map (
            O => \N__25790\,
            I => \N__25787\
        );

    \I__6063\ : Odrv4
    port map (
            O => \N__25787\,
            I => \tok.n14_adj_769\
        );

    \I__6062\ : CascadeMux
    port map (
            O => \N__25784\,
            I => \tok.n13_adj_772_cascade_\
        );

    \I__6061\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25778\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__25778\,
            I => \tok.n5412\
        );

    \I__6059\ : CascadeMux
    port map (
            O => \N__25775\,
            I => \tok.n22_adj_773_cascade_\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__25772\,
            I => \N__25768\
        );

    \I__6057\ : InMux
    port map (
            O => \N__25771\,
            I => \N__25758\
        );

    \I__6056\ : InMux
    port map (
            O => \N__25768\,
            I => \N__25755\
        );

    \I__6055\ : InMux
    port map (
            O => \N__25767\,
            I => \N__25752\
        );

    \I__6054\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25749\
        );

    \I__6053\ : CascadeMux
    port map (
            O => \N__25765\,
            I => \N__25746\
        );

    \I__6052\ : CascadeMux
    port map (
            O => \N__25764\,
            I => \N__25743\
        );

    \I__6051\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25735\
        );

    \I__6050\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25735\
        );

    \I__6049\ : InMux
    port map (
            O => \N__25761\,
            I => \N__25735\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__25758\,
            I => \N__25732\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__25755\,
            I => \N__25727\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__25752\,
            I => \N__25727\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__25749\,
            I => \N__25724\
        );

    \I__6044\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25721\
        );

    \I__6043\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25716\
        );

    \I__6042\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25716\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__25735\,
            I => \N__25713\
        );

    \I__6040\ : Span4Mux_v
    port map (
            O => \N__25732\,
            I => \N__25708\
        );

    \I__6039\ : Span4Mux_v
    port map (
            O => \N__25727\,
            I => \N__25708\
        );

    \I__6038\ : Span12Mux_s5_h
    port map (
            O => \N__25724\,
            I => \N__25703\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__25721\,
            I => \N__25703\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__25716\,
            I => \tok.A_14\
        );

    \I__6035\ : Odrv4
    port map (
            O => \N__25713\,
            I => \tok.A_14\
        );

    \I__6034\ : Odrv4
    port map (
            O => \N__25708\,
            I => \tok.A_14\
        );

    \I__6033\ : Odrv12
    port map (
            O => \N__25703\,
            I => \tok.A_14\
        );

    \I__6032\ : InMux
    port map (
            O => \N__25694\,
            I => \N__25689\
        );

    \I__6031\ : InMux
    port map (
            O => \N__25693\,
            I => \N__25685\
        );

    \I__6030\ : InMux
    port map (
            O => \N__25692\,
            I => \N__25682\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__25689\,
            I => \N__25676\
        );

    \I__6028\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25673\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__25685\,
            I => \N__25668\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__25682\,
            I => \N__25668\
        );

    \I__6025\ : InMux
    port map (
            O => \N__25681\,
            I => \N__25665\
        );

    \I__6024\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25662\
        );

    \I__6023\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25657\
        );

    \I__6022\ : Span4Mux_v
    port map (
            O => \N__25676\,
            I => \N__25652\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__25673\,
            I => \N__25652\
        );

    \I__6020\ : Span4Mux_h
    port map (
            O => \N__25668\,
            I => \N__25645\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__25665\,
            I => \N__25645\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__25662\,
            I => \N__25645\
        );

    \I__6017\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25642\
        );

    \I__6016\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25639\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__25657\,
            I => \N__25634\
        );

    \I__6014\ : Span4Mux_h
    port map (
            O => \N__25652\,
            I => \N__25634\
        );

    \I__6013\ : Span4Mux_h
    port map (
            O => \N__25645\,
            I => \N__25631\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__25642\,
            I => \N__25628\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__25639\,
            I => \N__25623\
        );

    \I__6010\ : Span4Mux_v
    port map (
            O => \N__25634\,
            I => \N__25623\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__25631\,
            I => \rx_data_7__N_511\
        );

    \I__6008\ : Odrv12
    port map (
            O => \N__25628\,
            I => \rx_data_7__N_511\
        );

    \I__6007\ : Odrv4
    port map (
            O => \N__25623\,
            I => \rx_data_7__N_511\
        );

    \I__6006\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25612\
        );

    \I__6005\ : CascadeMux
    port map (
            O => \N__25615\,
            I => \N__25608\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__25612\,
            I => \N__25605\
        );

    \I__6003\ : InMux
    port map (
            O => \N__25611\,
            I => \N__25600\
        );

    \I__6002\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25600\
        );

    \I__6001\ : Odrv4
    port map (
            O => \N__25605\,
            I => capture_6
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__25600\,
            I => capture_6
        );

    \I__5999\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25589\
        );

    \I__5998\ : InMux
    port map (
            O => \N__25594\,
            I => \N__25589\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__25589\,
            I => \tok.A_stk.tail_11\
        );

    \I__5996\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25580\
        );

    \I__5995\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25580\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__25580\,
            I => \tok.A_stk.tail_27\
        );

    \I__5993\ : InMux
    port map (
            O => \N__25577\,
            I => \N__25571\
        );

    \I__5992\ : InMux
    port map (
            O => \N__25576\,
            I => \N__25571\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__25571\,
            I => \tok.A_stk.tail_43\
        );

    \I__5990\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25565\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__25565\,
            I => \N__25561\
        );

    \I__5988\ : InMux
    port map (
            O => \N__25564\,
            I => \N__25558\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__25561\,
            I => \tok.A_stk.tail_75\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__25558\,
            I => \tok.A_stk.tail_75\
        );

    \I__5985\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25550\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__25550\,
            I => \N__25546\
        );

    \I__5983\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25543\
        );

    \I__5982\ : Span4Mux_h
    port map (
            O => \N__25546\,
            I => \N__25540\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__25543\,
            I => \tok.A_stk.tail_59\
        );

    \I__5980\ : Odrv4
    port map (
            O => \N__25540\,
            I => \tok.A_stk.tail_59\
        );

    \I__5979\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25532\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__25532\,
            I => \tok.n20_adj_648\
        );

    \I__5977\ : CascadeMux
    port map (
            O => \N__25529\,
            I => \N__25526\
        );

    \I__5976\ : InMux
    port map (
            O => \N__25526\,
            I => \N__25523\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__5974\ : Span4Mux_v
    port map (
            O => \N__25520\,
            I => \N__25517\
        );

    \I__5973\ : Odrv4
    port map (
            O => \N__25517\,
            I => \tok.n299\
        );

    \I__5972\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25508\
        );

    \I__5971\ : CascadeMux
    port map (
            O => \N__25513\,
            I => \N__25505\
        );

    \I__5970\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25495\
        );

    \I__5969\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25492\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__25508\,
            I => \N__25489\
        );

    \I__5967\ : InMux
    port map (
            O => \N__25505\,
            I => \N__25484\
        );

    \I__5966\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25484\
        );

    \I__5965\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25479\
        );

    \I__5964\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25479\
        );

    \I__5963\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25474\
        );

    \I__5962\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25474\
        );

    \I__5961\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25468\
        );

    \I__5960\ : InMux
    port map (
            O => \N__25498\,
            I => \N__25468\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__25495\,
            I => \N__25461\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__25492\,
            I => \N__25461\
        );

    \I__5957\ : Span4Mux_v
    port map (
            O => \N__25489\,
            I => \N__25452\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__25484\,
            I => \N__25452\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__25479\,
            I => \N__25452\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__25474\,
            I => \N__25452\
        );

    \I__5953\ : InMux
    port map (
            O => \N__25473\,
            I => \N__25447\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__25468\,
            I => \N__25444\
        );

    \I__5951\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25441\
        );

    \I__5950\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25438\
        );

    \I__5949\ : Span4Mux_s3_v
    port map (
            O => \N__25461\,
            I => \N__25433\
        );

    \I__5948\ : Span4Mux_v
    port map (
            O => \N__25452\,
            I => \N__25433\
        );

    \I__5947\ : InMux
    port map (
            O => \N__25451\,
            I => \N__25430\
        );

    \I__5946\ : InMux
    port map (
            O => \N__25450\,
            I => \N__25427\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__25447\,
            I => \N__25424\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__25444\,
            I => \N__25421\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__25441\,
            I => \N__25418\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__25438\,
            I => \N__25415\
        );

    \I__5941\ : Sp12to4
    port map (
            O => \N__25433\,
            I => \N__25408\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__25430\,
            I => \N__25408\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__25427\,
            I => \N__25408\
        );

    \I__5938\ : Span4Mux_h
    port map (
            O => \N__25424\,
            I => \N__25399\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__25421\,
            I => \N__25399\
        );

    \I__5936\ : Span4Mux_h
    port map (
            O => \N__25418\,
            I => \N__25399\
        );

    \I__5935\ : Span4Mux_s1_v
    port map (
            O => \N__25415\,
            I => \N__25399\
        );

    \I__5934\ : Odrv12
    port map (
            O => \N__25408\,
            I => \tok.n238\
        );

    \I__5933\ : Odrv4
    port map (
            O => \N__25399\,
            I => \tok.n238\
        );

    \I__5932\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__25391\,
            I => \N__25387\
        );

    \I__5930\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25384\
        );

    \I__5929\ : Odrv4
    port map (
            O => \N__25387\,
            I => \tok.A_stk.tail_5\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__25384\,
            I => \tok.A_stk.tail_5\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__5926\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25370\
        );

    \I__5925\ : CascadeMux
    port map (
            O => \N__25375\,
            I => \N__25366\
        );

    \I__5924\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25363\
        );

    \I__5923\ : CascadeMux
    port map (
            O => \N__25373\,
            I => \N__25360\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__25370\,
            I => \N__25357\
        );

    \I__5921\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25354\
        );

    \I__5920\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25351\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__25363\,
            I => \N__25348\
        );

    \I__5918\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25345\
        );

    \I__5917\ : Span4Mux_v
    port map (
            O => \N__25357\,
            I => \N__25340\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__25354\,
            I => \N__25340\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__25351\,
            I => \N__25336\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__25348\,
            I => \N__25330\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__25345\,
            I => \N__25330\
        );

    \I__5912\ : Span4Mux_h
    port map (
            O => \N__25340\,
            I => \N__25325\
        );

    \I__5911\ : InMux
    port map (
            O => \N__25339\,
            I => \N__25322\
        );

    \I__5910\ : Span4Mux_v
    port map (
            O => \N__25336\,
            I => \N__25319\
        );

    \I__5909\ : InMux
    port map (
            O => \N__25335\,
            I => \N__25316\
        );

    \I__5908\ : Span4Mux_h
    port map (
            O => \N__25330\,
            I => \N__25313\
        );

    \I__5907\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25308\
        );

    \I__5906\ : InMux
    port map (
            O => \N__25328\,
            I => \N__25308\
        );

    \I__5905\ : Span4Mux_h
    port map (
            O => \N__25325\,
            I => \N__25303\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25303\
        );

    \I__5903\ : Span4Mux_h
    port map (
            O => \N__25319\,
            I => \N__25298\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__25316\,
            I => \N__25298\
        );

    \I__5901\ : Span4Mux_s1_h
    port map (
            O => \N__25313\,
            I => \N__25295\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__25308\,
            I => \tok.S_3\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__25303\,
            I => \tok.S_3\
        );

    \I__5898\ : Odrv4
    port map (
            O => \N__25298\,
            I => \tok.S_3\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__25295\,
            I => \tok.S_3\
        );

    \I__5896\ : CascadeMux
    port map (
            O => \N__25286\,
            I => \N__25283\
        );

    \I__5895\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25277\
        );

    \I__5894\ : InMux
    port map (
            O => \N__25282\,
            I => \N__25277\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__25277\,
            I => \tok.A_stk.tail_3\
        );

    \I__5892\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25268\
        );

    \I__5891\ : InMux
    port map (
            O => \N__25273\,
            I => \N__25268\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__25268\,
            I => \tok.A_stk.tail_53\
        );

    \I__5889\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25259\
        );

    \I__5888\ : InMux
    port map (
            O => \N__25264\,
            I => \N__25259\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__25259\,
            I => \tok.A_stk.tail_37\
        );

    \I__5886\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25250\
        );

    \I__5885\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25250\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__25250\,
            I => \tok.A_stk.tail_21\
        );

    \I__5883\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25243\
        );

    \I__5882\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25240\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__25243\,
            I => \tok.A_stk.tail_90\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__25240\,
            I => \tok.A_stk.tail_90\
        );

    \I__5879\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25232\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__25232\,
            I => \N__25229\
        );

    \I__5877\ : IoSpan4Mux
    port map (
            O => \N__25229\,
            I => \N__25225\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__25228\,
            I => \N__25222\
        );

    \I__5875\ : Span4Mux_s1_v
    port map (
            O => \N__25225\,
            I => \N__25219\
        );

    \I__5874\ : InMux
    port map (
            O => \N__25222\,
            I => \N__25216\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__25219\,
            I => tail_122
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__25216\,
            I => tail_122
        );

    \I__5871\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25208\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__25208\,
            I => \N__25204\
        );

    \I__5869\ : InMux
    port map (
            O => \N__25207\,
            I => \N__25201\
        );

    \I__5868\ : Span4Mux_h
    port map (
            O => \N__25204\,
            I => \N__25198\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25195\
        );

    \I__5866\ : Odrv4
    port map (
            O => \N__25198\,
            I => tail_106
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__25195\,
            I => tail_106
        );

    \I__5864\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__25187\,
            I => \tok.n23_adj_642\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__25184\,
            I => \N__25181\
        );

    \I__5861\ : InMux
    port map (
            O => \N__25181\,
            I => \N__25178\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__25178\,
            I => \N__25175\
        );

    \I__5859\ : Span4Mux_v
    port map (
            O => \N__25175\,
            I => \N__25172\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__25172\,
            I => \tok.n288\
        );

    \I__5857\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25161\
        );

    \I__5856\ : InMux
    port map (
            O => \N__25168\,
            I => \N__25161\
        );

    \I__5855\ : InMux
    port map (
            O => \N__25167\,
            I => \N__25153\
        );

    \I__5854\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25150\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__25161\,
            I => \N__25147\
        );

    \I__5852\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25142\
        );

    \I__5851\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25139\
        );

    \I__5850\ : InMux
    port map (
            O => \N__25158\,
            I => \N__25136\
        );

    \I__5849\ : InMux
    port map (
            O => \N__25157\,
            I => \N__25131\
        );

    \I__5848\ : InMux
    port map (
            O => \N__25156\,
            I => \N__25131\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__25153\,
            I => \N__25126\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__25150\,
            I => \N__25126\
        );

    \I__5845\ : Span4Mux_v
    port map (
            O => \N__25147\,
            I => \N__25123\
        );

    \I__5844\ : InMux
    port map (
            O => \N__25146\,
            I => \N__25120\
        );

    \I__5843\ : CascadeMux
    port map (
            O => \N__25145\,
            I => \N__25117\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__25142\,
            I => \N__25109\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__25139\,
            I => \N__25109\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__25136\,
            I => \N__25109\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__25131\,
            I => \N__25106\
        );

    \I__5838\ : Span4Mux_s3_v
    port map (
            O => \N__25126\,
            I => \N__25099\
        );

    \I__5837\ : Span4Mux_h
    port map (
            O => \N__25123\,
            I => \N__25099\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__25120\,
            I => \N__25099\
        );

    \I__5835\ : InMux
    port map (
            O => \N__25117\,
            I => \N__25094\
        );

    \I__5834\ : InMux
    port map (
            O => \N__25116\,
            I => \N__25094\
        );

    \I__5833\ : Span4Mux_h
    port map (
            O => \N__25109\,
            I => \N__25091\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__25106\,
            I => \tok.A_11\
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__25099\,
            I => \tok.A_11\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__25094\,
            I => \tok.A_11\
        );

    \I__5829\ : Odrv4
    port map (
            O => \N__25091\,
            I => \tok.A_11\
        );

    \I__5828\ : InMux
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__5826\ : Span4Mux_s1_h
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__5825\ : Span4Mux_h
    port map (
            O => \N__25073\,
            I => \N__25069\
        );

    \I__5824\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25066\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__25069\,
            I => \tok.A_stk.tail_14\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__25066\,
            I => \tok.A_stk.tail_14\
        );

    \I__5821\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25056\
        );

    \I__5820\ : InMux
    port map (
            O => \N__25060\,
            I => \N__25051\
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__25059\,
            I => \N__25048\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__25056\,
            I => \N__25045\
        );

    \I__5817\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25042\
        );

    \I__5816\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25038\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__25051\,
            I => \N__25035\
        );

    \I__5814\ : InMux
    port map (
            O => \N__25048\,
            I => \N__25032\
        );

    \I__5813\ : Span4Mux_h
    port map (
            O => \N__25045\,
            I => \N__25027\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__25042\,
            I => \N__25027\
        );

    \I__5811\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25024\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__25038\,
            I => \N__25021\
        );

    \I__5809\ : Span4Mux_v
    port map (
            O => \N__25035\,
            I => \N__25016\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__25032\,
            I => \N__25016\
        );

    \I__5807\ : Span4Mux_h
    port map (
            O => \N__25027\,
            I => \N__25011\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__25024\,
            I => \N__25011\
        );

    \I__5805\ : Span4Mux_v
    port map (
            O => \N__25021\,
            I => \N__25004\
        );

    \I__5804\ : Span4Mux_h
    port map (
            O => \N__25016\,
            I => \N__25004\
        );

    \I__5803\ : Span4Mux_v
    port map (
            O => \N__25011\,
            I => \N__25001\
        );

    \I__5802\ : InMux
    port map (
            O => \N__25010\,
            I => \N__24996\
        );

    \I__5801\ : InMux
    port map (
            O => \N__25009\,
            I => \N__24996\
        );

    \I__5800\ : Span4Mux_h
    port map (
            O => \N__25004\,
            I => \N__24993\
        );

    \I__5799\ : Odrv4
    port map (
            O => \N__25001\,
            I => \tok.S_11\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__24996\,
            I => \tok.S_11\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__24993\,
            I => \tok.S_11\
        );

    \I__5796\ : CascadeMux
    port map (
            O => \N__24986\,
            I => \N__24983\
        );

    \I__5795\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24977\
        );

    \I__5794\ : InMux
    port map (
            O => \N__24982\,
            I => \N__24977\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__24977\,
            I => \tok.A_stk.tail_74\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__24974\,
            I => \N__24971\
        );

    \I__5791\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24965\
        );

    \I__5790\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24965\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__24965\,
            I => \tok.A_stk.tail_58\
        );

    \I__5788\ : InMux
    port map (
            O => \N__24962\,
            I => \N__24956\
        );

    \I__5787\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24956\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__24956\,
            I => \tok.A_stk.tail_42\
        );

    \I__5785\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24947\
        );

    \I__5784\ : InMux
    port map (
            O => \N__24952\,
            I => \N__24947\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__24947\,
            I => \tok.A_stk.tail_26\
        );

    \I__5782\ : CascadeMux
    port map (
            O => \N__24944\,
            I => \N__24941\
        );

    \I__5781\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24935\
        );

    \I__5780\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24935\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__24935\,
            I => \tok.A_stk.tail_10\
        );

    \I__5778\ : InMux
    port map (
            O => \N__24932\,
            I => \N__24929\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__24929\,
            I => \N__24926\
        );

    \I__5776\ : Span4Mux_s2_h
    port map (
            O => \N__24926\,
            I => \N__24922\
        );

    \I__5775\ : InMux
    port map (
            O => \N__24925\,
            I => \N__24919\
        );

    \I__5774\ : Odrv4
    port map (
            O => \N__24922\,
            I => tail_117
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__24919\,
            I => tail_117
        );

    \I__5772\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24911\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__24911\,
            I => \N__24908\
        );

    \I__5770\ : Span4Mux_h
    port map (
            O => \N__24908\,
            I => \N__24905\
        );

    \I__5769\ : Span4Mux_h
    port map (
            O => \N__24905\,
            I => \N__24901\
        );

    \I__5768\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24898\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__24901\,
            I => tail_101
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__24898\,
            I => tail_101
        );

    \I__5765\ : InMux
    port map (
            O => \N__24893\,
            I => \N__24889\
        );

    \I__5764\ : InMux
    port map (
            O => \N__24892\,
            I => \N__24886\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__24889\,
            I => \tok.A_stk.tail_85\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__24886\,
            I => \tok.A_stk.tail_85\
        );

    \I__5761\ : InMux
    port map (
            O => \N__24881\,
            I => \N__24875\
        );

    \I__5760\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24875\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__24875\,
            I => \tok.A_stk.tail_69\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__24872\,
            I => \N__24869\
        );

    \I__5757\ : InMux
    port map (
            O => \N__24869\,
            I => \N__24866\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__24866\,
            I => \tok.n287\
        );

    \I__5755\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24857\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__24862\,
            I => \N__24854\
        );

    \I__5753\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24851\
        );

    \I__5752\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24848\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__24857\,
            I => \N__24840\
        );

    \I__5750\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24837\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__24851\,
            I => \N__24834\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__24848\,
            I => \N__24831\
        );

    \I__5747\ : InMux
    port map (
            O => \N__24847\,
            I => \N__24826\
        );

    \I__5746\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24826\
        );

    \I__5745\ : CascadeMux
    port map (
            O => \N__24845\,
            I => \N__24822\
        );

    \I__5744\ : CascadeMux
    port map (
            O => \N__24844\,
            I => \N__24819\
        );

    \I__5743\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24816\
        );

    \I__5742\ : Span4Mux_h
    port map (
            O => \N__24840\,
            I => \N__24811\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__24837\,
            I => \N__24811\
        );

    \I__5740\ : Span4Mux_h
    port map (
            O => \N__24834\,
            I => \N__24804\
        );

    \I__5739\ : Span4Mux_v
    port map (
            O => \N__24831\,
            I => \N__24804\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24804\
        );

    \I__5737\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24801\
        );

    \I__5736\ : InMux
    port map (
            O => \N__24822\,
            I => \N__24796\
        );

    \I__5735\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24796\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__24816\,
            I => \N__24791\
        );

    \I__5733\ : Span4Mux_h
    port map (
            O => \N__24811\,
            I => \N__24791\
        );

    \I__5732\ : Odrv4
    port map (
            O => \N__24804\,
            I => \tok.A_15\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__24801\,
            I => \tok.A_15\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__24796\,
            I => \tok.A_15\
        );

    \I__5729\ : Odrv4
    port map (
            O => \N__24791\,
            I => \tok.A_15\
        );

    \I__5728\ : CascadeMux
    port map (
            O => \N__24782\,
            I => \N__24779\
        );

    \I__5727\ : InMux
    port map (
            O => \N__24779\,
            I => \N__24774\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__24778\,
            I => \N__24771\
        );

    \I__5725\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24768\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__24774\,
            I => \N__24764\
        );

    \I__5723\ : InMux
    port map (
            O => \N__24771\,
            I => \N__24761\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__24768\,
            I => \N__24755\
        );

    \I__5721\ : InMux
    port map (
            O => \N__24767\,
            I => \N__24752\
        );

    \I__5720\ : Span4Mux_h
    port map (
            O => \N__24764\,
            I => \N__24747\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__24761\,
            I => \N__24747\
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__24760\,
            I => \N__24743\
        );

    \I__5717\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24738\
        );

    \I__5716\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24738\
        );

    \I__5715\ : Span4Mux_h
    port map (
            O => \N__24755\,
            I => \N__24735\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__24752\,
            I => \N__24732\
        );

    \I__5713\ : Span4Mux_h
    port map (
            O => \N__24747\,
            I => \N__24729\
        );

    \I__5712\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24724\
        );

    \I__5711\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24724\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__24738\,
            I => \N__24719\
        );

    \I__5709\ : Span4Mux_v
    port map (
            O => \N__24735\,
            I => \N__24719\
        );

    \I__5708\ : Span4Mux_h
    port map (
            O => \N__24732\,
            I => \N__24714\
        );

    \I__5707\ : Span4Mux_s1_h
    port map (
            O => \N__24729\,
            I => \N__24714\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__24724\,
            I => \N__24711\
        );

    \I__5705\ : Odrv4
    port map (
            O => \N__24719\,
            I => \tok.S_15\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__24714\,
            I => \tok.S_15\
        );

    \I__5703\ : Odrv12
    port map (
            O => \N__24711\,
            I => \tok.S_15\
        );

    \I__5702\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24698\
        );

    \I__5701\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24698\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__24698\,
            I => \tok.A_stk.tail_15\
        );

    \I__5699\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24689\
        );

    \I__5698\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24689\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__24689\,
            I => \tok.A_stk.tail_31\
        );

    \I__5696\ : InMux
    port map (
            O => \N__24686\,
            I => \N__24680\
        );

    \I__5695\ : InMux
    port map (
            O => \N__24685\,
            I => \N__24680\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__24680\,
            I => \tok.A_stk.tail_47\
        );

    \I__5693\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24674\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__24674\,
            I => \N__24671\
        );

    \I__5691\ : Span4Mux_v
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__24668\,
            I => \N__24664\
        );

    \I__5689\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24661\
        );

    \I__5688\ : Span4Mux_h
    port map (
            O => \N__24664\,
            I => \N__24658\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__24661\,
            I => \N__24655\
        );

    \I__5686\ : Odrv4
    port map (
            O => \N__24658\,
            I => \tok.A_stk.tail_95\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__24655\,
            I => \tok.A_stk.tail_95\
        );

    \I__5684\ : InMux
    port map (
            O => \N__24650\,
            I => \N__24644\
        );

    \I__5683\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24644\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__24644\,
            I => \tok.A_stk.tail_63\
        );

    \I__5681\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__24638\,
            I => \N__24635\
        );

    \I__5679\ : Span4Mux_h
    port map (
            O => \N__24635\,
            I => \N__24631\
        );

    \I__5678\ : InMux
    port map (
            O => \N__24634\,
            I => \N__24628\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__24631\,
            I => \N__24625\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__24628\,
            I => \tok.A_stk.tail_79\
        );

    \I__5675\ : Odrv4
    port map (
            O => \N__24625\,
            I => \tok.A_stk.tail_79\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__5673\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24614\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__24614\,
            I => \N__24611\
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__24611\,
            I => \tok.n293\
        );

    \I__5670\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__24605\,
            I => \N__24602\
        );

    \I__5668\ : Span4Mux_v
    port map (
            O => \N__24602\,
            I => \N__24599\
        );

    \I__5667\ : Odrv4
    port map (
            O => \N__24599\,
            I => \tok.n28\
        );

    \I__5666\ : InMux
    port map (
            O => \N__24596\,
            I => \tok.n4777\
        );

    \I__5665\ : InMux
    port map (
            O => \N__24593\,
            I => \N__24585\
        );

    \I__5664\ : InMux
    port map (
            O => \N__24592\,
            I => \N__24580\
        );

    \I__5663\ : InMux
    port map (
            O => \N__24591\,
            I => \N__24580\
        );

    \I__5662\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24577\
        );

    \I__5661\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24572\
        );

    \I__5660\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24572\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24567\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__24580\,
            I => \N__24567\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__24577\,
            I => \N__24562\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__24572\,
            I => \N__24562\
        );

    \I__5655\ : Span4Mux_v
    port map (
            O => \N__24567\,
            I => \N__24559\
        );

    \I__5654\ : Span4Mux_v
    port map (
            O => \N__24562\,
            I => \N__24556\
        );

    \I__5653\ : Span4Mux_h
    port map (
            O => \N__24559\,
            I => \N__24551\
        );

    \I__5652\ : Span4Mux_h
    port map (
            O => \N__24556\,
            I => \N__24551\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__24551\,
            I => \tok.n8_adj_792\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__24548\,
            I => \N__24545\
        );

    \I__5649\ : InMux
    port map (
            O => \N__24545\,
            I => \N__24542\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__5647\ : Odrv12
    port map (
            O => \N__24539\,
            I => \tok.n292\
        );

    \I__5646\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24533\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__5644\ : Odrv4
    port map (
            O => \N__24530\,
            I => \tok.n27_adj_704\
        );

    \I__5643\ : InMux
    port map (
            O => \N__24527\,
            I => \tok.n4778\
        );

    \I__5642\ : CascadeMux
    port map (
            O => \N__24524\,
            I => \N__24521\
        );

    \I__5641\ : InMux
    port map (
            O => \N__24521\,
            I => \N__24518\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__5639\ : Span4Mux_s2_h
    port map (
            O => \N__24515\,
            I => \N__24512\
        );

    \I__5638\ : Odrv4
    port map (
            O => \N__24512\,
            I => \tok.n291\
        );

    \I__5637\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24506\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24503\
        );

    \I__5635\ : Odrv12
    port map (
            O => \N__24503\,
            I => \tok.n6_adj_728\
        );

    \I__5634\ : InMux
    port map (
            O => \N__24500\,
            I => \tok.n4779\
        );

    \I__5633\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24494\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__24494\,
            I => \N__24491\
        );

    \I__5631\ : Odrv12
    port map (
            O => \N__24491\,
            I => \tok.n290\
        );

    \I__5630\ : CascadeMux
    port map (
            O => \N__24488\,
            I => \N__24485\
        );

    \I__5629\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__24482\,
            I => \N__24474\
        );

    \I__5627\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24471\
        );

    \I__5626\ : InMux
    port map (
            O => \N__24480\,
            I => \N__24468\
        );

    \I__5625\ : InMux
    port map (
            O => \N__24479\,
            I => \N__24465\
        );

    \I__5624\ : CascadeMux
    port map (
            O => \N__24478\,
            I => \N__24461\
        );

    \I__5623\ : CascadeMux
    port map (
            O => \N__24477\,
            I => \N__24458\
        );

    \I__5622\ : Span4Mux_h
    port map (
            O => \N__24474\,
            I => \N__24452\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__24471\,
            I => \N__24452\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__24468\,
            I => \N__24447\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__24465\,
            I => \N__24447\
        );

    \I__5618\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24444\
        );

    \I__5617\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24441\
        );

    \I__5616\ : InMux
    port map (
            O => \N__24458\,
            I => \N__24438\
        );

    \I__5615\ : InMux
    port map (
            O => \N__24457\,
            I => \N__24435\
        );

    \I__5614\ : Span4Mux_v
    port map (
            O => \N__24452\,
            I => \N__24432\
        );

    \I__5613\ : Span4Mux_v
    port map (
            O => \N__24447\,
            I => \N__24427\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__24444\,
            I => \N__24427\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__24441\,
            I => \N__24424\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__24438\,
            I => \N__24421\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__24435\,
            I => \N__24414\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__24432\,
            I => \N__24414\
        );

    \I__5607\ : Span4Mux_v
    port map (
            O => \N__24427\,
            I => \N__24414\
        );

    \I__5606\ : Span4Mux_v
    port map (
            O => \N__24424\,
            I => \N__24409\
        );

    \I__5605\ : Span4Mux_h
    port map (
            O => \N__24421\,
            I => \N__24409\
        );

    \I__5604\ : Odrv4
    port map (
            O => \N__24414\,
            I => \tok.S_12\
        );

    \I__5603\ : Odrv4
    port map (
            O => \N__24409\,
            I => \tok.S_12\
        );

    \I__5602\ : InMux
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__24401\,
            I => \N__24398\
        );

    \I__5600\ : Span4Mux_v
    port map (
            O => \N__24398\,
            I => \N__24395\
        );

    \I__5599\ : Odrv4
    port map (
            O => \N__24395\,
            I => \tok.n6_adj_742\
        );

    \I__5598\ : InMux
    port map (
            O => \N__24392\,
            I => \tok.n4780\
        );

    \I__5597\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24386\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__24386\,
            I => \N__24383\
        );

    \I__5595\ : Span4Mux_s3_h
    port map (
            O => \N__24383\,
            I => \N__24380\
        );

    \I__5594\ : Span4Mux_h
    port map (
            O => \N__24380\,
            I => \N__24377\
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__24377\,
            I => \tok.n289\
        );

    \I__5592\ : CascadeMux
    port map (
            O => \N__24374\,
            I => \N__24371\
        );

    \I__5591\ : InMux
    port map (
            O => \N__24371\,
            I => \N__24366\
        );

    \I__5590\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24361\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__24369\,
            I => \N__24358\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__24366\,
            I => \N__24355\
        );

    \I__5587\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24352\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__24364\,
            I => \N__24348\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__24361\,
            I => \N__24345\
        );

    \I__5584\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24342\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__24355\,
            I => \N__24338\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__24352\,
            I => \N__24335\
        );

    \I__5581\ : InMux
    port map (
            O => \N__24351\,
            I => \N__24332\
        );

    \I__5580\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24329\
        );

    \I__5579\ : Span4Mux_h
    port map (
            O => \N__24345\,
            I => \N__24326\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__24342\,
            I => \N__24323\
        );

    \I__5577\ : CascadeMux
    port map (
            O => \N__24341\,
            I => \N__24320\
        );

    \I__5576\ : Span4Mux_v
    port map (
            O => \N__24338\,
            I => \N__24314\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__24335\,
            I => \N__24314\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__24332\,
            I => \N__24311\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24308\
        );

    \I__5572\ : Span4Mux_v
    port map (
            O => \N__24326\,
            I => \N__24303\
        );

    \I__5571\ : Span4Mux_h
    port map (
            O => \N__24323\,
            I => \N__24303\
        );

    \I__5570\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24300\
        );

    \I__5569\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24297\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__24314\,
            I => \N__24294\
        );

    \I__5567\ : Span12Mux_s11_h
    port map (
            O => \N__24311\,
            I => \N__24285\
        );

    \I__5566\ : Span12Mux_s5_v
    port map (
            O => \N__24308\,
            I => \N__24285\
        );

    \I__5565\ : Sp12to4
    port map (
            O => \N__24303\,
            I => \N__24285\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__24300\,
            I => \N__24285\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__24297\,
            I => \tok.S_13\
        );

    \I__5562\ : Odrv4
    port map (
            O => \N__24294\,
            I => \tok.S_13\
        );

    \I__5561\ : Odrv12
    port map (
            O => \N__24285\,
            I => \tok.S_13\
        );

    \I__5560\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24275\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__24275\,
            I => \N__24272\
        );

    \I__5558\ : Span4Mux_h
    port map (
            O => \N__24272\,
            I => \N__24269\
        );

    \I__5557\ : Odrv4
    port map (
            O => \N__24269\,
            I => \tok.n6_adj_752\
        );

    \I__5556\ : InMux
    port map (
            O => \N__24266\,
            I => \tok.n4781\
        );

    \I__5555\ : InMux
    port map (
            O => \N__24263\,
            I => \tok.n4782\
        );

    \I__5554\ : SRMux
    port map (
            O => \N__24260\,
            I => \N__24255\
        );

    \I__5553\ : DummyBuf
    port map (
            O => \N__24259\,
            I => \N__24251\
        );

    \I__5552\ : DummyBuf
    port map (
            O => \N__24258\,
            I => \N__24248\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__24255\,
            I => \N__24244\
        );

    \I__5550\ : SRMux
    port map (
            O => \N__24254\,
            I => \N__24241\
        );

    \I__5549\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24238\
        );

    \I__5548\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24235\
        );

    \I__5547\ : SRMux
    port map (
            O => \N__24247\,
            I => \N__24232\
        );

    \I__5546\ : Span4Mux_v
    port map (
            O => \N__24244\,
            I => \N__24227\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__24241\,
            I => \N__24227\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__24238\,
            I => \N__24221\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__24235\,
            I => \N__24221\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24216\
        );

    \I__5541\ : Span4Mux_h
    port map (
            O => \N__24227\,
            I => \N__24213\
        );

    \I__5540\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24210\
        );

    \I__5539\ : Span4Mux_h
    port map (
            O => \N__24221\,
            I => \N__24206\
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__24220\,
            I => \N__24203\
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__24219\,
            I => \N__24200\
        );

    \I__5536\ : Span4Mux_h
    port map (
            O => \N__24216\,
            I => \N__24197\
        );

    \I__5535\ : Span4Mux_v
    port map (
            O => \N__24213\,
            I => \N__24194\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__24210\,
            I => \N__24191\
        );

    \I__5533\ : CascadeMux
    port map (
            O => \N__24209\,
            I => \N__24186\
        );

    \I__5532\ : Sp12to4
    port map (
            O => \N__24206\,
            I => \N__24183\
        );

    \I__5531\ : InMux
    port map (
            O => \N__24203\,
            I => \N__24178\
        );

    \I__5530\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24178\
        );

    \I__5529\ : Span4Mux_h
    port map (
            O => \N__24197\,
            I => \N__24175\
        );

    \I__5528\ : Span4Mux_s1_v
    port map (
            O => \N__24194\,
            I => \N__24170\
        );

    \I__5527\ : Span4Mux_v
    port map (
            O => \N__24191\,
            I => \N__24170\
        );

    \I__5526\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24167\
        );

    \I__5525\ : InMux
    port map (
            O => \N__24189\,
            I => \N__24164\
        );

    \I__5524\ : InMux
    port map (
            O => \N__24186\,
            I => \N__24161\
        );

    \I__5523\ : Span12Mux_v
    port map (
            O => \N__24183\,
            I => \N__24156\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__24178\,
            I => \N__24156\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__24175\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5520\ : Odrv4
    port map (
            O => \N__24170\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__24167\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__24164\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__24161\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5516\ : Odrv12
    port map (
            O => \N__24156\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5515\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24131\
        );

    \I__5514\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24126\
        );

    \I__5513\ : InMux
    port map (
            O => \N__24141\,
            I => \N__24126\
        );

    \I__5512\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24119\
        );

    \I__5511\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24119\
        );

    \I__5510\ : InMux
    port map (
            O => \N__24138\,
            I => \N__24119\
        );

    \I__5509\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24114\
        );

    \I__5508\ : InMux
    port map (
            O => \N__24136\,
            I => \N__24114\
        );

    \I__5507\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24109\
        );

    \I__5506\ : InMux
    port map (
            O => \N__24134\,
            I => \N__24109\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__24131\,
            I => \N__24106\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__24126\,
            I => \N__24103\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__24119\,
            I => \N__24098\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__24114\,
            I => \N__24098\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__24109\,
            I => \N__24095\
        );

    \I__5500\ : Span4Mux_v
    port map (
            O => \N__24106\,
            I => \N__24090\
        );

    \I__5499\ : Span4Mux_v
    port map (
            O => \N__24103\,
            I => \N__24090\
        );

    \I__5498\ : Span4Mux_s3_h
    port map (
            O => \N__24098\,
            I => \N__24087\
        );

    \I__5497\ : Sp12to4
    port map (
            O => \N__24095\,
            I => \N__24082\
        );

    \I__5496\ : Sp12to4
    port map (
            O => \N__24090\,
            I => \N__24082\
        );

    \I__5495\ : Span4Mux_h
    port map (
            O => \N__24087\,
            I => \N__24079\
        );

    \I__5494\ : Odrv12
    port map (
            O => \N__24082\,
            I => \tok.n400\
        );

    \I__5493\ : Odrv4
    port map (
            O => \N__24079\,
            I => \tok.n400\
        );

    \I__5492\ : InMux
    port map (
            O => \N__24074\,
            I => \bfn_11_11_0_\
        );

    \I__5491\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24068\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__24065\
        );

    \I__5489\ : Span4Mux_h
    port map (
            O => \N__24065\,
            I => \N__24062\
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__24062\,
            I => \tok.n6_adj_783\
        );

    \I__5487\ : InMux
    port map (
            O => \N__24059\,
            I => \N__24056\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__24056\,
            I => \N__24053\
        );

    \I__5485\ : Odrv12
    port map (
            O => \N__24053\,
            I => \tok.n301\
        );

    \I__5484\ : CascadeMux
    port map (
            O => \N__24050\,
            I => \N__24047\
        );

    \I__5483\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24044\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__24044\,
            I => \N__24040\
        );

    \I__5481\ : CascadeMux
    port map (
            O => \N__24043\,
            I => \N__24036\
        );

    \I__5480\ : Span4Mux_v
    port map (
            O => \N__24040\,
            I => \N__24032\
        );

    \I__5479\ : InMux
    port map (
            O => \N__24039\,
            I => \N__24025\
        );

    \I__5478\ : InMux
    port map (
            O => \N__24036\,
            I => \N__24022\
        );

    \I__5477\ : CascadeMux
    port map (
            O => \N__24035\,
            I => \N__24019\
        );

    \I__5476\ : Span4Mux_s3_h
    port map (
            O => \N__24032\,
            I => \N__24016\
        );

    \I__5475\ : InMux
    port map (
            O => \N__24031\,
            I => \N__24011\
        );

    \I__5474\ : InMux
    port map (
            O => \N__24030\,
            I => \N__24011\
        );

    \I__5473\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24008\
        );

    \I__5472\ : CascadeMux
    port map (
            O => \N__24028\,
            I => \N__24005\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__24025\,
            I => \N__24000\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__24022\,
            I => \N__24000\
        );

    \I__5469\ : InMux
    port map (
            O => \N__24019\,
            I => \N__23997\
        );

    \I__5468\ : Span4Mux_h
    port map (
            O => \N__24016\,
            I => \N__23992\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__23992\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__24008\,
            I => \N__23989\
        );

    \I__5465\ : InMux
    port map (
            O => \N__24005\,
            I => \N__23986\
        );

    \I__5464\ : Span4Mux_h
    port map (
            O => \N__24000\,
            I => \N__23981\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__23997\,
            I => \N__23981\
        );

    \I__5462\ : Span4Mux_v
    port map (
            O => \N__23992\,
            I => \N__23975\
        );

    \I__5461\ : Span4Mux_h
    port map (
            O => \N__23989\,
            I => \N__23975\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__23986\,
            I => \N__23972\
        );

    \I__5459\ : Span4Mux_v
    port map (
            O => \N__23981\,
            I => \N__23969\
        );

    \I__5458\ : InMux
    port map (
            O => \N__23980\,
            I => \N__23966\
        );

    \I__5457\ : Span4Mux_v
    port map (
            O => \N__23975\,
            I => \N__23963\
        );

    \I__5456\ : Span4Mux_v
    port map (
            O => \N__23972\,
            I => \N__23958\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__23969\,
            I => \N__23958\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__23966\,
            I => \tok.S_1\
        );

    \I__5453\ : Odrv4
    port map (
            O => \N__23963\,
            I => \tok.S_1\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__23958\,
            I => \tok.S_1\
        );

    \I__5451\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__23948\,
            I => \N__23945\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__23945\,
            I => \tok.n20_adj_799\
        );

    \I__5448\ : InMux
    port map (
            O => \N__23942\,
            I => \tok.n4769\
        );

    \I__5447\ : CascadeMux
    port map (
            O => \N__23939\,
            I => \N__23936\
        );

    \I__5446\ : InMux
    port map (
            O => \N__23936\,
            I => \N__23933\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__23933\,
            I => \N__23928\
        );

    \I__5444\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23925\
        );

    \I__5443\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23921\
        );

    \I__5442\ : Span4Mux_h
    port map (
            O => \N__23928\,
            I => \N__23917\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__23925\,
            I => \N__23914\
        );

    \I__5440\ : InMux
    port map (
            O => \N__23924\,
            I => \N__23910\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__23921\,
            I => \N__23907\
        );

    \I__5438\ : CascadeMux
    port map (
            O => \N__23920\,
            I => \N__23903\
        );

    \I__5437\ : Span4Mux_h
    port map (
            O => \N__23917\,
            I => \N__23900\
        );

    \I__5436\ : Span4Mux_h
    port map (
            O => \N__23914\,
            I => \N__23897\
        );

    \I__5435\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23894\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__23910\,
            I => \N__23891\
        );

    \I__5433\ : Span4Mux_s3_v
    port map (
            O => \N__23907\,
            I => \N__23888\
        );

    \I__5432\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23885\
        );

    \I__5431\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23882\
        );

    \I__5430\ : Span4Mux_v
    port map (
            O => \N__23900\,
            I => \N__23873\
        );

    \I__5429\ : Span4Mux_h
    port map (
            O => \N__23897\,
            I => \N__23873\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__23894\,
            I => \N__23873\
        );

    \I__5427\ : Span4Mux_v
    port map (
            O => \N__23891\,
            I => \N__23870\
        );

    \I__5426\ : Span4Mux_h
    port map (
            O => \N__23888\,
            I => \N__23865\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__23885\,
            I => \N__23865\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__23882\,
            I => \N__23862\
        );

    \I__5423\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23857\
        );

    \I__5422\ : InMux
    port map (
            O => \N__23880\,
            I => \N__23857\
        );

    \I__5421\ : Span4Mux_v
    port map (
            O => \N__23873\,
            I => \N__23854\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__23870\,
            I => \N__23847\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__23865\,
            I => \N__23847\
        );

    \I__5418\ : Span4Mux_h
    port map (
            O => \N__23862\,
            I => \N__23847\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__23857\,
            I => \tok.S_2\
        );

    \I__5416\ : Odrv4
    port map (
            O => \N__23854\,
            I => \tok.S_2\
        );

    \I__5415\ : Odrv4
    port map (
            O => \N__23847\,
            I => \tok.S_2\
        );

    \I__5414\ : CascadeMux
    port map (
            O => \N__23840\,
            I => \N__23837\
        );

    \I__5413\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23834\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__23834\,
            I => \N__23831\
        );

    \I__5411\ : Span4Mux_s3_h
    port map (
            O => \N__23831\,
            I => \N__23828\
        );

    \I__5410\ : Odrv4
    port map (
            O => \N__23828\,
            I => \tok.n300\
        );

    \I__5409\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23822\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__23822\,
            I => \N__23819\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__23819\,
            I => \tok.n22_adj_797\
        );

    \I__5406\ : InMux
    port map (
            O => \N__23816\,
            I => \tok.n4770\
        );

    \I__5405\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23810\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__23810\,
            I => \N__23807\
        );

    \I__5403\ : Span4Mux_h
    port map (
            O => \N__23807\,
            I => \N__23804\
        );

    \I__5402\ : Span4Mux_h
    port map (
            O => \N__23804\,
            I => \N__23801\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__23801\,
            I => \tok.n10_adj_791\
        );

    \I__5400\ : InMux
    port map (
            O => \N__23798\,
            I => \tok.n4771\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__23795\,
            I => \N__23789\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__23794\,
            I => \N__23786\
        );

    \I__5397\ : InMux
    port map (
            O => \N__23793\,
            I => \N__23783\
        );

    \I__5396\ : CascadeMux
    port map (
            O => \N__23792\,
            I => \N__23780\
        );

    \I__5395\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23777\
        );

    \I__5394\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23772\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__23783\,
            I => \N__23769\
        );

    \I__5392\ : InMux
    port map (
            O => \N__23780\,
            I => \N__23766\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__23777\,
            I => \N__23763\
        );

    \I__5390\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23759\
        );

    \I__5389\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23756\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__23772\,
            I => \N__23749\
        );

    \I__5387\ : Span4Mux_v
    port map (
            O => \N__23769\,
            I => \N__23749\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__23766\,
            I => \N__23749\
        );

    \I__5385\ : Span4Mux_h
    port map (
            O => \N__23763\,
            I => \N__23746\
        );

    \I__5384\ : CascadeMux
    port map (
            O => \N__23762\,
            I => \N__23743\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__23759\,
            I => \N__23739\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__23756\,
            I => \N__23736\
        );

    \I__5381\ : Span4Mux_h
    port map (
            O => \N__23749\,
            I => \N__23733\
        );

    \I__5380\ : Span4Mux_h
    port map (
            O => \N__23746\,
            I => \N__23729\
        );

    \I__5379\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23726\
        );

    \I__5378\ : InMux
    port map (
            O => \N__23742\,
            I => \N__23723\
        );

    \I__5377\ : Span4Mux_v
    port map (
            O => \N__23739\,
            I => \N__23718\
        );

    \I__5376\ : Span4Mux_v
    port map (
            O => \N__23736\,
            I => \N__23718\
        );

    \I__5375\ : Span4Mux_v
    port map (
            O => \N__23733\,
            I => \N__23715\
        );

    \I__5374\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23712\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__23729\,
            I => \N__23707\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__23726\,
            I => \N__23707\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__23723\,
            I => \tok.S_4\
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__23718\,
            I => \tok.S_4\
        );

    \I__5369\ : Odrv4
    port map (
            O => \N__23715\,
            I => \tok.S_4\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__23712\,
            I => \tok.S_4\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__23707\,
            I => \tok.S_4\
        );

    \I__5366\ : InMux
    port map (
            O => \N__23696\,
            I => \N__23693\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__23693\,
            I => \N__23690\
        );

    \I__5364\ : Span4Mux_h
    port map (
            O => \N__23690\,
            I => \N__23687\
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__23687\,
            I => \tok.n6_adj_762\
        );

    \I__5362\ : InMux
    port map (
            O => \N__23684\,
            I => \tok.n4772\
        );

    \I__5361\ : InMux
    port map (
            O => \N__23681\,
            I => \tok.n4773\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__23678\,
            I => \N__23674\
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__23677\,
            I => \N__23671\
        );

    \I__5358\ : InMux
    port map (
            O => \N__23674\,
            I => \N__23668\
        );

    \I__5357\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23661\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__23668\,
            I => \N__23658\
        );

    \I__5355\ : InMux
    port map (
            O => \N__23667\,
            I => \N__23655\
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__23666\,
            I => \N__23652\
        );

    \I__5353\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23649\
        );

    \I__5352\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23645\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__23661\,
            I => \N__23642\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__23658\,
            I => \N__23637\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__23655\,
            I => \N__23637\
        );

    \I__5348\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23634\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__23649\,
            I => \N__23630\
        );

    \I__5346\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23626\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__23645\,
            I => \N__23623\
        );

    \I__5344\ : Span4Mux_v
    port map (
            O => \N__23642\,
            I => \N__23620\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__23637\,
            I => \N__23615\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__23634\,
            I => \N__23615\
        );

    \I__5341\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23612\
        );

    \I__5340\ : Span4Mux_h
    port map (
            O => \N__23630\,
            I => \N__23609\
        );

    \I__5339\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23606\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__23626\,
            I => \N__23597\
        );

    \I__5337\ : Span4Mux_v
    port map (
            O => \N__23623\,
            I => \N__23597\
        );

    \I__5336\ : Span4Mux_s1_h
    port map (
            O => \N__23620\,
            I => \N__23597\
        );

    \I__5335\ : Span4Mux_v
    port map (
            O => \N__23615\,
            I => \N__23597\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__23612\,
            I => \tok.S_6\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__23609\,
            I => \tok.S_6\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__23606\,
            I => \tok.S_6\
        );

    \I__5331\ : Odrv4
    port map (
            O => \N__23597\,
            I => \tok.S_6\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__23588\,
            I => \N__23585\
        );

    \I__5329\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__23582\,
            I => \N__23579\
        );

    \I__5327\ : Span4Mux_v
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__5326\ : Odrv4
    port map (
            O => \N__23576\,
            I => \tok.n296\
        );

    \I__5325\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__23567\,
            I => \N__23564\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__23564\,
            I => \tok.n6\
        );

    \I__5321\ : InMux
    port map (
            O => \N__23561\,
            I => \tok.n4774\
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__23558\,
            I => \N__23555\
        );

    \I__5319\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23550\
        );

    \I__5318\ : CascadeMux
    port map (
            O => \N__23554\,
            I => \N__23547\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__23553\,
            I => \N__23544\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__23550\,
            I => \N__23540\
        );

    \I__5315\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23537\
        );

    \I__5314\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23534\
        );

    \I__5313\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23530\
        );

    \I__5312\ : Span4Mux_s3_v
    port map (
            O => \N__23540\,
            I => \N__23527\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__23537\,
            I => \N__23524\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23520\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__23533\,
            I => \N__23516\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__23530\,
            I => \N__23513\
        );

    \I__5307\ : Span4Mux_h
    port map (
            O => \N__23527\,
            I => \N__23508\
        );

    \I__5306\ : Span4Mux_s3_v
    port map (
            O => \N__23524\,
            I => \N__23508\
        );

    \I__5305\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23503\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__23520\,
            I => \N__23500\
        );

    \I__5303\ : InMux
    port map (
            O => \N__23519\,
            I => \N__23497\
        );

    \I__5302\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23494\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__23513\,
            I => \N__23491\
        );

    \I__5300\ : Span4Mux_h
    port map (
            O => \N__23508\,
            I => \N__23488\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__23507\,
            I => \N__23485\
        );

    \I__5298\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23482\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__23503\,
            I => \N__23475\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__23500\,
            I => \N__23475\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__23497\,
            I => \N__23475\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__23494\,
            I => \N__23472\
        );

    \I__5293\ : Span4Mux_h
    port map (
            O => \N__23491\,
            I => \N__23467\
        );

    \I__5292\ : Span4Mux_v
    port map (
            O => \N__23488\,
            I => \N__23467\
        );

    \I__5291\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23464\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__23482\,
            I => \N__23461\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__23475\,
            I => \N__23458\
        );

    \I__5288\ : Span12Mux_s11_h
    port map (
            O => \N__23472\,
            I => \N__23455\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__23467\,
            I => \tok.S_7\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__23464\,
            I => \tok.S_7\
        );

    \I__5285\ : Odrv12
    port map (
            O => \N__23461\,
            I => \tok.S_7\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__23458\,
            I => \tok.S_7\
        );

    \I__5283\ : Odrv12
    port map (
            O => \N__23455\,
            I => \tok.S_7\
        );

    \I__5282\ : CascadeMux
    port map (
            O => \N__23444\,
            I => \N__23441\
        );

    \I__5281\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23438\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__23438\,
            I => \N__23435\
        );

    \I__5279\ : Odrv12
    port map (
            O => \N__23435\,
            I => \tok.n295\
        );

    \I__5278\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23429\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__23429\,
            I => \N__23426\
        );

    \I__5276\ : Span4Mux_h
    port map (
            O => \N__23426\,
            I => \N__23423\
        );

    \I__5275\ : Span4Mux_v
    port map (
            O => \N__23423\,
            I => \N__23420\
        );

    \I__5274\ : Odrv4
    port map (
            O => \N__23420\,
            I => \tok.n6_adj_657\
        );

    \I__5273\ : InMux
    port map (
            O => \N__23417\,
            I => \tok.n4775\
        );

    \I__5272\ : InMux
    port map (
            O => \N__23414\,
            I => \bfn_11_10_0_\
        );

    \I__5271\ : InMux
    port map (
            O => \N__23411\,
            I => \N__23407\
        );

    \I__5270\ : InMux
    port map (
            O => \N__23410\,
            I => \N__23403\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__23407\,
            I => \N__23399\
        );

    \I__5268\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23396\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__23403\,
            I => \N__23393\
        );

    \I__5266\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23390\
        );

    \I__5265\ : Span4Mux_v
    port map (
            O => \N__23399\,
            I => \N__23385\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__23396\,
            I => \N__23385\
        );

    \I__5263\ : Span4Mux_v
    port map (
            O => \N__23393\,
            I => \N__23378\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__23390\,
            I => \N__23378\
        );

    \I__5261\ : Span4Mux_h
    port map (
            O => \N__23385\,
            I => \N__23378\
        );

    \I__5260\ : Span4Mux_h
    port map (
            O => \N__23378\,
            I => \N__23374\
        );

    \I__5259\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23371\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__23374\,
            I => \tok.n11_adj_706\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__23371\,
            I => \tok.n11_adj_706\
        );

    \I__5256\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23362\
        );

    \I__5255\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23359\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__23362\,
            I => \N__23356\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__23359\,
            I => uart_rx_data_2
        );

    \I__5252\ : Odrv12
    port map (
            O => \N__23356\,
            I => uart_rx_data_2
        );

    \I__5251\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__5249\ : Span4Mux_v
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__5248\ : Odrv4
    port map (
            O => \N__23342\,
            I => \tok.n12_adj_832\
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__23339\,
            I => \tok.n6_adj_839_cascade_\
        );

    \I__5246\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23327\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__23335\,
            I => \N__23324\
        );

    \I__5244\ : InMux
    port map (
            O => \N__23334\,
            I => \N__23321\
        );

    \I__5243\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23318\
        );

    \I__5242\ : InMux
    port map (
            O => \N__23332\,
            I => \N__23315\
        );

    \I__5241\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23309\
        );

    \I__5240\ : InMux
    port map (
            O => \N__23330\,
            I => \N__23309\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__23327\,
            I => \N__23303\
        );

    \I__5238\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23300\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23297\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__23318\,
            I => \N__23292\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23292\
        );

    \I__5234\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23289\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__23309\,
            I => \N__23286\
        );

    \I__5232\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23279\
        );

    \I__5231\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23279\
        );

    \I__5230\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23279\
        );

    \I__5229\ : Span4Mux_h
    port map (
            O => \N__23303\,
            I => \N__23275\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__23300\,
            I => \N__23268\
        );

    \I__5227\ : Span4Mux_v
    port map (
            O => \N__23297\,
            I => \N__23268\
        );

    \I__5226\ : Span4Mux_h
    port map (
            O => \N__23292\,
            I => \N__23268\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__23289\,
            I => \N__23263\
        );

    \I__5224\ : Span4Mux_h
    port map (
            O => \N__23286\,
            I => \N__23263\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23260\
        );

    \I__5222\ : CascadeMux
    port map (
            O => \N__23278\,
            I => \N__23255\
        );

    \I__5221\ : Span4Mux_h
    port map (
            O => \N__23275\,
            I => \N__23252\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__23268\,
            I => \N__23249\
        );

    \I__5219\ : Span4Mux_h
    port map (
            O => \N__23263\,
            I => \N__23244\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__23260\,
            I => \N__23244\
        );

    \I__5217\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23239\
        );

    \I__5216\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23239\
        );

    \I__5215\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23236\
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__23252\,
            I => \tok.n11_adj_681\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__23249\,
            I => \tok.n11_adj_681\
        );

    \I__5212\ : Odrv4
    port map (
            O => \N__23244\,
            I => \tok.n11_adj_681\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__23239\,
            I => \tok.n11_adj_681\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__23236\,
            I => \tok.n11_adj_681\
        );

    \I__5209\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23222\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__23222\,
            I => \N__23219\
        );

    \I__5207\ : Span4Mux_h
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__5206\ : Odrv4
    port map (
            O => \N__23216\,
            I => \tok.n32\
        );

    \I__5205\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23209\
        );

    \I__5204\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23205\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__23209\,
            I => \N__23201\
        );

    \I__5202\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23198\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__23205\,
            I => \N__23195\
        );

    \I__5200\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23192\
        );

    \I__5199\ : Span4Mux_v
    port map (
            O => \N__23201\,
            I => \N__23189\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__23198\,
            I => \N__23186\
        );

    \I__5197\ : Span4Mux_v
    port map (
            O => \N__23195\,
            I => \N__23183\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__23192\,
            I => \N__23180\
        );

    \I__5195\ : Span4Mux_v
    port map (
            O => \N__23189\,
            I => \N__23177\
        );

    \I__5194\ : Span4Mux_v
    port map (
            O => \N__23186\,
            I => \N__23172\
        );

    \I__5193\ : Span4Mux_s3_v
    port map (
            O => \N__23183\,
            I => \N__23172\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__23180\,
            I => \N__23169\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__23177\,
            I => \tok.n15_adj_655\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__23172\,
            I => \tok.n15_adj_655\
        );

    \I__5189\ : Odrv4
    port map (
            O => \N__23169\,
            I => \tok.n15_adj_655\
        );

    \I__5188\ : InMux
    port map (
            O => \N__23162\,
            I => \N__23159\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__23159\,
            I => \N__23151\
        );

    \I__5186\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23147\
        );

    \I__5185\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23144\
        );

    \I__5184\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23141\
        );

    \I__5183\ : InMux
    port map (
            O => \N__23155\,
            I => \N__23138\
        );

    \I__5182\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23135\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__23151\,
            I => \N__23132\
        );

    \I__5180\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23129\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__23147\,
            I => \N__23126\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__23144\,
            I => \N__23123\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__23141\,
            I => \N__23120\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__23138\,
            I => \N__23117\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__23135\,
            I => \N__23113\
        );

    \I__5174\ : Span4Mux_v
    port map (
            O => \N__23132\,
            I => \N__23102\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__23129\,
            I => \N__23102\
        );

    \I__5172\ : Span4Mux_h
    port map (
            O => \N__23126\,
            I => \N__23102\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__23123\,
            I => \N__23102\
        );

    \I__5170\ : Span12Mux_s10_v
    port map (
            O => \N__23120\,
            I => \N__23099\
        );

    \I__5169\ : Span4Mux_s3_h
    port map (
            O => \N__23117\,
            I => \N__23096\
        );

    \I__5168\ : InMux
    port map (
            O => \N__23116\,
            I => \N__23093\
        );

    \I__5167\ : Span4Mux_s3_v
    port map (
            O => \N__23113\,
            I => \N__23090\
        );

    \I__5166\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23085\
        );

    \I__5165\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23085\
        );

    \I__5164\ : Span4Mux_v
    port map (
            O => \N__23102\,
            I => \N__23082\
        );

    \I__5163\ : Odrv12
    port map (
            O => \N__23099\,
            I => \tok.A_13\
        );

    \I__5162\ : Odrv4
    port map (
            O => \N__23096\,
            I => \tok.A_13\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__23093\,
            I => \tok.A_13\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__23090\,
            I => \tok.A_13\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__23085\,
            I => \tok.A_13\
        );

    \I__5158\ : Odrv4
    port map (
            O => \N__23082\,
            I => \tok.A_13\
        );

    \I__5157\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__23066\,
            I => \N__23063\
        );

    \I__5155\ : Span4Mux_v
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__5154\ : Span4Mux_h
    port map (
            O => \N__23060\,
            I => \N__23057\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__23057\,
            I => \tok.n211\
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \N__23051\
        );

    \I__5151\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23048\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__23048\,
            I => \N__23045\
        );

    \I__5149\ : Span4Mux_h
    port map (
            O => \N__23045\,
            I => \N__23042\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__23042\,
            I => \tok.n184\
        );

    \I__5147\ : InMux
    port map (
            O => \N__23039\,
            I => \N__23036\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__23036\,
            I => \N__23032\
        );

    \I__5145\ : InMux
    port map (
            O => \N__23035\,
            I => \N__23029\
        );

    \I__5144\ : Span4Mux_v
    port map (
            O => \N__23032\,
            I => \N__23024\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__23029\,
            I => \N__23024\
        );

    \I__5142\ : Span4Mux_h
    port map (
            O => \N__23024\,
            I => \N__23020\
        );

    \I__5141\ : InMux
    port map (
            O => \N__23023\,
            I => \N__23017\
        );

    \I__5140\ : Odrv4
    port map (
            O => \N__23020\,
            I => capture_5
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__23017\,
            I => capture_5
        );

    \I__5138\ : InMux
    port map (
            O => \N__23012\,
            I => \N__23009\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__23009\,
            I => \N__23005\
        );

    \I__5136\ : InMux
    port map (
            O => \N__23008\,
            I => \N__23002\
        );

    \I__5135\ : Span4Mux_s2_h
    port map (
            O => \N__23005\,
            I => \N__22997\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__23002\,
            I => \N__22997\
        );

    \I__5133\ : Span4Mux_h
    port map (
            O => \N__22997\,
            I => \N__22994\
        );

    \I__5132\ : Span4Mux_h
    port map (
            O => \N__22994\,
            I => \N__22990\
        );

    \I__5131\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22987\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__22990\,
            I => capture_8
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__22987\,
            I => capture_8
        );

    \I__5128\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22979\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__22979\,
            I => \N__22967\
        );

    \I__5126\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22964\
        );

    \I__5125\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22957\
        );

    \I__5124\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22957\
        );

    \I__5123\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22957\
        );

    \I__5122\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22952\
        );

    \I__5121\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22952\
        );

    \I__5120\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22945\
        );

    \I__5119\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22945\
        );

    \I__5118\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22945\
        );

    \I__5117\ : Span4Mux_v
    port map (
            O => \N__22967\,
            I => \N__22938\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__22964\,
            I => \N__22938\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__22957\,
            I => \N__22938\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__22952\,
            I => \N__22935\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__22945\,
            I => \N__22932\
        );

    \I__5112\ : Span4Mux_v
    port map (
            O => \N__22938\,
            I => \N__22927\
        );

    \I__5111\ : Span4Mux_h
    port map (
            O => \N__22935\,
            I => \N__22927\
        );

    \I__5110\ : Span12Mux_s9_v
    port map (
            O => \N__22932\,
            I => \N__22924\
        );

    \I__5109\ : Span4Mux_h
    port map (
            O => \N__22927\,
            I => \N__22921\
        );

    \I__5108\ : Odrv12
    port map (
            O => \N__22924\,
            I => n4858
        );

    \I__5107\ : Odrv4
    port map (
            O => \N__22921\,
            I => n4858
        );

    \I__5106\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__5104\ : Span4Mux_v
    port map (
            O => \N__22910\,
            I => \N__22907\
        );

    \I__5103\ : Span4Mux_h
    port map (
            O => \N__22907\,
            I => \N__22902\
        );

    \I__5102\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22897\
        );

    \I__5101\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22897\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__22902\,
            I => capture_7
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__22897\,
            I => capture_7
        );

    \I__5098\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22889\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__22889\,
            I => \tok.n17_adj_711\
        );

    \I__5096\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22883\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__22883\,
            I => \N__22876\
        );

    \I__5094\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22873\
        );

    \I__5093\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22868\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__22880\,
            I => \N__22865\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__22879\,
            I => \N__22862\
        );

    \I__5090\ : Span4Mux_h
    port map (
            O => \N__22876\,
            I => \N__22857\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__22873\,
            I => \N__22857\
        );

    \I__5088\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22854\
        );

    \I__5087\ : CascadeMux
    port map (
            O => \N__22871\,
            I => \N__22850\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__22868\,
            I => \N__22847\
        );

    \I__5085\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22844\
        );

    \I__5084\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22841\
        );

    \I__5083\ : Span4Mux_v
    port map (
            O => \N__22857\,
            I => \N__22835\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__22854\,
            I => \N__22835\
        );

    \I__5081\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22832\
        );

    \I__5080\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22829\
        );

    \I__5079\ : Span4Mux_v
    port map (
            O => \N__22847\,
            I => \N__22824\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__22844\,
            I => \N__22824\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__22841\,
            I => \N__22821\
        );

    \I__5076\ : InMux
    port map (
            O => \N__22840\,
            I => \N__22818\
        );

    \I__5075\ : Span4Mux_h
    port map (
            O => \N__22835\,
            I => \N__22815\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__22832\,
            I => \N__22812\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__22829\,
            I => \N__22809\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__22824\,
            I => \N__22806\
        );

    \I__5071\ : Span12Mux_v
    port map (
            O => \N__22821\,
            I => \N__22803\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__22818\,
            I => \N__22798\
        );

    \I__5069\ : Span4Mux_v
    port map (
            O => \N__22815\,
            I => \N__22798\
        );

    \I__5068\ : Span12Mux_s6_h
    port map (
            O => \N__22812\,
            I => \N__22793\
        );

    \I__5067\ : Span12Mux_s7_h
    port map (
            O => \N__22809\,
            I => \N__22793\
        );

    \I__5066\ : Span4Mux_v
    port map (
            O => \N__22806\,
            I => \N__22790\
        );

    \I__5065\ : Odrv12
    port map (
            O => \N__22803\,
            I => \tok.S_0\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__22798\,
            I => \tok.S_0\
        );

    \I__5063\ : Odrv12
    port map (
            O => \N__22793\,
            I => \tok.S_0\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__22790\,
            I => \tok.S_0\
        );

    \I__5061\ : InMux
    port map (
            O => \N__22781\,
            I => \N__22778\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__22778\,
            I => \N__22775\
        );

    \I__5059\ : Span4Mux_h
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__22772\,
            I => \tok.n11_adj_809\
        );

    \I__5057\ : InMux
    port map (
            O => \N__22769\,
            I => \bfn_11_9_0_\
        );

    \I__5056\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22754\
        );

    \I__5055\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22751\
        );

    \I__5054\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22747\
        );

    \I__5053\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22742\
        );

    \I__5052\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22742\
        );

    \I__5051\ : InMux
    port map (
            O => \N__22761\,
            I => \N__22739\
        );

    \I__5050\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22736\
        );

    \I__5049\ : InMux
    port map (
            O => \N__22759\,
            I => \N__22733\
        );

    \I__5048\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22728\
        );

    \I__5047\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22725\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__22754\,
            I => \N__22722\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__22751\,
            I => \N__22719\
        );

    \I__5044\ : InMux
    port map (
            O => \N__22750\,
            I => \N__22716\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__22747\,
            I => \N__22711\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__22742\,
            I => \N__22711\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__22739\,
            I => \N__22702\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__22736\,
            I => \N__22702\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__22733\,
            I => \N__22702\
        );

    \I__5038\ : InMux
    port map (
            O => \N__22732\,
            I => \N__22699\
        );

    \I__5037\ : CascadeMux
    port map (
            O => \N__22731\,
            I => \N__22696\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__22728\,
            I => \N__22693\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__22725\,
            I => \N__22690\
        );

    \I__5034\ : Span4Mux_h
    port map (
            O => \N__22722\,
            I => \N__22685\
        );

    \I__5033\ : Span4Mux_h
    port map (
            O => \N__22719\,
            I => \N__22685\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22682\
        );

    \I__5031\ : Span12Mux_s9_v
    port map (
            O => \N__22711\,
            I => \N__22679\
        );

    \I__5030\ : InMux
    port map (
            O => \N__22710\,
            I => \N__22674\
        );

    \I__5029\ : InMux
    port map (
            O => \N__22709\,
            I => \N__22674\
        );

    \I__5028\ : Span4Mux_v
    port map (
            O => \N__22702\,
            I => \N__22669\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__22699\,
            I => \N__22669\
        );

    \I__5026\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22666\
        );

    \I__5025\ : Span4Mux_v
    port map (
            O => \N__22693\,
            I => \N__22661\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__22690\,
            I => \N__22661\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__22685\,
            I => \tok.A_low_2\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__22682\,
            I => \tok.A_low_2\
        );

    \I__5021\ : Odrv12
    port map (
            O => \N__22679\,
            I => \tok.A_low_2\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__22674\,
            I => \tok.A_low_2\
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__22669\,
            I => \tok.A_low_2\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__22666\,
            I => \tok.A_low_2\
        );

    \I__5017\ : Odrv4
    port map (
            O => \N__22661\,
            I => \tok.A_low_2\
        );

    \I__5016\ : InMux
    port map (
            O => \N__22646\,
            I => \N__22643\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__22643\,
            I => \N__22640\
        );

    \I__5014\ : Span4Mux_s3_h
    port map (
            O => \N__22640\,
            I => \N__22637\
        );

    \I__5013\ : Odrv4
    port map (
            O => \N__22637\,
            I => \tok.n22_adj_698\
        );

    \I__5012\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22631\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__22631\,
            I => \N__22628\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__22628\,
            I => \N__22625\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__22625\,
            I => \N__22622\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__22622\,
            I => \tok.n24_adj_703\
        );

    \I__5007\ : CascadeMux
    port map (
            O => \N__22619\,
            I => \tok.n4_adj_699_cascade_\
        );

    \I__5006\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22613\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__22613\,
            I => \N__22610\
        );

    \I__5004\ : Span4Mux_h
    port map (
            O => \N__22610\,
            I => \N__22607\
        );

    \I__5003\ : Odrv4
    port map (
            O => \N__22607\,
            I => \tok.n9_adj_705\
        );

    \I__5002\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22601\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22597\
        );

    \I__5000\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22594\
        );

    \I__4999\ : Span4Mux_s3_h
    port map (
            O => \N__22597\,
            I => \N__22591\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__22594\,
            I => uart_rx_data_1
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__22591\,
            I => uart_rx_data_1
        );

    \I__4996\ : InMux
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__4994\ : Span12Mux_s4_h
    port map (
            O => \N__22580\,
            I => \N__22577\
        );

    \I__4993\ : Odrv12
    port map (
            O => \N__22577\,
            I => \tok.n14_adj_662\
        );

    \I__4992\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22571\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__22571\,
            I => \tok.n6_adj_834\
        );

    \I__4990\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__4988\ : Span4Mux_v
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__4987\ : Span4Mux_h
    port map (
            O => \N__22559\,
            I => \N__22556\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__22556\,
            I => \tok.n23_adj_718\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__22553\,
            I => \tok.n5_adj_835_cascade_\
        );

    \I__4984\ : InMux
    port map (
            O => \N__22550\,
            I => \N__22536\
        );

    \I__4983\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22533\
        );

    \I__4982\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22530\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__22547\,
            I => \N__22524\
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__22546\,
            I => \N__22520\
        );

    \I__4979\ : CascadeMux
    port map (
            O => \N__22545\,
            I => \N__22517\
        );

    \I__4978\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22512\
        );

    \I__4977\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22512\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__22542\,
            I => \N__22498\
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__22541\,
            I => \N__22493\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__22540\,
            I => \N__22489\
        );

    \I__4973\ : InMux
    port map (
            O => \N__22539\,
            I => \N__22486\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__22536\,
            I => \N__22482\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__22533\,
            I => \N__22474\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__22530\,
            I => \N__22474\
        );

    \I__4969\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22469\
        );

    \I__4968\ : InMux
    port map (
            O => \N__22528\,
            I => \N__22469\
        );

    \I__4967\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22466\
        );

    \I__4966\ : InMux
    port map (
            O => \N__22524\,
            I => \N__22457\
        );

    \I__4965\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22457\
        );

    \I__4964\ : InMux
    port map (
            O => \N__22520\,
            I => \N__22457\
        );

    \I__4963\ : InMux
    port map (
            O => \N__22517\,
            I => \N__22457\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__22512\,
            I => \N__22454\
        );

    \I__4961\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22451\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__22510\,
            I => \N__22447\
        );

    \I__4959\ : InMux
    port map (
            O => \N__22509\,
            I => \N__22432\
        );

    \I__4958\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22432\
        );

    \I__4957\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22432\
        );

    \I__4956\ : InMux
    port map (
            O => \N__22506\,
            I => \N__22432\
        );

    \I__4955\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22432\
        );

    \I__4954\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22432\
        );

    \I__4953\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22432\
        );

    \I__4952\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22415\
        );

    \I__4951\ : InMux
    port map (
            O => \N__22501\,
            I => \N__22415\
        );

    \I__4950\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22415\
        );

    \I__4949\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22415\
        );

    \I__4948\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22415\
        );

    \I__4947\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22415\
        );

    \I__4946\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22415\
        );

    \I__4945\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22415\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22412\
        );

    \I__4943\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22408\
        );

    \I__4942\ : Span4Mux_v
    port map (
            O => \N__22482\,
            I => \N__22405\
        );

    \I__4941\ : InMux
    port map (
            O => \N__22481\,
            I => \N__22398\
        );

    \I__4940\ : InMux
    port map (
            O => \N__22480\,
            I => \N__22398\
        );

    \I__4939\ : InMux
    port map (
            O => \N__22479\,
            I => \N__22398\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__22474\,
            I => \N__22389\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__22469\,
            I => \N__22389\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__22466\,
            I => \N__22389\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__22457\,
            I => \N__22389\
        );

    \I__4934\ : Span4Mux_h
    port map (
            O => \N__22454\,
            I => \N__22384\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__22451\,
            I => \N__22384\
        );

    \I__4932\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22379\
        );

    \I__4931\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22379\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__22432\,
            I => \N__22374\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__22415\,
            I => \N__22374\
        );

    \I__4928\ : Span4Mux_v
    port map (
            O => \N__22412\,
            I => \N__22371\
        );

    \I__4927\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22368\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__22408\,
            I => \N__22361\
        );

    \I__4925\ : Span4Mux_v
    port map (
            O => \N__22405\,
            I => \N__22361\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__22398\,
            I => \N__22361\
        );

    \I__4923\ : Span4Mux_h
    port map (
            O => \N__22389\,
            I => \N__22358\
        );

    \I__4922\ : Span4Mux_h
    port map (
            O => \N__22384\,
            I => \N__22353\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__22379\,
            I => \N__22353\
        );

    \I__4920\ : Odrv4
    port map (
            O => \N__22374\,
            I => \tok.n14_adj_644\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__22371\,
            I => \tok.n14_adj_644\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__22368\,
            I => \tok.n14_adj_644\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__22361\,
            I => \tok.n14_adj_644\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__22358\,
            I => \tok.n14_adj_644\
        );

    \I__4915\ : Odrv4
    port map (
            O => \N__22353\,
            I => \tok.n14_adj_644\
        );

    \I__4914\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__4912\ : Span4Mux_h
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__4911\ : Odrv4
    port map (
            O => \N__22331\,
            I => \tok.n10_adj_836\
        );

    \I__4910\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22323\
        );

    \I__4909\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22317\
        );

    \I__4908\ : InMux
    port map (
            O => \N__22326\,
            I => \N__22314\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N__22307\
        );

    \I__4906\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22304\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__22321\,
            I => \N__22300\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__22320\,
            I => \N__22296\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__22317\,
            I => \N__22293\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__22314\,
            I => \N__22290\
        );

    \I__4901\ : CascadeMux
    port map (
            O => \N__22313\,
            I => \N__22287\
        );

    \I__4900\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22282\
        );

    \I__4899\ : InMux
    port map (
            O => \N__22311\,
            I => \N__22282\
        );

    \I__4898\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22279\
        );

    \I__4897\ : Span4Mux_v
    port map (
            O => \N__22307\,
            I => \N__22276\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__22304\,
            I => \N__22273\
        );

    \I__4895\ : InMux
    port map (
            O => \N__22303\,
            I => \N__22270\
        );

    \I__4894\ : InMux
    port map (
            O => \N__22300\,
            I => \N__22265\
        );

    \I__4893\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22262\
        );

    \I__4892\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22259\
        );

    \I__4891\ : Span4Mux_v
    port map (
            O => \N__22293\,
            I => \N__22253\
        );

    \I__4890\ : Span4Mux_v
    port map (
            O => \N__22290\,
            I => \N__22253\
        );

    \I__4889\ : InMux
    port map (
            O => \N__22287\,
            I => \N__22250\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__22282\,
            I => \N__22247\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__22279\,
            I => \N__22244\
        );

    \I__4886\ : Span4Mux_h
    port map (
            O => \N__22276\,
            I => \N__22237\
        );

    \I__4885\ : Span4Mux_h
    port map (
            O => \N__22273\,
            I => \N__22237\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22237\
        );

    \I__4883\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22234\
        );

    \I__4882\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22231\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__22265\,
            I => \N__22228\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__22262\,
            I => \N__22225\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__22259\,
            I => \N__22222\
        );

    \I__4878\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22219\
        );

    \I__4877\ : Span4Mux_h
    port map (
            O => \N__22253\,
            I => \N__22210\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22210\
        );

    \I__4875\ : Span4Mux_v
    port map (
            O => \N__22247\,
            I => \N__22210\
        );

    \I__4874\ : Span4Mux_v
    port map (
            O => \N__22244\,
            I => \N__22210\
        );

    \I__4873\ : Sp12to4
    port map (
            O => \N__22237\,
            I => \N__22203\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__22234\,
            I => \N__22203\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__22231\,
            I => \N__22203\
        );

    \I__4870\ : Span4Mux_v
    port map (
            O => \N__22228\,
            I => \N__22196\
        );

    \I__4869\ : Span4Mux_v
    port map (
            O => \N__22225\,
            I => \N__22196\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__22222\,
            I => \N__22196\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__22219\,
            I => \A_low_7\
        );

    \I__4866\ : Odrv4
    port map (
            O => \N__22210\,
            I => \A_low_7\
        );

    \I__4865\ : Odrv12
    port map (
            O => \N__22203\,
            I => \A_low_7\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__22196\,
            I => \A_low_7\
        );

    \I__4863\ : CascadeMux
    port map (
            O => \N__22187\,
            I => \N__22183\
        );

    \I__4862\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22179\
        );

    \I__4861\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22174\
        );

    \I__4860\ : InMux
    port map (
            O => \N__22182\,
            I => \N__22174\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__22179\,
            I => \N__22171\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__22174\,
            I => \N__22167\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__22171\,
            I => \N__22164\
        );

    \I__4856\ : InMux
    port map (
            O => \N__22170\,
            I => \N__22161\
        );

    \I__4855\ : Span4Mux_v
    port map (
            O => \N__22167\,
            I => \N__22158\
        );

    \I__4854\ : Odrv4
    port map (
            O => \N__22164\,
            I => \tok.n6_adj_650\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__22161\,
            I => \tok.n6_adj_650\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__22158\,
            I => \tok.n6_adj_650\
        );

    \I__4851\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22147\
        );

    \I__4850\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22136\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__22147\,
            I => \N__22131\
        );

    \I__4848\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22126\
        );

    \I__4847\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22126\
        );

    \I__4846\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22123\
        );

    \I__4845\ : InMux
    port map (
            O => \N__22143\,
            I => \N__22116\
        );

    \I__4844\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22116\
        );

    \I__4843\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22116\
        );

    \I__4842\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22111\
        );

    \I__4841\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22111\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__22136\,
            I => \N__22104\
        );

    \I__4839\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22099\
        );

    \I__4838\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22099\
        );

    \I__4837\ : Span4Mux_v
    port map (
            O => \N__22131\,
            I => \N__22094\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__22126\,
            I => \N__22094\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__22123\,
            I => \N__22089\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__22116\,
            I => \N__22089\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__22111\,
            I => \N__22086\
        );

    \I__4832\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22083\
        );

    \I__4831\ : InMux
    port map (
            O => \N__22109\,
            I => \N__22078\
        );

    \I__4830\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22078\
        );

    \I__4829\ : CascadeMux
    port map (
            O => \N__22107\,
            I => \N__22074\
        );

    \I__4828\ : Span4Mux_s3_v
    port map (
            O => \N__22104\,
            I => \N__22069\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__22099\,
            I => \N__22069\
        );

    \I__4826\ : Span4Mux_h
    port map (
            O => \N__22094\,
            I => \N__22064\
        );

    \I__4825\ : Span4Mux_v
    port map (
            O => \N__22089\,
            I => \N__22064\
        );

    \I__4824\ : Span4Mux_h
    port map (
            O => \N__22086\,
            I => \N__22060\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__22083\,
            I => \N__22057\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__22078\,
            I => \N__22054\
        );

    \I__4821\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22049\
        );

    \I__4820\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22049\
        );

    \I__4819\ : Span4Mux_v
    port map (
            O => \N__22069\,
            I => \N__22044\
        );

    \I__4818\ : Span4Mux_h
    port map (
            O => \N__22064\,
            I => \N__22044\
        );

    \I__4817\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22041\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__22060\,
            I => \N__22038\
        );

    \I__4815\ : Span4Mux_s3_v
    port map (
            O => \N__22057\,
            I => \N__22033\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__22054\,
            I => \N__22033\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__22049\,
            I => \N__22030\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__22044\,
            I => \tok.T_7\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__22041\,
            I => \tok.T_7\
        );

    \I__4810\ : Odrv4
    port map (
            O => \N__22038\,
            I => \tok.T_7\
        );

    \I__4809\ : Odrv4
    port map (
            O => \N__22033\,
            I => \tok.T_7\
        );

    \I__4808\ : Odrv12
    port map (
            O => \N__22030\,
            I => \tok.T_7\
        );

    \I__4807\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22013\
        );

    \I__4806\ : InMux
    port map (
            O => \N__22018\,
            I => \N__22013\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__22013\,
            I => \tok.A_stk.tail_8\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__22010\,
            I => \N__22006\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__22009\,
            I => \N__22003\
        );

    \I__4802\ : InMux
    port map (
            O => \N__22006\,
            I => \N__21998\
        );

    \I__4801\ : InMux
    port map (
            O => \N__22003\,
            I => \N__21998\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__21998\,
            I => \tok.A_stk.tail_24\
        );

    \I__4799\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__21992\,
            I => \N__21989\
        );

    \I__4797\ : Span4Mux_v
    port map (
            O => \N__21989\,
            I => \N__21985\
        );

    \I__4796\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21982\
        );

    \I__4795\ : Odrv4
    port map (
            O => \N__21985\,
            I => \tok.A_stk.tail_56\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__21982\,
            I => \tok.A_stk.tail_56\
        );

    \I__4793\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21970\
        );

    \I__4791\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21967\
        );

    \I__4790\ : Span4Mux_h
    port map (
            O => \N__21970\,
            I => \N__21964\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__21967\,
            I => \tok.A_stk.tail_40\
        );

    \I__4788\ : Odrv4
    port map (
            O => \N__21964\,
            I => \tok.A_stk.tail_40\
        );

    \I__4787\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__21953\,
            I => \tok.n22\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__4783\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__4781\ : Span4Mux_s3_h
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__4780\ : Span4Mux_v
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__4779\ : Odrv4
    port map (
            O => \N__21935\,
            I => \tok.n24\
        );

    \I__4778\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__4776\ : Span4Mux_s3_h
    port map (
            O => \N__21926\,
            I => \N__21923\
        );

    \I__4775\ : Span4Mux_h
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__21920\,
            I => \tok.n21\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__21917\,
            I => \tok.n30_cascade_\
        );

    \I__4772\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21911\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__21911\,
            I => \N__21907\
        );

    \I__4770\ : InMux
    port map (
            O => \N__21910\,
            I => \N__21904\
        );

    \I__4769\ : Span12Mux_s8_v
    port map (
            O => \N__21907\,
            I => \N__21899\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__21904\,
            I => \N__21899\
        );

    \I__4767\ : Odrv12
    port map (
            O => \N__21899\,
            I => \tok.n15_adj_671\
        );

    \I__4766\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21890\
        );

    \I__4765\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21887\
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__21894\,
            I => \N__21883\
        );

    \I__4763\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21880\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__21890\,
            I => \N__21877\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__21887\,
            I => \N__21872\
        );

    \I__4760\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21869\
        );

    \I__4759\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21861\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__21880\,
            I => \N__21856\
        );

    \I__4757\ : Span4Mux_h
    port map (
            O => \N__21877\,
            I => \N__21856\
        );

    \I__4756\ : InMux
    port map (
            O => \N__21876\,
            I => \N__21851\
        );

    \I__4755\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21851\
        );

    \I__4754\ : Span4Mux_v
    port map (
            O => \N__21872\,
            I => \N__21846\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__21869\,
            I => \N__21846\
        );

    \I__4752\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21841\
        );

    \I__4751\ : InMux
    port map (
            O => \N__21867\,
            I => \N__21841\
        );

    \I__4750\ : InMux
    port map (
            O => \N__21866\,
            I => \N__21836\
        );

    \I__4749\ : InMux
    port map (
            O => \N__21865\,
            I => \N__21836\
        );

    \I__4748\ : InMux
    port map (
            O => \N__21864\,
            I => \N__21831\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__21861\,
            I => \N__21827\
        );

    \I__4746\ : Span4Mux_h
    port map (
            O => \N__21856\,
            I => \N__21818\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__21851\,
            I => \N__21818\
        );

    \I__4744\ : Span4Mux_h
    port map (
            O => \N__21846\,
            I => \N__21818\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__21841\,
            I => \N__21818\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__21836\,
            I => \N__21815\
        );

    \I__4741\ : InMux
    port map (
            O => \N__21835\,
            I => \N__21812\
        );

    \I__4740\ : InMux
    port map (
            O => \N__21834\,
            I => \N__21809\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__21831\,
            I => \N__21806\
        );

    \I__4738\ : InMux
    port map (
            O => \N__21830\,
            I => \N__21803\
        );

    \I__4737\ : Span4Mux_h
    port map (
            O => \N__21827\,
            I => \N__21798\
        );

    \I__4736\ : Span4Mux_v
    port map (
            O => \N__21818\,
            I => \N__21798\
        );

    \I__4735\ : Span4Mux_v
    port map (
            O => \N__21815\,
            I => \N__21795\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__21812\,
            I => \tok.A_low_6\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__21809\,
            I => \tok.A_low_6\
        );

    \I__4732\ : Odrv12
    port map (
            O => \N__21806\,
            I => \tok.A_low_6\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__21803\,
            I => \tok.A_low_6\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__21798\,
            I => \tok.A_low_6\
        );

    \I__4729\ : Odrv4
    port map (
            O => \N__21795\,
            I => \tok.A_low_6\
        );

    \I__4728\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__4726\ : Span4Mux_s3_h
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__4725\ : Span4Mux_v
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__4724\ : Odrv4
    port map (
            O => \N__21770\,
            I => \tok.n18\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__21767\,
            I => \tok.n17_adj_661_cascade_\
        );

    \I__4722\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__21761\,
            I => \tok.n19\
        );

    \I__4720\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__21755\,
            I => \tok.n29\
        );

    \I__4718\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__21749\,
            I => \N__21746\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__21746\,
            I => \N__21742\
        );

    \I__4715\ : InMux
    port map (
            O => \N__21745\,
            I => \N__21739\
        );

    \I__4714\ : Odrv4
    port map (
            O => \N__21742\,
            I => \tok.A_stk.tail_7\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__21739\,
            I => \tok.A_stk.tail_7\
        );

    \I__4712\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21728\
        );

    \I__4711\ : InMux
    port map (
            O => \N__21733\,
            I => \N__21728\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__21728\,
            I => \tok.A_stk.tail_2\
        );

    \I__4709\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21719\
        );

    \I__4708\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21719\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__21719\,
            I => \tok.A_stk.tail_18\
        );

    \I__4706\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21710\
        );

    \I__4705\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21710\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__21710\,
            I => \tok.A_stk.tail_34\
        );

    \I__4703\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21704\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__21704\,
            I => \N__21700\
        );

    \I__4701\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21697\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__21700\,
            I => \tok.A_stk.tail_66\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__21697\,
            I => \tok.A_stk.tail_66\
        );

    \I__4698\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21688\
        );

    \I__4697\ : InMux
    port map (
            O => \N__21691\,
            I => \N__21685\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__21688\,
            I => \N__21682\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__21685\,
            I => \tok.A_stk.tail_50\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__21682\,
            I => \tok.A_stk.tail_50\
        );

    \I__4693\ : InMux
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__21674\,
            I => \N__21670\
        );

    \I__4691\ : InMux
    port map (
            O => \N__21673\,
            I => \N__21667\
        );

    \I__4690\ : Odrv4
    port map (
            O => \N__21670\,
            I => \tok.A_stk.tail_44\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__21667\,
            I => \tok.A_stk.tail_44\
        );

    \I__4688\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21658\
        );

    \I__4687\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21655\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__21658\,
            I => \N__21652\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__21655\,
            I => \tok.A_stk.tail_28\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__21652\,
            I => \tok.A_stk.tail_28\
        );

    \I__4683\ : CascadeMux
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__4682\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21638\
        );

    \I__4681\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21638\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__21638\,
            I => \tok.A_stk.tail_12\
        );

    \I__4679\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21626\
        );

    \I__4678\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21626\
        );

    \I__4677\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21623\
        );

    \I__4676\ : InMux
    port map (
            O => \N__21632\,
            I => \N__21620\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__21631\,
            I => \N__21616\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__21626\,
            I => \N__21613\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__21623\,
            I => \N__21608\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__21620\,
            I => \N__21605\
        );

    \I__4671\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21600\
        );

    \I__4670\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21600\
        );

    \I__4669\ : Span4Mux_s3_h
    port map (
            O => \N__21613\,
            I => \N__21596\
        );

    \I__4668\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21592\
        );

    \I__4667\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21589\
        );

    \I__4666\ : Span4Mux_h
    port map (
            O => \N__21608\,
            I => \N__21582\
        );

    \I__4665\ : Span4Mux_v
    port map (
            O => \N__21605\,
            I => \N__21582\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__21600\,
            I => \N__21582\
        );

    \I__4663\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21579\
        );

    \I__4662\ : Span4Mux_v
    port map (
            O => \N__21596\,
            I => \N__21576\
        );

    \I__4661\ : InMux
    port map (
            O => \N__21595\,
            I => \N__21573\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__21592\,
            I => \N__21566\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__21589\,
            I => \N__21566\
        );

    \I__4658\ : Span4Mux_h
    port map (
            O => \N__21582\,
            I => \N__21566\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__21579\,
            I => \tok.A_12\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__21576\,
            I => \tok.A_12\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__21573\,
            I => \tok.A_12\
        );

    \I__4654\ : Odrv4
    port map (
            O => \N__21566\,
            I => \tok.A_12\
        );

    \I__4653\ : InMux
    port map (
            O => \N__21557\,
            I => \N__21554\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__21554\,
            I => \N__21550\
        );

    \I__4651\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21547\
        );

    \I__4650\ : Odrv4
    port map (
            O => \N__21550\,
            I => tail_107
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__21547\,
            I => tail_107
        );

    \I__4648\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21538\
        );

    \I__4647\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21535\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__21538\,
            I => \tok.A_stk.tail_91\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__21535\,
            I => \tok.A_stk.tail_91\
        );

    \I__4644\ : CascadeMux
    port map (
            O => \N__21530\,
            I => \N__21526\
        );

    \I__4643\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21523\
        );

    \I__4642\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21520\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__21523\,
            I => \N__21517\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__21520\,
            I => \N__21514\
        );

    \I__4639\ : Odrv4
    port map (
            O => \N__21517\,
            I => tail_124
        );

    \I__4638\ : Odrv4
    port map (
            O => \N__21514\,
            I => tail_124
        );

    \I__4637\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21506\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__21506\,
            I => \N__21502\
        );

    \I__4635\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21499\
        );

    \I__4634\ : Odrv4
    port map (
            O => \N__21502\,
            I => tail_108
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__21499\,
            I => tail_108
        );

    \I__4632\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21488\
        );

    \I__4631\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21488\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__21488\,
            I => \tok.A_stk.tail_92\
        );

    \I__4629\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21479\
        );

    \I__4628\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21479\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__21479\,
            I => \tok.A_stk.tail_76\
        );

    \I__4626\ : InMux
    port map (
            O => \N__21476\,
            I => \N__21470\
        );

    \I__4625\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21470\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__21470\,
            I => \tok.A_stk.tail_60\
        );

    \I__4623\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21464\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__21464\,
            I => \N__21461\
        );

    \I__4621\ : Span4Mux_s2_v
    port map (
            O => \N__21461\,
            I => \N__21457\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__21460\,
            I => \N__21454\
        );

    \I__4619\ : Span4Mux_s1_h
    port map (
            O => \N__21457\,
            I => \N__21451\
        );

    \I__4618\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21448\
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__21451\,
            I => tail_125
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__21448\,
            I => tail_125
        );

    \I__4615\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21440\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__4613\ : Span4Mux_h
    port map (
            O => \N__21437\,
            I => \N__21433\
        );

    \I__4612\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21430\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__21433\,
            I => tail_109
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__21430\,
            I => tail_109
        );

    \I__4609\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21421\
        );

    \I__4608\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21418\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__21421\,
            I => \tok.A_stk.tail_93\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__21418\,
            I => \tok.A_stk.tail_93\
        );

    \I__4605\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21407\
        );

    \I__4604\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21407\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__21407\,
            I => \tok.A_stk.tail_77\
        );

    \I__4602\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21398\
        );

    \I__4601\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21398\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__21398\,
            I => \tok.A_stk.tail_61\
        );

    \I__4599\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21389\
        );

    \I__4598\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21389\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__21389\,
            I => \tok.A_stk.tail_45\
        );

    \I__4596\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21380\
        );

    \I__4595\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21380\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__21380\,
            I => \tok.A_stk.tail_29\
        );

    \I__4593\ : CascadeMux
    port map (
            O => \N__21377\,
            I => \N__21374\
        );

    \I__4592\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21368\
        );

    \I__4591\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21368\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__21368\,
            I => \tok.A_stk.tail_13\
        );

    \I__4589\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21362\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__21362\,
            I => \N__21358\
        );

    \I__4587\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21355\
        );

    \I__4586\ : Odrv12
    port map (
            O => \N__21358\,
            I => tail_123
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__21355\,
            I => tail_123
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__21350\,
            I => \tok.n13_adj_746_cascade_\
        );

    \I__4583\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__21344\,
            I => \tok.n12_adj_745\
        );

    \I__4581\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21338\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__21338\,
            I => \N__21335\
        );

    \I__4579\ : Span4Mux_v
    port map (
            O => \N__21335\,
            I => \N__21332\
        );

    \I__4578\ : Odrv4
    port map (
            O => \N__21332\,
            I => \tok.n5525\
        );

    \I__4577\ : InMux
    port map (
            O => \N__21329\,
            I => \N__21326\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__21326\,
            I => \tok.n16_adj_749\
        );

    \I__4575\ : CascadeMux
    port map (
            O => \N__21323\,
            I => \tok.n20_adj_753_cascade_\
        );

    \I__4574\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21317\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__21317\,
            I => \tok.n5522\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__21314\,
            I => \N__21308\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__21313\,
            I => \N__21305\
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__21312\,
            I => \N__21301\
        );

    \I__4569\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21298\
        );

    \I__4568\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21295\
        );

    \I__4567\ : InMux
    port map (
            O => \N__21305\,
            I => \N__21292\
        );

    \I__4566\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21289\
        );

    \I__4565\ : InMux
    port map (
            O => \N__21301\,
            I => \N__21286\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__21298\,
            I => \N__21275\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__21295\,
            I => \N__21275\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__21292\,
            I => \N__21275\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__21289\,
            I => \N__21275\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__21286\,
            I => \N__21275\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__21275\,
            I => \N__21272\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__21272\,
            I => \tok.n8\
        );

    \I__4557\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21266\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__21266\,
            I => \tok.n14_adj_744\
        );

    \I__4555\ : InMux
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__21260\,
            I => \tok.n9_adj_748\
        );

    \I__4553\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__21254\,
            I => \tok.n2_adj_743\
        );

    \I__4551\ : CascadeMux
    port map (
            O => \N__21251\,
            I => \tok.n204_cascade_\
        );

    \I__4550\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__21245\,
            I => \N__21242\
        );

    \I__4548\ : Odrv12
    port map (
            O => \N__21242\,
            I => \tok.n16_adj_741\
        );

    \I__4547\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21236\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__21236\,
            I => \N__21233\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__21233\,
            I => \tok.n2\
        );

    \I__4544\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21227\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__21227\,
            I => \tok.n14_adj_722\
        );

    \I__4542\ : InMux
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__4540\ : Odrv12
    port map (
            O => \N__21218\,
            I => \tok.n20_adj_740\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__21215\,
            I => \tok.n5527_cascade_\
        );

    \I__4538\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21209\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__21209\,
            I => \tok.n5513\
        );

    \I__4536\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21203\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__4534\ : Odrv4
    port map (
            O => \N__21200\,
            I => \tok.n5539\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__4532\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__21191\,
            I => \tok.n5348\
        );

    \I__4530\ : InMux
    port map (
            O => \N__21188\,
            I => \N__21185\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__21185\,
            I => \N__21180\
        );

    \I__4528\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21177\
        );

    \I__4527\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21174\
        );

    \I__4526\ : Span4Mux_v
    port map (
            O => \N__21180\,
            I => \N__21171\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__21177\,
            I => \N__21168\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__21174\,
            I => \N__21165\
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__21171\,
            I => capture_2
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__21168\,
            I => capture_2
        );

    \I__4521\ : Odrv4
    port map (
            O => \N__21165\,
            I => capture_2
        );

    \I__4520\ : InMux
    port map (
            O => \N__21158\,
            I => \N__21155\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__21155\,
            I => \tok.n9\
        );

    \I__4518\ : CascadeMux
    port map (
            O => \N__21152\,
            I => \tok.n5342_cascade_\
        );

    \I__4517\ : InMux
    port map (
            O => \N__21149\,
            I => \N__21146\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__21146\,
            I => \tok.n10_adj_686\
        );

    \I__4515\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21137\
        );

    \I__4514\ : InMux
    port map (
            O => \N__21142\,
            I => \N__21132\
        );

    \I__4513\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21128\
        );

    \I__4512\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21125\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__21137\,
            I => \N__21122\
        );

    \I__4510\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21119\
        );

    \I__4509\ : InMux
    port map (
            O => \N__21135\,
            I => \N__21116\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__21132\,
            I => \N__21112\
        );

    \I__4507\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21104\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__21128\,
            I => \N__21100\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__21125\,
            I => \N__21097\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__21122\,
            I => \N__21094\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__21119\,
            I => \N__21091\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__21116\,
            I => \N__21088\
        );

    \I__4501\ : InMux
    port map (
            O => \N__21115\,
            I => \N__21085\
        );

    \I__4500\ : Span4Mux_h
    port map (
            O => \N__21112\,
            I => \N__21081\
        );

    \I__4499\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21076\
        );

    \I__4498\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21076\
        );

    \I__4497\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21073\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__21108\,
            I => \N__21070\
        );

    \I__4495\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21067\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21064\
        );

    \I__4493\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21061\
        );

    \I__4492\ : Span4Mux_v
    port map (
            O => \N__21100\,
            I => \N__21056\
        );

    \I__4491\ : Span4Mux_v
    port map (
            O => \N__21097\,
            I => \N__21056\
        );

    \I__4490\ : Span4Mux_v
    port map (
            O => \N__21094\,
            I => \N__21047\
        );

    \I__4489\ : Span4Mux_h
    port map (
            O => \N__21091\,
            I => \N__21047\
        );

    \I__4488\ : Span4Mux_h
    port map (
            O => \N__21088\,
            I => \N__21047\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__21085\,
            I => \N__21047\
        );

    \I__4486\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21044\
        );

    \I__4485\ : Span4Mux_v
    port map (
            O => \N__21081\,
            I => \N__21037\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__21076\,
            I => \N__21037\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__21073\,
            I => \N__21037\
        );

    \I__4482\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21034\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__21067\,
            I => \N__21031\
        );

    \I__4480\ : Span4Mux_h
    port map (
            O => \N__21064\,
            I => \N__21026\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__21061\,
            I => \N__21026\
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__21056\,
            I => \tok.A_low_1\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__21047\,
            I => \tok.A_low_1\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__21044\,
            I => \tok.A_low_1\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__21037\,
            I => \tok.A_low_1\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__21034\,
            I => \tok.A_low_1\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__21031\,
            I => \tok.A_low_1\
        );

    \I__4472\ : Odrv4
    port map (
            O => \N__21026\,
            I => \tok.A_low_1\
        );

    \I__4471\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21008\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__21008\,
            I => \tok.n5336\
        );

    \I__4469\ : InMux
    port map (
            O => \N__21005\,
            I => \N__21002\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__21002\,
            I => \N__20999\
        );

    \I__4467\ : Span4Mux_v
    port map (
            O => \N__20999\,
            I => \N__20996\
        );

    \I__4466\ : Span4Mux_h
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__4465\ : Sp12to4
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__4464\ : Odrv12
    port map (
            O => \N__20990\,
            I => \tok.table_rd_11\
        );

    \I__4463\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__20984\,
            I => \N__20981\
        );

    \I__4461\ : Span4Mux_v
    port map (
            O => \N__20981\,
            I => \N__20978\
        );

    \I__4460\ : Odrv4
    port map (
            O => \N__20978\,
            I => \tok.n5_adj_726\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__20975\,
            I => \tok.n13_adj_724_cascade_\
        );

    \I__4458\ : InMux
    port map (
            O => \N__20972\,
            I => \N__20969\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__20969\,
            I => \tok.n12_adj_723\
        );

    \I__4456\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20963\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__4454\ : Odrv12
    port map (
            O => \N__20960\,
            I => \tok.n5534\
        );

    \I__4453\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__20954\,
            I => \tok.n16\
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__20951\,
            I => \tok.n20_adj_729_cascade_\
        );

    \I__4450\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20945\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__20945\,
            I => \tok.n9_adj_725\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__20942\,
            I => \N__20939\
        );

    \I__4447\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__20936\,
            I => \N__20933\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__20933\,
            I => \tok.n5531\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__20930\,
            I => \tok.n1_cascade_\
        );

    \I__4443\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20924\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__20924\,
            I => \N__20921\
        );

    \I__4441\ : Span4Mux_h
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__20918\,
            I => \tok.n17_adj_656\
        );

    \I__4439\ : InMux
    port map (
            O => \N__20915\,
            I => \N__20912\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__20912\,
            I => \tok.n12\
        );

    \I__4437\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20903\
        );

    \I__4436\ : InMux
    port map (
            O => \N__20908\,
            I => \N__20903\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__20903\,
            I => uart_rx_data_7
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__4433\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__20894\,
            I => \tok.n177\
        );

    \I__4431\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__20888\,
            I => \N__20885\
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__20885\,
            I => \tok.n17_adj_812\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__4427\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__20876\,
            I => \tok.n9_adj_838\
        );

    \I__4425\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__4423\ : Span4Mux_v
    port map (
            O => \N__20867\,
            I => \N__20864\
        );

    \I__4422\ : Odrv4
    port map (
            O => \N__20864\,
            I => \tok.n23_adj_682\
        );

    \I__4421\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20858\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__20858\,
            I => \tok.n25\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__20855\,
            I => \tok.n4_cascade_\
        );

    \I__4418\ : InMux
    port map (
            O => \N__20852\,
            I => \N__20849\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__20849\,
            I => \tok.n5350\
        );

    \I__4416\ : InMux
    port map (
            O => \N__20846\,
            I => \tok.n4807\
        );

    \I__4415\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20833\
        );

    \I__4414\ : InMux
    port map (
            O => \N__20842\,
            I => \N__20833\
        );

    \I__4413\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20830\
        );

    \I__4412\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20827\
        );

    \I__4411\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20822\
        );

    \I__4410\ : InMux
    port map (
            O => \N__20838\,
            I => \N__20822\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20813\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__20830\,
            I => \N__20813\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__20827\,
            I => \N__20813\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__20822\,
            I => \N__20813\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__4404\ : Span4Mux_h
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__20807\,
            I => \tok.n20_adj_663\
        );

    \I__4402\ : InMux
    port map (
            O => \N__20804\,
            I => \tok.n4808\
        );

    \I__4401\ : InMux
    port map (
            O => \N__20801\,
            I => \tok.n4809\
        );

    \I__4400\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20795\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__20795\,
            I => \N__20792\
        );

    \I__4398\ : Odrv4
    port map (
            O => \N__20792\,
            I => \tok.n10_adj_738\
        );

    \I__4397\ : InMux
    port map (
            O => \N__20789\,
            I => \tok.n4810\
        );

    \I__4396\ : InMux
    port map (
            O => \N__20786\,
            I => \tok.n4811\
        );

    \I__4395\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__4393\ : Span4Mux_v
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__20774\,
            I => \tok.n10_adj_768\
        );

    \I__4391\ : InMux
    port map (
            O => \N__20771\,
            I => \tok.n4812\
        );

    \I__4390\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20757\
        );

    \I__4389\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20757\
        );

    \I__4388\ : InMux
    port map (
            O => \N__20766\,
            I => \N__20752\
        );

    \I__4387\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20752\
        );

    \I__4386\ : SRMux
    port map (
            O => \N__20764\,
            I => \N__20745\
        );

    \I__4385\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20740\
        );

    \I__4384\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20740\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__20757\,
            I => \N__20737\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__20752\,
            I => \N__20734\
        );

    \I__4381\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20725\
        );

    \I__4380\ : InMux
    port map (
            O => \N__20750\,
            I => \N__20725\
        );

    \I__4379\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20725\
        );

    \I__4378\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20725\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__20745\,
            I => \N__20722\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__20740\,
            I => \N__20713\
        );

    \I__4375\ : Span4Mux_v
    port map (
            O => \N__20737\,
            I => \N__20713\
        );

    \I__4374\ : Span4Mux_v
    port map (
            O => \N__20734\,
            I => \N__20713\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__20725\,
            I => \N__20713\
        );

    \I__4372\ : Span4Mux_v
    port map (
            O => \N__20722\,
            I => \N__20710\
        );

    \I__4371\ : Span4Mux_h
    port map (
            O => \N__20713\,
            I => \N__20707\
        );

    \I__4370\ : Odrv4
    port map (
            O => \N__20710\,
            I => \tok.write_flag\
        );

    \I__4369\ : Odrv4
    port map (
            O => \N__20707\,
            I => \tok.write_flag\
        );

    \I__4368\ : InMux
    port map (
            O => \N__20702\,
            I => \tok.n4813\
        );

    \I__4367\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20696\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__20696\,
            I => \N__20693\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__20693\,
            I => \N__20690\
        );

    \I__4364\ : Span4Mux_v
    port map (
            O => \N__20690\,
            I => \N__20687\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__20687\,
            I => \tok.n5516\
        );

    \I__4362\ : InMux
    port map (
            O => \N__20684\,
            I => \N__20681\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__20681\,
            I => \N__20678\
        );

    \I__4360\ : Span4Mux_v
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__4359\ : Sp12to4
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__4358\ : Odrv12
    port map (
            O => \N__20672\,
            I => \tok.n18_adj_739\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__20669\,
            I => \tok.n12_adj_737_cascade_\
        );

    \I__4356\ : InMux
    port map (
            O => \N__20666\,
            I => \bfn_9_6_0_\
        );

    \I__4355\ : InMux
    port map (
            O => \N__20663\,
            I => \tok.n4799\
        );

    \I__4354\ : InMux
    port map (
            O => \N__20660\,
            I => \tok.n4800\
        );

    \I__4353\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20654\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__20654\,
            I => \N__20651\
        );

    \I__4351\ : Span4Mux_h
    port map (
            O => \N__20651\,
            I => \N__20648\
        );

    \I__4350\ : Odrv4
    port map (
            O => \N__20648\,
            I => \tok.n22_adj_829\
        );

    \I__4349\ : InMux
    port map (
            O => \N__20645\,
            I => \tok.n4801\
        );

    \I__4348\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20639\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__20639\,
            I => \N__20636\
        );

    \I__4346\ : Span4Mux_h
    port map (
            O => \N__20636\,
            I => \N__20633\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__20633\,
            I => \tok.n10_adj_827\
        );

    \I__4344\ : InMux
    port map (
            O => \N__20630\,
            I => \tok.n4802\
        );

    \I__4343\ : InMux
    port map (
            O => \N__20627\,
            I => \tok.n4803\
        );

    \I__4342\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20621\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__20621\,
            I => \tok.n10_adj_820\
        );

    \I__4340\ : InMux
    port map (
            O => \N__20618\,
            I => \tok.n4804\
        );

    \I__4339\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__20612\,
            I => \tok.n10_adj_653\
        );

    \I__4337\ : InMux
    port map (
            O => \N__20609\,
            I => \tok.n4805\
        );

    \I__4336\ : InMux
    port map (
            O => \N__20606\,
            I => \bfn_9_7_0_\
        );

    \I__4335\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20599\
        );

    \I__4334\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20596\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__20599\,
            I => \N__20593\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__20596\,
            I => \tok.A_stk.tail_86\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__20593\,
            I => \tok.A_stk.tail_86\
        );

    \I__4330\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20584\
        );

    \I__4329\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20581\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__20584\,
            I => \tok.A_stk.tail_55\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__20581\,
            I => \tok.A_stk.tail_55\
        );

    \I__4326\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20572\
        );

    \I__4325\ : InMux
    port map (
            O => \N__20575\,
            I => \N__20569\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__20572\,
            I => \tok.A_stk.tail_39\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__20569\,
            I => \tok.A_stk.tail_39\
        );

    \I__4322\ : InMux
    port map (
            O => \N__20564\,
            I => \N__20561\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__20561\,
            I => \N__20557\
        );

    \I__4320\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20554\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__20557\,
            I => \tok.A_stk.tail_83\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__20554\,
            I => \tok.A_stk.tail_83\
        );

    \I__4317\ : InMux
    port map (
            O => \N__20549\,
            I => \N__20545\
        );

    \I__4316\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20542\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__20545\,
            I => \tok.A_stk.tail_4\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__20542\,
            I => \tok.A_stk.tail_4\
        );

    \I__4313\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20531\
        );

    \I__4312\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20531\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__20531\,
            I => \tok.A_stk.tail_6\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__20528\,
            I => \N__20525\
        );

    \I__4309\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20521\
        );

    \I__4308\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20518\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__20521\,
            I => \tok.A_stk.tail_54\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__20518\,
            I => \tok.A_stk.tail_54\
        );

    \I__4305\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20507\
        );

    \I__4304\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20507\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__20507\,
            I => \tok.A_stk.tail_22\
        );

    \I__4302\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20501\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__20501\,
            I => \N__20497\
        );

    \I__4300\ : InMux
    port map (
            O => \N__20500\,
            I => \N__20494\
        );

    \I__4299\ : Odrv4
    port map (
            O => \N__20497\,
            I => \tok.A_stk.tail_38\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__20494\,
            I => \tok.A_stk.tail_38\
        );

    \I__4297\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20485\
        );

    \I__4296\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20482\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__20485\,
            I => \tok.A_stk.tail_23\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__20482\,
            I => \tok.A_stk.tail_23\
        );

    \I__4293\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20474\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__20474\,
            I => \N__20471\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__20471\,
            I => \tok.n3_adj_692\
        );

    \I__4290\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20465\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__20465\,
            I => \N__20461\
        );

    \I__4288\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20458\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__20461\,
            I => tail_100
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__20458\,
            I => tail_100
        );

    \I__4285\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20450\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__20450\,
            I => \N__20446\
        );

    \I__4283\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20443\
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__20446\,
            I => tail_116
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__20443\,
            I => tail_116
        );

    \I__4280\ : InMux
    port map (
            O => \N__20438\,
            I => \N__20434\
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__20437\,
            I => \N__20431\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__20434\,
            I => \N__20428\
        );

    \I__4277\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20425\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__20428\,
            I => tail_114
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__20425\,
            I => tail_114
        );

    \I__4274\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20416\
        );

    \I__4273\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20413\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__20416\,
            I => \N__20410\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__20413\,
            I => tail_98
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__20410\,
            I => tail_98
        );

    \I__4269\ : CascadeMux
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__4268\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20396\
        );

    \I__4267\ : InMux
    port map (
            O => \N__20401\,
            I => \N__20396\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__20396\,
            I => \tok.A_stk.tail_82\
        );

    \I__4265\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20389\
        );

    \I__4264\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20386\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__20389\,
            I => \tok.A_stk.tail_72\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__20386\,
            I => \tok.A_stk.tail_72\
        );

    \I__4261\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20377\
        );

    \I__4260\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20374\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__20377\,
            I => \N__20371\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__20374\,
            I => tail_102
        );

    \I__4257\ : Odrv12
    port map (
            O => \N__20371\,
            I => tail_102
        );

    \I__4256\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20360\
        );

    \I__4255\ : InMux
    port map (
            O => \N__20365\,
            I => \N__20360\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__20360\,
            I => \tok.A_stk.tail_70\
        );

    \I__4253\ : InMux
    port map (
            O => \N__20357\,
            I => \N__20354\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__20354\,
            I => \tok.n209\
        );

    \I__4251\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__4249\ : Odrv12
    port map (
            O => \N__20345\,
            I => \tok.n14_adj_658\
        );

    \I__4248\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__20336\,
            I => \tok.n2_adj_775\
        );

    \I__4245\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20329\
        );

    \I__4244\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20326\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__20329\,
            I => tail_118
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__20326\,
            I => tail_118
        );

    \I__4241\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20318\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__20318\,
            I => \tok.n14_adj_764\
        );

    \I__4239\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20304\
        );

    \I__4238\ : InMux
    port map (
            O => \N__20314\,
            I => \N__20304\
        );

    \I__4237\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20304\
        );

    \I__4236\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20299\
        );

    \I__4235\ : InMux
    port map (
            O => \N__20311\,
            I => \N__20299\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__20304\,
            I => \N__20286\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__20299\,
            I => \N__20286\
        );

    \I__4232\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20281\
        );

    \I__4231\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20281\
        );

    \I__4230\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20273\
        );

    \I__4229\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20254\
        );

    \I__4228\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20254\
        );

    \I__4227\ : InMux
    port map (
            O => \N__20293\,
            I => \N__20254\
        );

    \I__4226\ : InMux
    port map (
            O => \N__20292\,
            I => \N__20254\
        );

    \I__4225\ : InMux
    port map (
            O => \N__20291\,
            I => \N__20254\
        );

    \I__4224\ : Span4Mux_v
    port map (
            O => \N__20286\,
            I => \N__20249\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__20281\,
            I => \N__20249\
        );

    \I__4222\ : CascadeMux
    port map (
            O => \N__20280\,
            I => \N__20246\
        );

    \I__4221\ : CascadeMux
    port map (
            O => \N__20279\,
            I => \N__20241\
        );

    \I__4220\ : InMux
    port map (
            O => \N__20278\,
            I => \N__20233\
        );

    \I__4219\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20233\
        );

    \I__4218\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20224\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__20273\,
            I => \N__20221\
        );

    \I__4216\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20218\
        );

    \I__4215\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20213\
        );

    \I__4214\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20213\
        );

    \I__4213\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20208\
        );

    \I__4212\ : InMux
    port map (
            O => \N__20268\,
            I => \N__20208\
        );

    \I__4211\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20201\
        );

    \I__4210\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20201\
        );

    \I__4209\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20201\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__20254\,
            I => \N__20196\
        );

    \I__4207\ : Span4Mux_h
    port map (
            O => \N__20249\,
            I => \N__20196\
        );

    \I__4206\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20183\
        );

    \I__4205\ : InMux
    port map (
            O => \N__20245\,
            I => \N__20183\
        );

    \I__4204\ : InMux
    port map (
            O => \N__20244\,
            I => \N__20183\
        );

    \I__4203\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20183\
        );

    \I__4202\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20183\
        );

    \I__4201\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20178\
        );

    \I__4200\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20178\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__20233\,
            I => \N__20175\
        );

    \I__4198\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20172\
        );

    \I__4197\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20169\
        );

    \I__4196\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20159\
        );

    \I__4195\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20156\
        );

    \I__4194\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20151\
        );

    \I__4193\ : InMux
    port map (
            O => \N__20227\,
            I => \N__20151\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__20224\,
            I => \N__20146\
        );

    \I__4191\ : Span4Mux_v
    port map (
            O => \N__20221\,
            I => \N__20146\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__20218\,
            I => \N__20140\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__20213\,
            I => \N__20140\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__20208\,
            I => \N__20133\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__20201\,
            I => \N__20133\
        );

    \I__4186\ : Span4Mux_v
    port map (
            O => \N__20196\,
            I => \N__20133\
        );

    \I__4185\ : CascadeMux
    port map (
            O => \N__20195\,
            I => \N__20129\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__20194\,
            I => \N__20126\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__20183\,
            I => \N__20115\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20108\
        );

    \I__4181\ : Span4Mux_h
    port map (
            O => \N__20175\,
            I => \N__20108\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__20172\,
            I => \N__20108\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__20169\,
            I => \N__20105\
        );

    \I__4178\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20090\
        );

    \I__4177\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20090\
        );

    \I__4176\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20090\
        );

    \I__4175\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20090\
        );

    \I__4174\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20090\
        );

    \I__4173\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20090\
        );

    \I__4172\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20090\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__20159\,
            I => \N__20085\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__20156\,
            I => \N__20085\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__20151\,
            I => \N__20082\
        );

    \I__4168\ : Span4Mux_h
    port map (
            O => \N__20146\,
            I => \N__20079\
        );

    \I__4167\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20076\
        );

    \I__4166\ : Span4Mux_h
    port map (
            O => \N__20140\,
            I => \N__20071\
        );

    \I__4165\ : Span4Mux_v
    port map (
            O => \N__20133\,
            I => \N__20071\
        );

    \I__4164\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20060\
        );

    \I__4163\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20060\
        );

    \I__4162\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20060\
        );

    \I__4161\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20060\
        );

    \I__4160\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20060\
        );

    \I__4159\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20051\
        );

    \I__4158\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20051\
        );

    \I__4157\ : InMux
    port map (
            O => \N__20121\,
            I => \N__20051\
        );

    \I__4156\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20051\
        );

    \I__4155\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20046\
        );

    \I__4154\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20046\
        );

    \I__4153\ : Span4Mux_h
    port map (
            O => \N__20115\,
            I => \N__20043\
        );

    \I__4152\ : Span4Mux_v
    port map (
            O => \N__20108\,
            I => \N__20034\
        );

    \I__4151\ : Span4Mux_h
    port map (
            O => \N__20105\,
            I => \N__20034\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__20090\,
            I => \N__20034\
        );

    \I__4149\ : Span4Mux_h
    port map (
            O => \N__20085\,
            I => \N__20034\
        );

    \I__4148\ : Span12Mux_s11_v
    port map (
            O => \N__20082\,
            I => \N__20031\
        );

    \I__4147\ : Odrv4
    port map (
            O => \N__20079\,
            I => \tok.T_0\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__20076\,
            I => \tok.T_0\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__20071\,
            I => \tok.T_0\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__20060\,
            I => \tok.T_0\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__20051\,
            I => \tok.T_0\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__20046\,
            I => \tok.T_0\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__20043\,
            I => \tok.T_0\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__20034\,
            I => \tok.T_0\
        );

    \I__4139\ : Odrv12
    port map (
            O => \N__20031\,
            I => \tok.T_0\
        );

    \I__4138\ : InMux
    port map (
            O => \N__20012\,
            I => \N__20009\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__20009\,
            I => \N__20006\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__20006\,
            I => \tok.n10_adj_858\
        );

    \I__4135\ : InMux
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__20000\,
            I => \N__19997\
        );

    \I__4133\ : Span4Mux_h
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__4132\ : Span4Mux_h
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__4131\ : Odrv4
    port map (
            O => \N__19991\,
            I => \tok.table_rd_13\
        );

    \I__4130\ : InMux
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__4128\ : Odrv12
    port map (
            O => \N__19982\,
            I => \tok.n5_adj_732\
        );

    \I__4127\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__19976\,
            I => \tok.n12_adj_779\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__19973\,
            I => \tok.n14_adj_776_cascade_\
        );

    \I__4124\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__19967\,
            I => \tok.n13_adj_780\
        );

    \I__4122\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \tok.n20_adj_784_cascade_\
        );

    \I__4121\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__19958\,
            I => \tok.n9_adj_781\
        );

    \I__4119\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19952\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__4117\ : Odrv12
    port map (
            O => \N__19949\,
            I => \tok.n5_adj_713\
        );

    \I__4116\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__4114\ : Span4Mux_v
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__4113\ : Span4Mux_h
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__4112\ : Span4Mux_h
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__19931\,
            I => \tok.table_rd_15\
        );

    \I__4110\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__19925\,
            I => \tok.n16_adj_782\
        );

    \I__4108\ : CascadeMux
    port map (
            O => \N__19922\,
            I => \tok.n10_adj_700_cascade_\
        );

    \I__4107\ : InMux
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__19916\,
            I => \tok.n5536\
        );

    \I__4105\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__19910\,
            I => \tok.n11_adj_730\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__19907\,
            I => \tok.n26_cascade_\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__19904\,
            I => \N__19898\
        );

    \I__4101\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19892\
        );

    \I__4100\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19889\
        );

    \I__4099\ : InMux
    port map (
            O => \N__19901\,
            I => \N__19885\
        );

    \I__4098\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19882\
        );

    \I__4097\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19879\
        );

    \I__4096\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19876\
        );

    \I__4095\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19873\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__19892\,
            I => \N__19870\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__19889\,
            I => \N__19867\
        );

    \I__4092\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19864\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__19885\,
            I => \N__19861\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__19882\,
            I => \N__19856\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__19879\,
            I => \N__19856\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__19876\,
            I => \N__19853\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__19873\,
            I => \N__19848\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__19870\,
            I => \N__19848\
        );

    \I__4085\ : Span4Mux_v
    port map (
            O => \N__19867\,
            I => \N__19845\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__19864\,
            I => \N__19842\
        );

    \I__4083\ : Span4Mux_v
    port map (
            O => \N__19861\,
            I => \N__19839\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__19856\,
            I => \N__19836\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__19853\,
            I => \N__19831\
        );

    \I__4080\ : Span4Mux_v
    port map (
            O => \N__19848\,
            I => \N__19831\
        );

    \I__4079\ : Span4Mux_h
    port map (
            O => \N__19845\,
            I => \N__19828\
        );

    \I__4078\ : Span4Mux_h
    port map (
            O => \N__19842\,
            I => \N__19823\
        );

    \I__4077\ : Span4Mux_h
    port map (
            O => \N__19839\,
            I => \N__19823\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__19836\,
            I => \N__19818\
        );

    \I__4075\ : Span4Mux_h
    port map (
            O => \N__19831\,
            I => \N__19818\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__19828\,
            I => \tok.tc__7__N_134\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__19823\,
            I => \tok.tc__7__N_134\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__19818\,
            I => \tok.tc__7__N_134\
        );

    \I__4071\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__19808\,
            I => \tok.n25_adj_710\
        );

    \I__4069\ : InMux
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__19799\,
            I => \tok.n28_adj_708\
        );

    \I__4066\ : InMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__19793\,
            I => \tok.n27_adj_709\
        );

    \I__4064\ : InMux
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__4062\ : Span4Mux_v
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__4061\ : Span4Mux_h
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__19778\,
            I => \tok.n16_adj_810\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__19775\,
            I => \tok.n14_adj_841_cascade_\
        );

    \I__4058\ : InMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__4056\ : Span4Mux_h
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__19763\,
            I => \tok.n5571\
        );

    \I__4054\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__19757\,
            I => \tok.n5569\
        );

    \I__4052\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__19748\,
            I => \tok.n45_adj_849\
        );

    \I__4049\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19739\
        );

    \I__4048\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19739\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__19739\,
            I => \N__19735\
        );

    \I__4046\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19732\
        );

    \I__4045\ : Span4Mux_v
    port map (
            O => \N__19735\,
            I => \N__19727\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__19732\,
            I => \N__19727\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__19727\,
            I => \tok.n4848\
        );

    \I__4042\ : InMux
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__4040\ : Span4Mux_h
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__4039\ : Span4Mux_h
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__19712\,
            I => \tok.table_rd_9\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__19709\,
            I => \tok.n45_cascade_\
        );

    \I__4036\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__19703\,
            I => \tok.n39\
        );

    \I__4034\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19694\
        );

    \I__4033\ : InMux
    port map (
            O => \N__19699\,
            I => \N__19694\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__19694\,
            I => \N__19690\
        );

    \I__4031\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19687\
        );

    \I__4030\ : Span4Mux_v
    port map (
            O => \N__19690\,
            I => \N__19682\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__19687\,
            I => \N__19682\
        );

    \I__4028\ : Span4Mux_h
    port map (
            O => \N__19682\,
            I => \N__19677\
        );

    \I__4027\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19672\
        );

    \I__4026\ : InMux
    port map (
            O => \N__19680\,
            I => \N__19672\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__19677\,
            I => \tok.n11_adj_680\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__19672\,
            I => \tok.n11_adj_680\
        );

    \I__4023\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__4021\ : Span4Mux_v
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__4020\ : Span4Mux_h
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__4019\ : Span4Mux_h
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__4018\ : Span4Mux_s0_h
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__19649\,
            I => \tok.table_rd_10\
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__4015\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19637\
        );

    \I__4014\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19637\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__19637\,
            I => \tok.n14_adj_679\
        );

    \I__4012\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__19631\,
            I => \tok.n45_adj_696\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__19628\,
            I => \tok.n39_adj_697_cascade_\
        );

    \I__4009\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__19622\,
            I => \tok.n5_adj_734\
        );

    \I__4007\ : InMux
    port map (
            O => \N__19619\,
            I => \tok.n4795\
        );

    \I__4006\ : InMux
    port map (
            O => \N__19616\,
            I => \tok.n4796\
        );

    \I__4005\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__4003\ : Odrv4
    port map (
            O => \N__19607\,
            I => \tok.n5_adj_716\
        );

    \I__4002\ : InMux
    port map (
            O => \N__19604\,
            I => \tok.n4797\
        );

    \I__4001\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19579\
        );

    \I__4000\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19579\
        );

    \I__3999\ : InMux
    port map (
            O => \N__19599\,
            I => \N__19579\
        );

    \I__3998\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19568\
        );

    \I__3997\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19568\
        );

    \I__3996\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19568\
        );

    \I__3995\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19568\
        );

    \I__3994\ : InMux
    port map (
            O => \N__19594\,
            I => \N__19568\
        );

    \I__3993\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19561\
        );

    \I__3992\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19561\
        );

    \I__3991\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19561\
        );

    \I__3990\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19550\
        );

    \I__3989\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19550\
        );

    \I__3988\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19550\
        );

    \I__3987\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19550\
        );

    \I__3986\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19550\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__19579\,
            I => \N__19545\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__19568\,
            I => \N__19545\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__19561\,
            I => \N__19540\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__19550\,
            I => \N__19540\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__19545\,
            I => \N__19537\
        );

    \I__3980\ : Span4Mux_v
    port map (
            O => \N__19540\,
            I => \N__19534\
        );

    \I__3979\ : Span4Mux_h
    port map (
            O => \N__19537\,
            I => \N__19529\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__19534\,
            I => \N__19529\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__19529\,
            I => \tok.n399\
        );

    \I__3976\ : InMux
    port map (
            O => \N__19526\,
            I => \tok.n4798\
        );

    \I__3975\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__19520\,
            I => \tok.n8_adj_837\
        );

    \I__3973\ : InMux
    port map (
            O => \N__19517\,
            I => \N__19514\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__19514\,
            I => \tok.n5574\
        );

    \I__3971\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19507\
        );

    \I__3970\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19504\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__19507\,
            I => \tok.n5334\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__19504\,
            I => \tok.n5334\
        );

    \I__3967\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__3965\ : Span4Mux_v
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__19490\,
            I => \tok.n5254\
        );

    \I__3963\ : CascadeMux
    port map (
            O => \N__19487\,
            I => \tok.n5414_cascade_\
        );

    \I__3962\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__19481\,
            I => \tok.n8_adj_767\
        );

    \I__3960\ : CascadeMux
    port map (
            O => \N__19478\,
            I => \tok.n904_cascade_\
        );

    \I__3959\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19472\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__19472\,
            I => \N__19469\
        );

    \I__3957\ : Span4Mux_v
    port map (
            O => \N__19469\,
            I => \N__19466\
        );

    \I__3956\ : Span4Mux_s2_v
    port map (
            O => \N__19466\,
            I => \N__19463\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__19463\,
            I => \tok.n11_adj_840\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__19460\,
            I => \tok.n5346_cascade_\
        );

    \I__3953\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19454\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__3951\ : Sp12to4
    port map (
            O => \N__19451\,
            I => \N__19448\
        );

    \I__3950\ : Odrv12
    port map (
            O => \N__19448\,
            I => \tok.n4_adj_806\
        );

    \I__3949\ : InMux
    port map (
            O => \N__19445\,
            I => \tok.n4786\
        );

    \I__3948\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19439\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__19439\,
            I => \tok.n5564\
        );

    \I__3946\ : InMux
    port map (
            O => \N__19436\,
            I => \tok.n4787\
        );

    \I__3945\ : InMux
    port map (
            O => \N__19433\,
            I => \tok.n4788\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__3943\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__19424\,
            I => \tok.n5554\
        );

    \I__3941\ : InMux
    port map (
            O => \N__19421\,
            I => \tok.n4789\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__3939\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__19412\,
            I => \N__19409\
        );

    \I__3937\ : Odrv12
    port map (
            O => \N__19409\,
            I => \tok.n5549\
        );

    \I__3936\ : InMux
    port map (
            O => \N__19406\,
            I => \tok.n4790\
        );

    \I__3935\ : InMux
    port map (
            O => \N__19403\,
            I => \bfn_8_8_0_\
        );

    \I__3934\ : InMux
    port map (
            O => \N__19400\,
            I => \tok.n4792\
        );

    \I__3933\ : InMux
    port map (
            O => \N__19397\,
            I => \tok.n4793\
        );

    \I__3932\ : InMux
    port map (
            O => \N__19394\,
            I => \tok.n4794\
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__19391\,
            I => \tok.n13_adj_654_cascade_\
        );

    \I__3930\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__19385\,
            I => \tok.n5547\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__19382\,
            I => \tok.n5546_cascade_\
        );

    \I__3927\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__3925\ : Span4Mux_h
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__3924\ : Odrv4
    port map (
            O => \N__19370\,
            I => \tok.n14\
        );

    \I__3923\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__19364\,
            I => \tok.n17\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__19361\,
            I => \tok.n13_adj_641_cascade_\
        );

    \I__3920\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__19355\,
            I => \tok.n5552\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__19352\,
            I => \tok.n5551_cascade_\
        );

    \I__3917\ : InMux
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__19343\,
            I => \tok.n5465\
        );

    \I__3914\ : InMux
    port map (
            O => \N__19340\,
            I => \tok.n4784\
        );

    \I__3913\ : InMux
    port map (
            O => \N__19337\,
            I => \tok.n4785\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__19334\,
            I => \N__19330\
        );

    \I__3911\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19325\
        );

    \I__3910\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19325\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__19325\,
            I => \N__19320\
        );

    \I__3908\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19315\
        );

    \I__3907\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19315\
        );

    \I__3906\ : Span12Mux_s4_v
    port map (
            O => \N__19320\,
            I => \N__19312\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__19315\,
            I => \tok.n9_adj_786\
        );

    \I__3904\ : Odrv12
    port map (
            O => \N__19312\,
            I => \tok.n9_adj_786\
        );

    \I__3903\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19304\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__3901\ : Span4Mux_v
    port map (
            O => \N__19301\,
            I => \N__19297\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__19300\,
            I => \N__19294\
        );

    \I__3899\ : Span4Mux_h
    port map (
            O => \N__19297\,
            I => \N__19291\
        );

    \I__3898\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19288\
        );

    \I__3897\ : Odrv4
    port map (
            O => \N__19291\,
            I => \tok.table_rd_7\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__19288\,
            I => \tok.table_rd_7\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__19283\,
            I => \tok.n5548_cascade_\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__19280\,
            I => \tok.n285_cascade_\
        );

    \I__3893\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__19274\,
            I => \N__19271\
        );

    \I__3891\ : Span4Mux_v
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__3890\ : Span4Mux_h
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__3889\ : Odrv4
    port map (
            O => \N__19265\,
            I => \tok.n12_adj_824\
        );

    \I__3888\ : CascadeMux
    port map (
            O => \N__19262\,
            I => \tok.n1_adj_862_cascade_\
        );

    \I__3887\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19252\
        );

    \I__3886\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19247\
        );

    \I__3885\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19247\
        );

    \I__3884\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19241\
        );

    \I__3883\ : CascadeMux
    port map (
            O => \N__19255\,
            I => \N__19233\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__19252\,
            I => \N__19227\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__19247\,
            I => \N__19227\
        );

    \I__3880\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19224\
        );

    \I__3879\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19221\
        );

    \I__3878\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19218\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__19241\,
            I => \N__19211\
        );

    \I__3876\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19208\
        );

    \I__3875\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19205\
        );

    \I__3874\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19200\
        );

    \I__3873\ : InMux
    port map (
            O => \N__19237\,
            I => \N__19200\
        );

    \I__3872\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19191\
        );

    \I__3871\ : InMux
    port map (
            O => \N__19233\,
            I => \N__19191\
        );

    \I__3870\ : InMux
    port map (
            O => \N__19232\,
            I => \N__19191\
        );

    \I__3869\ : Span4Mux_v
    port map (
            O => \N__19227\,
            I => \N__19186\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__19224\,
            I => \N__19186\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__19221\,
            I => \N__19183\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__19218\,
            I => \N__19180\
        );

    \I__3865\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19175\
        );

    \I__3864\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19175\
        );

    \I__3863\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19172\
        );

    \I__3862\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19169\
        );

    \I__3861\ : Span4Mux_v
    port map (
            O => \N__19211\,
            I => \N__19163\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__19208\,
            I => \N__19158\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__19205\,
            I => \N__19158\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__19200\,
            I => \N__19155\
        );

    \I__3857\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19148\
        );

    \I__3856\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19148\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__19191\,
            I => \N__19143\
        );

    \I__3854\ : Span4Mux_h
    port map (
            O => \N__19186\,
            I => \N__19143\
        );

    \I__3853\ : Span4Mux_h
    port map (
            O => \N__19183\,
            I => \N__19140\
        );

    \I__3852\ : Span4Mux_v
    port map (
            O => \N__19180\,
            I => \N__19135\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__19175\,
            I => \N__19135\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__19172\,
            I => \N__19130\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__19169\,
            I => \N__19130\
        );

    \I__3848\ : InMux
    port map (
            O => \N__19168\,
            I => \N__19125\
        );

    \I__3847\ : InMux
    port map (
            O => \N__19167\,
            I => \N__19125\
        );

    \I__3846\ : InMux
    port map (
            O => \N__19166\,
            I => \N__19122\
        );

    \I__3845\ : Span4Mux_v
    port map (
            O => \N__19163\,
            I => \N__19119\
        );

    \I__3844\ : Span4Mux_v
    port map (
            O => \N__19158\,
            I => \N__19116\
        );

    \I__3843\ : Span12Mux_s10_v
    port map (
            O => \N__19155\,
            I => \N__19113\
        );

    \I__3842\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19110\
        );

    \I__3841\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19107\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__19148\,
            I => \N__19102\
        );

    \I__3839\ : Span4Mux_v
    port map (
            O => \N__19143\,
            I => \N__19102\
        );

    \I__3838\ : Span4Mux_v
    port map (
            O => \N__19140\,
            I => \N__19097\
        );

    \I__3837\ : Span4Mux_h
    port map (
            O => \N__19135\,
            I => \N__19097\
        );

    \I__3836\ : Span4Mux_s3_v
    port map (
            O => \N__19130\,
            I => \N__19092\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__19125\,
            I => \N__19092\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__19122\,
            I => \tok.T_6\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__19119\,
            I => \tok.T_6\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__19116\,
            I => \tok.T_6\
        );

    \I__3831\ : Odrv12
    port map (
            O => \N__19113\,
            I => \tok.T_6\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__19110\,
            I => \tok.T_6\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__19107\,
            I => \tok.T_6\
        );

    \I__3828\ : Odrv4
    port map (
            O => \N__19102\,
            I => \tok.T_6\
        );

    \I__3827\ : Odrv4
    port map (
            O => \N__19097\,
            I => \tok.T_6\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__19092\,
            I => \tok.T_6\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__19073\,
            I => \N__19067\
        );

    \I__3824\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19061\
        );

    \I__3823\ : InMux
    port map (
            O => \N__19071\,
            I => \N__19061\
        );

    \I__3822\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19039\
        );

    \I__3821\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19032\
        );

    \I__3820\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19032\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__19061\,
            I => \N__19029\
        );

    \I__3818\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19024\
        );

    \I__3817\ : InMux
    port map (
            O => \N__19059\,
            I => \N__19024\
        );

    \I__3816\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19019\
        );

    \I__3815\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19019\
        );

    \I__3814\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19010\
        );

    \I__3813\ : InMux
    port map (
            O => \N__19055\,
            I => \N__19010\
        );

    \I__3812\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19010\
        );

    \I__3811\ : InMux
    port map (
            O => \N__19053\,
            I => \N__19007\
        );

    \I__3810\ : InMux
    port map (
            O => \N__19052\,
            I => \N__19004\
        );

    \I__3809\ : InMux
    port map (
            O => \N__19051\,
            I => \N__18999\
        );

    \I__3808\ : InMux
    port map (
            O => \N__19050\,
            I => \N__18999\
        );

    \I__3807\ : InMux
    port map (
            O => \N__19049\,
            I => \N__18994\
        );

    \I__3806\ : InMux
    port map (
            O => \N__19048\,
            I => \N__18994\
        );

    \I__3805\ : InMux
    port map (
            O => \N__19047\,
            I => \N__18987\
        );

    \I__3804\ : InMux
    port map (
            O => \N__19046\,
            I => \N__18987\
        );

    \I__3803\ : InMux
    port map (
            O => \N__19045\,
            I => \N__18987\
        );

    \I__3802\ : InMux
    port map (
            O => \N__19044\,
            I => \N__18984\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__19043\,
            I => \N__18980\
        );

    \I__3800\ : InMux
    port map (
            O => \N__19042\,
            I => \N__18976\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__19039\,
            I => \N__18973\
        );

    \I__3798\ : InMux
    port map (
            O => \N__19038\,
            I => \N__18970\
        );

    \I__3797\ : InMux
    port map (
            O => \N__19037\,
            I => \N__18967\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__19032\,
            I => \N__18964\
        );

    \I__3795\ : Span4Mux_v
    port map (
            O => \N__19029\,
            I => \N__18955\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__19024\,
            I => \N__18955\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__19019\,
            I => \N__18955\
        );

    \I__3792\ : InMux
    port map (
            O => \N__19018\,
            I => \N__18950\
        );

    \I__3791\ : InMux
    port map (
            O => \N__19017\,
            I => \N__18950\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__19010\,
            I => \N__18947\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__19007\,
            I => \N__18942\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__19004\,
            I => \N__18942\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__18999\,
            I => \N__18937\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__18994\,
            I => \N__18937\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__18987\,
            I => \N__18932\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__18984\,
            I => \N__18932\
        );

    \I__3783\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18925\
        );

    \I__3782\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18925\
        );

    \I__3781\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18925\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__18976\,
            I => \N__18921\
        );

    \I__3779\ : Span4Mux_h
    port map (
            O => \N__18973\,
            I => \N__18918\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__18970\,
            I => \N__18915\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__18967\,
            I => \N__18910\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__18964\,
            I => \N__18910\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__18963\,
            I => \N__18905\
        );

    \I__3774\ : CascadeMux
    port map (
            O => \N__18962\,
            I => \N__18902\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__18955\,
            I => \N__18897\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__18950\,
            I => \N__18897\
        );

    \I__3771\ : Span4Mux_s3_h
    port map (
            O => \N__18947\,
            I => \N__18894\
        );

    \I__3770\ : Span4Mux_v
    port map (
            O => \N__18942\,
            I => \N__18891\
        );

    \I__3769\ : Span4Mux_v
    port map (
            O => \N__18937\,
            I => \N__18884\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__18932\,
            I => \N__18884\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__18925\,
            I => \N__18884\
        );

    \I__3766\ : InMux
    port map (
            O => \N__18924\,
            I => \N__18881\
        );

    \I__3765\ : Span4Mux_h
    port map (
            O => \N__18921\,
            I => \N__18876\
        );

    \I__3764\ : Span4Mux_v
    port map (
            O => \N__18918\,
            I => \N__18876\
        );

    \I__3763\ : Span4Mux_v
    port map (
            O => \N__18915\,
            I => \N__18871\
        );

    \I__3762\ : Span4Mux_h
    port map (
            O => \N__18910\,
            I => \N__18871\
        );

    \I__3761\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18866\
        );

    \I__3760\ : InMux
    port map (
            O => \N__18908\,
            I => \N__18866\
        );

    \I__3759\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18863\
        );

    \I__3758\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18860\
        );

    \I__3757\ : Span4Mux_v
    port map (
            O => \N__18897\,
            I => \N__18851\
        );

    \I__3756\ : Span4Mux_v
    port map (
            O => \N__18894\,
            I => \N__18851\
        );

    \I__3755\ : Span4Mux_h
    port map (
            O => \N__18891\,
            I => \N__18851\
        );

    \I__3754\ : Span4Mux_h
    port map (
            O => \N__18884\,
            I => \N__18851\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__18881\,
            I => \tok.T_4\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__18876\,
            I => \tok.T_4\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__18871\,
            I => \tok.T_4\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__18866\,
            I => \tok.T_4\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__18863\,
            I => \tok.T_4\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__18860\,
            I => \tok.T_4\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__18851\,
            I => \tok.T_4\
        );

    \I__3746\ : CascadeMux
    port map (
            O => \N__18836\,
            I => \N__18827\
        );

    \I__3745\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18822\
        );

    \I__3744\ : InMux
    port map (
            O => \N__18834\,
            I => \N__18822\
        );

    \I__3743\ : InMux
    port map (
            O => \N__18833\,
            I => \N__18819\
        );

    \I__3742\ : InMux
    port map (
            O => \N__18832\,
            I => \N__18808\
        );

    \I__3741\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18808\
        );

    \I__3740\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18808\
        );

    \I__3739\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18805\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__18822\,
            I => \N__18799\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__18819\,
            I => \N__18799\
        );

    \I__3736\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18792\
        );

    \I__3735\ : InMux
    port map (
            O => \N__18817\,
            I => \N__18792\
        );

    \I__3734\ : InMux
    port map (
            O => \N__18816\,
            I => \N__18792\
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__18815\,
            I => \N__18788\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__18808\,
            I => \N__18785\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__18805\,
            I => \N__18782\
        );

    \I__3730\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18779\
        );

    \I__3729\ : Span4Mux_v
    port map (
            O => \N__18799\,
            I => \N__18774\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__18792\,
            I => \N__18771\
        );

    \I__3727\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18766\
        );

    \I__3726\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18766\
        );

    \I__3725\ : Span4Mux_v
    port map (
            O => \N__18785\,
            I => \N__18762\
        );

    \I__3724\ : Span4Mux_v
    port map (
            O => \N__18782\,
            I => \N__18758\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__18779\,
            I => \N__18755\
        );

    \I__3722\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18750\
        );

    \I__3721\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18750\
        );

    \I__3720\ : Span4Mux_v
    port map (
            O => \N__18774\,
            I => \N__18743\
        );

    \I__3719\ : Span4Mux_v
    port map (
            O => \N__18771\,
            I => \N__18743\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__18766\,
            I => \N__18743\
        );

    \I__3717\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18740\
        );

    \I__3716\ : Span4Mux_h
    port map (
            O => \N__18762\,
            I => \N__18737\
        );

    \I__3715\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18734\
        );

    \I__3714\ : Span4Mux_v
    port map (
            O => \N__18758\,
            I => \N__18727\
        );

    \I__3713\ : Span4Mux_s3_v
    port map (
            O => \N__18755\,
            I => \N__18727\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__18750\,
            I => \N__18727\
        );

    \I__3711\ : Span4Mux_h
    port map (
            O => \N__18743\,
            I => \N__18724\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__18740\,
            I => \tok.T_5\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__18737\,
            I => \tok.T_5\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__18734\,
            I => \tok.T_5\
        );

    \I__3707\ : Odrv4
    port map (
            O => \N__18727\,
            I => \tok.T_5\
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__18724\,
            I => \tok.T_5\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__18713\,
            I => \tok.n6_adj_650_cascade_\
        );

    \I__3704\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18704\
        );

    \I__3703\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18704\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__18704\,
            I => \tok.A_stk.tail_68\
        );

    \I__3701\ : InMux
    port map (
            O => \N__18701\,
            I => \N__18695\
        );

    \I__3700\ : InMux
    port map (
            O => \N__18700\,
            I => \N__18695\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__18695\,
            I => \tok.A_stk.tail_52\
        );

    \I__3698\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18686\
        );

    \I__3697\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18686\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__18686\,
            I => \tok.A_stk.tail_36\
        );

    \I__3695\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18679\
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__18682\,
            I => \N__18676\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__18679\,
            I => \N__18673\
        );

    \I__3692\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18670\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__18673\,
            I => tail_119
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__18670\,
            I => tail_119
        );

    \I__3689\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18661\
        );

    \I__3688\ : InMux
    port map (
            O => \N__18664\,
            I => \N__18658\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__18661\,
            I => \tok.A_stk.tail_20\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__18658\,
            I => \tok.A_stk.tail_20\
        );

    \I__3685\ : InMux
    port map (
            O => \N__18653\,
            I => \N__18649\
        );

    \I__3684\ : InMux
    port map (
            O => \N__18652\,
            I => \N__18646\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__18649\,
            I => tail_103
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__18646\,
            I => tail_103
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__3680\ : InMux
    port map (
            O => \N__18638\,
            I => \N__18632\
        );

    \I__3679\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18632\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__18632\,
            I => \tok.A_stk.tail_71\
        );

    \I__3677\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18625\
        );

    \I__3676\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18622\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__18625\,
            I => \tok.A_stk.tail_87\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__18622\,
            I => \tok.A_stk.tail_87\
        );

    \I__3673\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18613\
        );

    \I__3672\ : InMux
    port map (
            O => \N__18616\,
            I => \N__18610\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__18613\,
            I => tail_120
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__18610\,
            I => tail_120
        );

    \I__3669\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18599\
        );

    \I__3668\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18599\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__18599\,
            I => \tok.A_stk.tail_88\
        );

    \I__3666\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__18593\,
            I => \N__18589\
        );

    \I__3664\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18586\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__18589\,
            I => tail_104
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__18586\,
            I => tail_104
        );

    \I__3661\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18575\
        );

    \I__3660\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18575\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__18575\,
            I => \tok.A_stk.tail_41\
        );

    \I__3658\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18566\
        );

    \I__3657\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18566\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__18566\,
            I => \tok.A_stk.tail_25\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__3654\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18554\
        );

    \I__3653\ : InMux
    port map (
            O => \N__18559\,
            I => \N__18554\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__18554\,
            I => \tok.A_stk.tail_9\
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__18551\,
            I => \N__18547\
        );

    \I__3650\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18544\
        );

    \I__3649\ : InMux
    port map (
            O => \N__18547\,
            I => \N__18541\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__18544\,
            I => tail_115
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__18541\,
            I => tail_115
        );

    \I__3646\ : InMux
    port map (
            O => \N__18536\,
            I => \N__18532\
        );

    \I__3645\ : InMux
    port map (
            O => \N__18535\,
            I => \N__18529\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__18532\,
            I => tail_99
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__18529\,
            I => tail_99
        );

    \I__3642\ : InMux
    port map (
            O => \N__18524\,
            I => \N__18520\
        );

    \I__3641\ : InMux
    port map (
            O => \N__18523\,
            I => \N__18517\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__18520\,
            I => \tok.A_stk.tail_84\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__18517\,
            I => \tok.A_stk.tail_84\
        );

    \I__3638\ : InMux
    port map (
            O => \N__18512\,
            I => \tok.n4765\
        );

    \I__3637\ : CascadeMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__3636\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__3634\ : Sp12to4
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__3633\ : Odrv12
    port map (
            O => \N__18497\,
            I => \tok.n210\
        );

    \I__3632\ : InMux
    port map (
            O => \N__18494\,
            I => \tok.n4766\
        );

    \I__3631\ : InMux
    port map (
            O => \N__18491\,
            I => \tok.n4767\
        );

    \I__3630\ : InMux
    port map (
            O => \N__18488\,
            I => \bfn_7_14_0_\
        );

    \I__3629\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__18482\,
            I => \N__18478\
        );

    \I__3627\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18475\
        );

    \I__3626\ : Odrv4
    port map (
            O => \N__18478\,
            I => tail_121
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__18475\,
            I => tail_121
        );

    \I__3624\ : InMux
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__3622\ : Span4Mux_h
    port map (
            O => \N__18464\,
            I => \N__18460\
        );

    \I__3621\ : InMux
    port map (
            O => \N__18463\,
            I => \N__18457\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__18460\,
            I => tail_105
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__18457\,
            I => tail_105
        );

    \I__3618\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18446\
        );

    \I__3617\ : InMux
    port map (
            O => \N__18451\,
            I => \N__18446\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__18446\,
            I => \tok.A_stk.tail_89\
        );

    \I__3615\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18437\
        );

    \I__3614\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18437\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__18437\,
            I => \tok.A_stk.tail_73\
        );

    \I__3612\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18428\
        );

    \I__3611\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18428\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__18428\,
            I => \tok.A_stk.tail_57\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__18425\,
            I => \tok.n82_cascade_\
        );

    \I__3608\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18415\
        );

    \I__3607\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18415\
        );

    \I__3606\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18411\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__18415\,
            I => \N__18408\
        );

    \I__3604\ : InMux
    port map (
            O => \N__18414\,
            I => \N__18405\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__18411\,
            I => \tok.n878\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__18408\,
            I => \tok.n878\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__18405\,
            I => \tok.n878\
        );

    \I__3600\ : InMux
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__3598\ : Span4Mux_h
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__18389\,
            I => \tok.n8_adj_846\
        );

    \I__3596\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18380\
        );

    \I__3595\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18380\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__3592\ : Span4Mux_v
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__18371\,
            I => \tok.n41\
        );

    \I__3590\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18362\
        );

    \I__3589\ : InMux
    port map (
            O => \N__18367\,
            I => \N__18362\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__18362\,
            I => \N__18347\
        );

    \I__3587\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18342\
        );

    \I__3586\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18342\
        );

    \I__3585\ : CascadeMux
    port map (
            O => \N__18359\,
            I => \N__18336\
        );

    \I__3584\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18331\
        );

    \I__3583\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18322\
        );

    \I__3582\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18322\
        );

    \I__3581\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18322\
        );

    \I__3580\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18322\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \N__18319\
        );

    \I__3578\ : InMux
    port map (
            O => \N__18352\,
            I => \N__18308\
        );

    \I__3577\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18308\
        );

    \I__3576\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18301\
        );

    \I__3575\ : Span4Mux_v
    port map (
            O => \N__18347\,
            I => \N__18296\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18296\
        );

    \I__3573\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18284\
        );

    \I__3572\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18284\
        );

    \I__3571\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18284\
        );

    \I__3570\ : InMux
    port map (
            O => \N__18336\,
            I => \N__18284\
        );

    \I__3569\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18276\
        );

    \I__3568\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18273\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__18331\,
            I => \N__18268\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__18322\,
            I => \N__18268\
        );

    \I__3565\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18263\
        );

    \I__3564\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18263\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__18317\,
            I => \N__18259\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__18316\,
            I => \N__18255\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__18315\,
            I => \N__18252\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__18314\,
            I => \N__18247\
        );

    \I__3559\ : InMux
    port map (
            O => \N__18313\,
            I => \N__18244\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__18308\,
            I => \N__18241\
        );

    \I__3557\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18232\
        );

    \I__3556\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18232\
        );

    \I__3555\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18232\
        );

    \I__3554\ : InMux
    port map (
            O => \N__18304\,
            I => \N__18232\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__18301\,
            I => \N__18229\
        );

    \I__3552\ : Span4Mux_h
    port map (
            O => \N__18296\,
            I => \N__18226\
        );

    \I__3551\ : InMux
    port map (
            O => \N__18295\,
            I => \N__18223\
        );

    \I__3550\ : InMux
    port map (
            O => \N__18294\,
            I => \N__18218\
        );

    \I__3549\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18218\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__18284\,
            I => \N__18215\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__18283\,
            I => \N__18210\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__18282\,
            I => \N__18205\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__18281\,
            I => \N__18202\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__18280\,
            I => \N__18198\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__18279\,
            I => \N__18195\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__18276\,
            I => \N__18189\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__18273\,
            I => \N__18182\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__18268\,
            I => \N__18182\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__18263\,
            I => \N__18182\
        );

    \I__3538\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18179\
        );

    \I__3537\ : InMux
    port map (
            O => \N__18259\,
            I => \N__18164\
        );

    \I__3536\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18164\
        );

    \I__3535\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18164\
        );

    \I__3534\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18164\
        );

    \I__3533\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18164\
        );

    \I__3532\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18164\
        );

    \I__3531\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18164\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__18244\,
            I => \N__18157\
        );

    \I__3529\ : Span4Mux_h
    port map (
            O => \N__18241\,
            I => \N__18157\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__18232\,
            I => \N__18157\
        );

    \I__3527\ : Span12Mux_s10_h
    port map (
            O => \N__18229\,
            I => \N__18154\
        );

    \I__3526\ : Span4Mux_v
    port map (
            O => \N__18226\,
            I => \N__18151\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__18223\,
            I => \N__18144\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__18218\,
            I => \N__18144\
        );

    \I__3523\ : Span4Mux_v
    port map (
            O => \N__18215\,
            I => \N__18144\
        );

    \I__3522\ : InMux
    port map (
            O => \N__18214\,
            I => \N__18141\
        );

    \I__3521\ : InMux
    port map (
            O => \N__18213\,
            I => \N__18128\
        );

    \I__3520\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18128\
        );

    \I__3519\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18128\
        );

    \I__3518\ : InMux
    port map (
            O => \N__18208\,
            I => \N__18128\
        );

    \I__3517\ : InMux
    port map (
            O => \N__18205\,
            I => \N__18128\
        );

    \I__3516\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18128\
        );

    \I__3515\ : InMux
    port map (
            O => \N__18201\,
            I => \N__18115\
        );

    \I__3514\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18115\
        );

    \I__3513\ : InMux
    port map (
            O => \N__18195\,
            I => \N__18115\
        );

    \I__3512\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18115\
        );

    \I__3511\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18115\
        );

    \I__3510\ : InMux
    port map (
            O => \N__18192\,
            I => \N__18115\
        );

    \I__3509\ : Span4Mux_v
    port map (
            O => \N__18189\,
            I => \N__18110\
        );

    \I__3508\ : Span4Mux_s2_v
    port map (
            O => \N__18182\,
            I => \N__18110\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__18179\,
            I => \N__18103\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__18164\,
            I => \N__18103\
        );

    \I__3505\ : Span4Mux_v
    port map (
            O => \N__18157\,
            I => \N__18103\
        );

    \I__3504\ : Odrv12
    port map (
            O => \N__18154\,
            I => \tok.T_1\
        );

    \I__3503\ : Odrv4
    port map (
            O => \N__18151\,
            I => \tok.T_1\
        );

    \I__3502\ : Odrv4
    port map (
            O => \N__18144\,
            I => \tok.T_1\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__18141\,
            I => \tok.T_1\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__18128\,
            I => \tok.T_1\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__18115\,
            I => \tok.T_1\
        );

    \I__3498\ : Odrv4
    port map (
            O => \N__18110\,
            I => \tok.T_1\
        );

    \I__3497\ : Odrv4
    port map (
            O => \N__18103\,
            I => \tok.T_1\
        );

    \I__3496\ : InMux
    port map (
            O => \N__18086\,
            I => \tok.n4761\
        );

    \I__3495\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__18080\,
            I => \tok.n15_adj_664\
        );

    \I__3493\ : InMux
    port map (
            O => \N__18077\,
            I => \tok.n4762\
        );

    \I__3492\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18069\
        );

    \I__3491\ : InMux
    port map (
            O => \N__18073\,
            I => \N__18064\
        );

    \I__3490\ : InMux
    port map (
            O => \N__18072\,
            I => \N__18064\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__18069\,
            I => \tok.n82\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__18064\,
            I => \tok.n82\
        );

    \I__3487\ : InMux
    port map (
            O => \N__18059\,
            I => \N__18055\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__18058\,
            I => \N__18048\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__18055\,
            I => \N__18043\
        );

    \I__3484\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18038\
        );

    \I__3483\ : InMux
    port map (
            O => \N__18053\,
            I => \N__18038\
        );

    \I__3482\ : InMux
    port map (
            O => \N__18052\,
            I => \N__18035\
        );

    \I__3481\ : InMux
    port map (
            O => \N__18051\,
            I => \N__18031\
        );

    \I__3480\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18028\
        );

    \I__3479\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18013\
        );

    \I__3478\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18010\
        );

    \I__3477\ : Span4Mux_s3_v
    port map (
            O => \N__18043\,
            I => \N__18003\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__18038\,
            I => \N__18003\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__18035\,
            I => \N__18003\
        );

    \I__3474\ : InMux
    port map (
            O => \N__18034\,
            I => \N__17999\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__18031\,
            I => \N__17991\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__18028\,
            I => \N__17991\
        );

    \I__3471\ : InMux
    port map (
            O => \N__18027\,
            I => \N__17986\
        );

    \I__3470\ : InMux
    port map (
            O => \N__18026\,
            I => \N__17986\
        );

    \I__3469\ : InMux
    port map (
            O => \N__18025\,
            I => \N__17983\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__18024\,
            I => \N__17979\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__18023\,
            I => \N__17976\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__18022\,
            I => \N__17971\
        );

    \I__3465\ : InMux
    port map (
            O => \N__18021\,
            I => \N__17968\
        );

    \I__3464\ : InMux
    port map (
            O => \N__18020\,
            I => \N__17951\
        );

    \I__3463\ : InMux
    port map (
            O => \N__18019\,
            I => \N__17951\
        );

    \I__3462\ : InMux
    port map (
            O => \N__18018\,
            I => \N__17951\
        );

    \I__3461\ : InMux
    port map (
            O => \N__18017\,
            I => \N__17951\
        );

    \I__3460\ : InMux
    port map (
            O => \N__18016\,
            I => \N__17951\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__18013\,
            I => \N__17944\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__18010\,
            I => \N__17944\
        );

    \I__3457\ : Span4Mux_h
    port map (
            O => \N__18003\,
            I => \N__17944\
        );

    \I__3456\ : InMux
    port map (
            O => \N__18002\,
            I => \N__17941\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__17999\,
            I => \N__17938\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__17998\,
            I => \N__17935\
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__17997\,
            I => \N__17930\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__17996\,
            I => \N__17927\
        );

    \I__3451\ : Span4Mux_v
    port map (
            O => \N__17991\,
            I => \N__17921\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__17986\,
            I => \N__17921\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__17983\,
            I => \N__17918\
        );

    \I__3448\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17905\
        );

    \I__3447\ : InMux
    port map (
            O => \N__17979\,
            I => \N__17905\
        );

    \I__3446\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17905\
        );

    \I__3445\ : InMux
    port map (
            O => \N__17975\,
            I => \N__17905\
        );

    \I__3444\ : InMux
    port map (
            O => \N__17974\,
            I => \N__17905\
        );

    \I__3443\ : InMux
    port map (
            O => \N__17971\,
            I => \N__17905\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__17968\,
            I => \N__17902\
        );

    \I__3441\ : InMux
    port map (
            O => \N__17967\,
            I => \N__17889\
        );

    \I__3440\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17889\
        );

    \I__3439\ : InMux
    port map (
            O => \N__17965\,
            I => \N__17889\
        );

    \I__3438\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17889\
        );

    \I__3437\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17889\
        );

    \I__3436\ : InMux
    port map (
            O => \N__17962\,
            I => \N__17889\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__17951\,
            I => \N__17886\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__17944\,
            I => \N__17881\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__17941\,
            I => \N__17881\
        );

    \I__3432\ : Span12Mux_s10_h
    port map (
            O => \N__17938\,
            I => \N__17878\
        );

    \I__3431\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17869\
        );

    \I__3430\ : InMux
    port map (
            O => \N__17934\,
            I => \N__17869\
        );

    \I__3429\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17869\
        );

    \I__3428\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17869\
        );

    \I__3427\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17864\
        );

    \I__3426\ : InMux
    port map (
            O => \N__17926\,
            I => \N__17864\
        );

    \I__3425\ : Span4Mux_v
    port map (
            O => \N__17921\,
            I => \N__17857\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__17918\,
            I => \N__17857\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__17905\,
            I => \N__17857\
        );

    \I__3422\ : Span4Mux_h
    port map (
            O => \N__17902\,
            I => \N__17848\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__17889\,
            I => \N__17848\
        );

    \I__3420\ : Span4Mux_v
    port map (
            O => \N__17886\,
            I => \N__17848\
        );

    \I__3419\ : Span4Mux_v
    port map (
            O => \N__17881\,
            I => \N__17848\
        );

    \I__3418\ : Odrv12
    port map (
            O => \N__17878\,
            I => \tok.T_3\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__17869\,
            I => \tok.T_3\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__17864\,
            I => \tok.T_3\
        );

    \I__3415\ : Odrv4
    port map (
            O => \N__17857\,
            I => \tok.T_3\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__17848\,
            I => \tok.T_3\
        );

    \I__3413\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__17831\,
            I => \tok.n11_adj_830\
        );

    \I__3410\ : InMux
    port map (
            O => \N__17828\,
            I => \tok.n4763\
        );

    \I__3409\ : InMux
    port map (
            O => \N__17825\,
            I => \N__17822\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17819\
        );

    \I__3407\ : Odrv12
    port map (
            O => \N__17819\,
            I => \tok.n212\
        );

    \I__3406\ : InMux
    port map (
            O => \N__17816\,
            I => \tok.n4764\
        );

    \I__3405\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17809\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__17812\,
            I => \N__17804\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__17809\,
            I => \N__17801\
        );

    \I__3402\ : InMux
    port map (
            O => \N__17808\,
            I => \N__17794\
        );

    \I__3401\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17794\
        );

    \I__3400\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17794\
        );

    \I__3399\ : Span4Mux_v
    port map (
            O => \N__17801\,
            I => \N__17791\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__17794\,
            I => \N__17788\
        );

    \I__3397\ : Span4Mux_h
    port map (
            O => \N__17791\,
            I => \N__17785\
        );

    \I__3396\ : Span4Mux_h
    port map (
            O => \N__17788\,
            I => \N__17782\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__17785\,
            I => \N__17779\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__17782\,
            I => \tok.uart_tx_busy\
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__17779\,
            I => \tok.uart_tx_busy\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__17774\,
            I => \tok.n15_adj_655_cascade_\
        );

    \I__3391\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17759\
        );

    \I__3390\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17759\
        );

    \I__3389\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17759\
        );

    \I__3388\ : InMux
    port map (
            O => \N__17768\,
            I => \N__17759\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__17759\,
            I => \N__17756\
        );

    \I__3386\ : Sp12to4
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__3385\ : Odrv12
    port map (
            O => \N__17753\,
            I => \tok.uart_stall\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__17750\,
            I => \N__17746\
        );

    \I__3383\ : InMux
    port map (
            O => \N__17749\,
            I => \N__17742\
        );

    \I__3382\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17737\
        );

    \I__3381\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17737\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__17742\,
            I => \tok.uart_rx_valid\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__17737\,
            I => \tok.uart_rx_valid\
        );

    \I__3378\ : CEMux
    port map (
            O => \N__17732\,
            I => \N__17729\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__17729\,
            I => \N__17726\
        );

    \I__3376\ : Odrv4
    port map (
            O => \N__17726\,
            I => \tok.uart.n953\
        );

    \I__3375\ : CascadeMux
    port map (
            O => \N__17723\,
            I => \tok.n15_adj_667_cascade_\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__17720\,
            I => \N__17716\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__17719\,
            I => \N__17713\
        );

    \I__3372\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17710\
        );

    \I__3371\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17707\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__17710\,
            I => \N__17704\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__17707\,
            I => \N__17701\
        );

    \I__3368\ : Span4Mux_h
    port map (
            O => \N__17704\,
            I => \N__17698\
        );

    \I__3367\ : Span4Mux_s3_h
    port map (
            O => \N__17701\,
            I => \N__17695\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__17698\,
            I => \tok.table_rd_2\
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__17695\,
            I => \tok.table_rd_2\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__17690\,
            I => \tok.n28_adj_771_cascade_\
        );

    \I__3363\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__17684\,
            I => \tok.n5470\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__17681\,
            I => \tok.n5467_cascade_\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__17678\,
            I => \N__17674\
        );

    \I__3359\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17669\
        );

    \I__3358\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17669\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__17669\,
            I => \N__17666\
        );

    \I__3356\ : Odrv12
    port map (
            O => \N__17666\,
            I => \tok.n34\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__17663\,
            I => \N__17660\
        );

    \I__3354\ : InMux
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__17657\,
            I => \tok.n5462\
        );

    \I__3352\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17651\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__17651\,
            I => \tok.n5566\
        );

    \I__3350\ : InMux
    port map (
            O => \N__17648\,
            I => \N__17645\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__17645\,
            I => \N__17642\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__17642\,
            I => \tok.n5561\
        );

    \I__3347\ : InMux
    port map (
            O => \N__17639\,
            I => \N__17635\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__17638\,
            I => \N__17632\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__17635\,
            I => \N__17629\
        );

    \I__3344\ : InMux
    port map (
            O => \N__17632\,
            I => \N__17626\
        );

    \I__3343\ : Span4Mux_v
    port map (
            O => \N__17629\,
            I => \N__17621\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__17626\,
            I => \N__17621\
        );

    \I__3341\ : Span4Mux_v
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__17618\,
            I => \tok.n9_adj_766\
        );

    \I__3339\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17607\
        );

    \I__3338\ : InMux
    port map (
            O => \N__17614\,
            I => \N__17602\
        );

    \I__3337\ : InMux
    port map (
            O => \N__17613\,
            I => \N__17602\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__17612\,
            I => \N__17599\
        );

    \I__3335\ : InMux
    port map (
            O => \N__17611\,
            I => \N__17593\
        );

    \I__3334\ : InMux
    port map (
            O => \N__17610\,
            I => \N__17593\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__17607\,
            I => \N__17590\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__17602\,
            I => \N__17587\
        );

    \I__3331\ : InMux
    port map (
            O => \N__17599\,
            I => \N__17582\
        );

    \I__3330\ : InMux
    port map (
            O => \N__17598\,
            I => \N__17582\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__17593\,
            I => \N__17579\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__17590\,
            I => \tok.n10_adj_643\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__17587\,
            I => \tok.n10_adj_643\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__17582\,
            I => \tok.n10_adj_643\
        );

    \I__3325\ : Odrv4
    port map (
            O => \N__17579\,
            I => \tok.n10_adj_643\
        );

    \I__3324\ : CascadeMux
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__3323\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__3321\ : Span4Mux_h
    port map (
            O => \N__17561\,
            I => \N__17557\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__17560\,
            I => \N__17554\
        );

    \I__3319\ : Span4Mux_h
    port map (
            O => \N__17557\,
            I => \N__17551\
        );

    \I__3318\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17548\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__17551\,
            I => \tok.table_rd_0\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__17548\,
            I => \tok.table_rd_0\
        );

    \I__3315\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17540\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__3313\ : Odrv12
    port map (
            O => \N__17537\,
            I => \tok.n31\
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__17534\,
            I => \tok.n5463_cascade_\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__17531\,
            I => \N__17525\
        );

    \I__3310\ : InMux
    port map (
            O => \N__17530\,
            I => \N__17522\
        );

    \I__3309\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17517\
        );

    \I__3308\ : InMux
    port map (
            O => \N__17528\,
            I => \N__17517\
        );

    \I__3307\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17514\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__17522\,
            I => \N__17509\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__17517\,
            I => \N__17509\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__17514\,
            I => \N__17506\
        );

    \I__3303\ : Span4Mux_h
    port map (
            O => \N__17509\,
            I => \N__17503\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__17506\,
            I => \tok.n2607\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__17503\,
            I => \tok.n2607\
        );

    \I__3300\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17495\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__17495\,
            I => \N__17492\
        );

    \I__3298\ : Span4Mux_s2_h
    port map (
            O => \N__17492\,
            I => \N__17488\
        );

    \I__3297\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17484\
        );

    \I__3296\ : Span4Mux_h
    port map (
            O => \N__17488\,
            I => \N__17479\
        );

    \I__3295\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17476\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__17484\,
            I => \N__17473\
        );

    \I__3293\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17468\
        );

    \I__3292\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17468\
        );

    \I__3291\ : Odrv4
    port map (
            O => \N__17479\,
            I => \tok.n14_adj_765\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__17476\,
            I => \tok.n14_adj_765\
        );

    \I__3289\ : Odrv4
    port map (
            O => \N__17473\,
            I => \tok.n14_adj_765\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__17468\,
            I => \tok.n14_adj_765\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__17459\,
            I => \N__17455\
        );

    \I__3286\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17452\
        );

    \I__3285\ : InMux
    port map (
            O => \N__17455\,
            I => \N__17449\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__17452\,
            I => \N__17446\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__17449\,
            I => \N__17443\
        );

    \I__3282\ : Span4Mux_v
    port map (
            O => \N__17446\,
            I => \N__17440\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__17443\,
            I => \N__17437\
        );

    \I__3280\ : Span4Mux_h
    port map (
            O => \N__17440\,
            I => \N__17434\
        );

    \I__3279\ : Span4Mux_v
    port map (
            O => \N__17437\,
            I => \N__17431\
        );

    \I__3278\ : Odrv4
    port map (
            O => \N__17434\,
            I => \tok.table_rd_1\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__17431\,
            I => \tok.table_rd_1\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__17426\,
            I => \tok.n5334_cascade_\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__17423\,
            I => \tok.n14_adj_735_cascade_\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__17420\,
            I => \N__17417\
        );

    \I__3273\ : InMux
    port map (
            O => \N__17417\,
            I => \N__17411\
        );

    \I__3272\ : InMux
    port map (
            O => \N__17416\,
            I => \N__17411\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__3270\ : Span4Mux_h
    port map (
            O => \N__17408\,
            I => \N__17405\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__17405\,
            I => \tok.n6_adj_754\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__17402\,
            I => \N__17398\
        );

    \I__3267\ : InMux
    port map (
            O => \N__17401\,
            I => \N__17395\
        );

    \I__3266\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17392\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__17395\,
            I => \N__17389\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__17392\,
            I => \N__17386\
        );

    \I__3263\ : Span4Mux_v
    port map (
            O => \N__17389\,
            I => \N__17383\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__17386\,
            I => \N__17380\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__17383\,
            I => \tok.table_rd_4\
        );

    \I__3260\ : Odrv4
    port map (
            O => \N__17380\,
            I => \tok.table_rd_4\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__17375\,
            I => \tok.n16_adj_851_cascade_\
        );

    \I__3258\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17369\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__17369\,
            I => \N__17366\
        );

    \I__3256\ : Span4Mux_h
    port map (
            O => \N__17366\,
            I => \N__17363\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__17363\,
            I => \tok.n17_adj_853\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__17360\,
            I => \tok.n5562_cascade_\
        );

    \I__3253\ : InMux
    port map (
            O => \N__17357\,
            I => \N__17354\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__17354\,
            I => \tok.n13_adj_852\
        );

    \I__3251\ : InMux
    port map (
            O => \N__17351\,
            I => \N__17348\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__17348\,
            I => \tok.n14_adj_854\
        );

    \I__3249\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17340\
        );

    \I__3248\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17335\
        );

    \I__3247\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17335\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__17340\,
            I => capture_3
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__17335\,
            I => capture_3
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__17330\,
            I => \N__17327\
        );

    \I__3243\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__17324\,
            I => \N__17321\
        );

    \I__3241\ : Span4Mux_h
    port map (
            O => \N__17321\,
            I => \N__17317\
        );

    \I__3240\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17314\
        );

    \I__3239\ : Sp12to4
    port map (
            O => \N__17317\,
            I => \N__17311\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__17314\,
            I => capture_0
        );

    \I__3237\ : Odrv12
    port map (
            O => \N__17311\,
            I => capture_0
        );

    \I__3236\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17297\
        );

    \I__3235\ : InMux
    port map (
            O => \N__17305\,
            I => \N__17297\
        );

    \I__3234\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17297\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__17297\,
            I => capture_1
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__17294\,
            I => \N__17290\
        );

    \I__3231\ : InMux
    port map (
            O => \N__17293\,
            I => \N__17285\
        );

    \I__3230\ : InMux
    port map (
            O => \N__17290\,
            I => \N__17285\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__17285\,
            I => uart_rx_data_0
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__17282\,
            I => \tok.n6_adj_794_cascade_\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__17279\,
            I => \N__17276\
        );

    \I__3226\ : InMux
    port map (
            O => \N__17276\,
            I => \N__17272\
        );

    \I__3225\ : InMux
    port map (
            O => \N__17275\,
            I => \N__17269\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__17272\,
            I => \N__17266\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__17269\,
            I => \N__17263\
        );

    \I__3222\ : Span4Mux_v
    port map (
            O => \N__17266\,
            I => \N__17260\
        );

    \I__3221\ : Span4Mux_v
    port map (
            O => \N__17263\,
            I => \N__17257\
        );

    \I__3220\ : Span4Mux_v
    port map (
            O => \N__17260\,
            I => \N__17254\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__17257\,
            I => \tok.table_rd_6\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__17254\,
            I => \tok.table_rd_6\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__17249\,
            I => \tok.n5553_cascade_\
        );

    \I__3216\ : InMux
    port map (
            O => \N__17246\,
            I => \N__17243\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__17243\,
            I => \N__17240\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__17240\,
            I => \N__17237\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__17237\,
            I => \tok.table_rd_14\
        );

    \I__3212\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17231\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__17231\,
            I => \N__17228\
        );

    \I__3210\ : Span4Mux_v
    port map (
            O => \N__17228\,
            I => \N__17225\
        );

    \I__3209\ : Span4Mux_h
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__17222\,
            I => \tok.table_rd_12\
        );

    \I__3207\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17216\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__17216\,
            I => \N__17212\
        );

    \I__3205\ : InMux
    port map (
            O => \N__17215\,
            I => \N__17209\
        );

    \I__3204\ : Span4Mux_v
    port map (
            O => \N__17212\,
            I => \N__17206\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__17209\,
            I => tail_110
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__17206\,
            I => tail_110
        );

    \I__3201\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__17198\,
            I => \N__17194\
        );

    \I__3199\ : InMux
    port map (
            O => \N__17197\,
            I => \N__17191\
        );

    \I__3198\ : Odrv12
    port map (
            O => \N__17194\,
            I => tail_126
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__17191\,
            I => tail_126
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__17186\,
            I => \N__17183\
        );

    \I__3195\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17180\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__17180\,
            I => \N__17177\
        );

    \I__3193\ : Span4Mux_v
    port map (
            O => \N__17177\,
            I => \N__17173\
        );

    \I__3192\ : InMux
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__3191\ : Sp12to4
    port map (
            O => \N__17173\,
            I => \N__17167\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__17170\,
            I => \N__17164\
        );

    \I__3189\ : Odrv12
    port map (
            O => \N__17167\,
            I => tail_111
        );

    \I__3188\ : Odrv12
    port map (
            O => \N__17164\,
            I => tail_111
        );

    \I__3187\ : InMux
    port map (
            O => \N__17159\,
            I => \N__17155\
        );

    \I__3186\ : InMux
    port map (
            O => \N__17158\,
            I => \N__17152\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__17155\,
            I => \N__17148\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__17152\,
            I => \N__17145\
        );

    \I__3183\ : InMux
    port map (
            O => \N__17151\,
            I => \N__17142\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__17148\,
            I => \N__17137\
        );

    \I__3181\ : Span4Mux_h
    port map (
            O => \N__17145\,
            I => \N__17137\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__17142\,
            I => \N__17134\
        );

    \I__3179\ : Sp12to4
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__17134\,
            I => \N__17128\
        );

    \I__3177\ : Odrv12
    port map (
            O => \N__17131\,
            I => rx_c
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__17128\,
            I => rx_c
        );

    \I__3175\ : InMux
    port map (
            O => \N__17123\,
            I => \N__17120\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__3173\ : Span4Mux_h
    port map (
            O => \N__17117\,
            I => \N__17114\
        );

    \I__3172\ : Odrv4
    port map (
            O => \N__17114\,
            I => \tok.uart.n5235\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__3170\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17102\
        );

    \I__3169\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17102\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__17102\,
            I => \N__17098\
        );

    \I__3167\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17094\
        );

    \I__3166\ : Span4Mux_h
    port map (
            O => \N__17098\,
            I => \N__17091\
        );

    \I__3165\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17088\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__17094\,
            I => \N__17083\
        );

    \I__3163\ : Span4Mux_h
    port map (
            O => \N__17091\,
            I => \N__17083\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__17088\,
            I => \tok.uart.bytephase_5\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__17083\,
            I => \tok.uart.bytephase_5\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__17078\,
            I => \N__17073\
        );

    \I__3159\ : InMux
    port map (
            O => \N__17077\,
            I => \N__17068\
        );

    \I__3158\ : InMux
    port map (
            O => \N__17076\,
            I => \N__17068\
        );

    \I__3157\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17064\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__17068\,
            I => \N__17061\
        );

    \I__3155\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17058\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__17064\,
            I => \N__17053\
        );

    \I__3153\ : Span12Mux_s11_h
    port map (
            O => \N__17061\,
            I => \N__17053\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__17058\,
            I => \tok.uart.bytephase_3\
        );

    \I__3151\ : Odrv12
    port map (
            O => \N__17053\,
            I => \tok.uart.bytephase_3\
        );

    \I__3150\ : InMux
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__3148\ : Span4Mux_v
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__3147\ : Odrv4
    port map (
            O => \N__17039\,
            I => \tok.uart.n5374\
        );

    \I__3146\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17032\
        );

    \I__3145\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17029\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__17032\,
            I => \N__17024\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__17029\,
            I => \N__17024\
        );

    \I__3142\ : Span4Mux_h
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__17021\,
            I => \tok.key_rd_13\
        );

    \I__3140\ : InMux
    port map (
            O => \N__17018\,
            I => \N__17015\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__17012\,
            I => \tok.n14_adj_647\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__17009\,
            I => \tok.n27_adj_818_cascade_\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__17006\,
            I => \N__17002\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__17005\,
            I => \N__16999\
        );

    \I__3134\ : CascadeBuf
    port map (
            O => \N__17002\,
            I => \N__16996\
        );

    \I__3133\ : CascadeBuf
    port map (
            O => \N__16999\,
            I => \N__16993\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__16996\,
            I => \N__16990\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__16993\,
            I => \N__16987\
        );

    \I__3130\ : InMux
    port map (
            O => \N__16990\,
            I => \N__16984\
        );

    \I__3129\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16981\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__16984\,
            I => \N__16976\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__16981\,
            I => \N__16976\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__16976\,
            I => \N__16970\
        );

    \I__3125\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16967\
        );

    \I__3124\ : InMux
    port map (
            O => \N__16974\,
            I => \N__16964\
        );

    \I__3123\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16961\
        );

    \I__3122\ : Span4Mux_h
    port map (
            O => \N__16970\,
            I => \N__16958\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__16967\,
            I => \tok.idx_2\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__16964\,
            I => \tok.idx_2\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__16961\,
            I => \tok.idx_2\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__16958\,
            I => \tok.idx_2\
        );

    \I__3117\ : InMux
    port map (
            O => \N__16949\,
            I => \N__16945\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__16948\,
            I => \N__16936\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__16945\,
            I => \N__16927\
        );

    \I__3114\ : InMux
    port map (
            O => \N__16944\,
            I => \N__16924\
        );

    \I__3113\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16917\
        );

    \I__3112\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16917\
        );

    \I__3111\ : InMux
    port map (
            O => \N__16941\,
            I => \N__16912\
        );

    \I__3110\ : InMux
    port map (
            O => \N__16940\,
            I => \N__16912\
        );

    \I__3109\ : InMux
    port map (
            O => \N__16939\,
            I => \N__16909\
        );

    \I__3108\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16902\
        );

    \I__3107\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16902\
        );

    \I__3106\ : InMux
    port map (
            O => \N__16934\,
            I => \N__16902\
        );

    \I__3105\ : InMux
    port map (
            O => \N__16933\,
            I => \N__16893\
        );

    \I__3104\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16893\
        );

    \I__3103\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16893\
        );

    \I__3102\ : InMux
    port map (
            O => \N__16930\,
            I => \N__16893\
        );

    \I__3101\ : Span4Mux_v
    port map (
            O => \N__16927\,
            I => \N__16890\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__16924\,
            I => \N__16887\
        );

    \I__3099\ : InMux
    port map (
            O => \N__16923\,
            I => \N__16882\
        );

    \I__3098\ : InMux
    port map (
            O => \N__16922\,
            I => \N__16882\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__16917\,
            I => \tok.stall\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__16912\,
            I => \tok.stall\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__16909\,
            I => \tok.stall\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__16902\,
            I => \tok.stall\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__16893\,
            I => \tok.stall\
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__16890\,
            I => \tok.stall\
        );

    \I__3091\ : Odrv12
    port map (
            O => \N__16887\,
            I => \tok.stall\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__16882\,
            I => \tok.stall\
        );

    \I__3089\ : InMux
    port map (
            O => \N__16865\,
            I => \N__16862\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__16862\,
            I => \tok.n33_adj_821\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__16859\,
            I => \N__16850\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__16858\,
            I => \N__16845\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__16857\,
            I => \N__16841\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__16856\,
            I => \N__16838\
        );

    \I__3083\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16828\
        );

    \I__3082\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16828\
        );

    \I__3081\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16828\
        );

    \I__3080\ : InMux
    port map (
            O => \N__16850\,
            I => \N__16828\
        );

    \I__3079\ : InMux
    port map (
            O => \N__16849\,
            I => \N__16821\
        );

    \I__3078\ : InMux
    port map (
            O => \N__16848\,
            I => \N__16821\
        );

    \I__3077\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16821\
        );

    \I__3076\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16812\
        );

    \I__3075\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16812\
        );

    \I__3074\ : InMux
    port map (
            O => \N__16838\,
            I => \N__16812\
        );

    \I__3073\ : InMux
    port map (
            O => \N__16837\,
            I => \N__16812\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__16828\,
            I => \tok.search_clk\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__16821\,
            I => \tok.search_clk\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__16812\,
            I => \tok.search_clk\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__16805\,
            I => \tok.n27_adj_822_cascade_\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__16802\,
            I => \N__16799\
        );

    \I__3067\ : CascadeBuf
    port map (
            O => \N__16799\,
            I => \N__16795\
        );

    \I__3066\ : CascadeMux
    port map (
            O => \N__16798\,
            I => \N__16792\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__16795\,
            I => \N__16789\
        );

    \I__3064\ : CascadeBuf
    port map (
            O => \N__16792\,
            I => \N__16786\
        );

    \I__3063\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16783\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__16786\,
            I => \N__16780\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__16783\,
            I => \N__16777\
        );

    \I__3060\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16774\
        );

    \I__3059\ : Span4Mux_h
    port map (
            O => \N__16777\,
            I => \N__16771\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__16774\,
            I => \N__16765\
        );

    \I__3057\ : Span4Mux_h
    port map (
            O => \N__16771\,
            I => \N__16762\
        );

    \I__3056\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16759\
        );

    \I__3055\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16756\
        );

    \I__3054\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16753\
        );

    \I__3053\ : Span12Mux_s7_h
    port map (
            O => \N__16765\,
            I => \N__16750\
        );

    \I__3052\ : Span4Mux_v
    port map (
            O => \N__16762\,
            I => \N__16747\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__16759\,
            I => \tok.idx_3\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__16756\,
            I => \tok.idx_3\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__16753\,
            I => \tok.idx_3\
        );

    \I__3048\ : Odrv12
    port map (
            O => \N__16750\,
            I => \tok.idx_3\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__16747\,
            I => \tok.idx_3\
        );

    \I__3046\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16720\
        );

    \I__3045\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16720\
        );

    \I__3044\ : InMux
    port map (
            O => \N__16734\,
            I => \N__16720\
        );

    \I__3043\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16720\
        );

    \I__3042\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16713\
        );

    \I__3041\ : InMux
    port map (
            O => \N__16731\,
            I => \N__16713\
        );

    \I__3040\ : InMux
    port map (
            O => \N__16730\,
            I => \N__16713\
        );

    \I__3039\ : InMux
    port map (
            O => \N__16729\,
            I => \N__16710\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__16720\,
            I => \tok.n2699\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__16713\,
            I => \tok.n2699\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__16710\,
            I => \tok.n2699\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__16703\,
            I => \N__16694\
        );

    \I__3034\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16684\
        );

    \I__3033\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16684\
        );

    \I__3032\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16684\
        );

    \I__3031\ : InMux
    port map (
            O => \N__16699\,
            I => \N__16684\
        );

    \I__3030\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16677\
        );

    \I__3029\ : InMux
    port map (
            O => \N__16697\,
            I => \N__16677\
        );

    \I__3028\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16677\
        );

    \I__3027\ : InMux
    port map (
            O => \N__16693\,
            I => \N__16674\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__16684\,
            I => \tok.n5282\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__16677\,
            I => \tok.n5282\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__16674\,
            I => \tok.n5282\
        );

    \I__3023\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__16664\,
            I => \tok.n27_adj_815\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__3020\ : CascadeBuf
    port map (
            O => \N__16658\,
            I => \N__16654\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__16657\,
            I => \N__16651\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__16654\,
            I => \N__16648\
        );

    \I__3017\ : CascadeBuf
    port map (
            O => \N__16651\,
            I => \N__16645\
        );

    \I__3016\ : InMux
    port map (
            O => \N__16648\,
            I => \N__16642\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__16645\,
            I => \N__16639\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__16642\,
            I => \N__16636\
        );

    \I__3013\ : InMux
    port map (
            O => \N__16639\,
            I => \N__16633\
        );

    \I__3012\ : Span4Mux_h
    port map (
            O => \N__16636\,
            I => \N__16627\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__16633\,
            I => \N__16624\
        );

    \I__3010\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16621\
        );

    \I__3009\ : InMux
    port map (
            O => \N__16631\,
            I => \N__16618\
        );

    \I__3008\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16615\
        );

    \I__3007\ : Sp12to4
    port map (
            O => \N__16627\,
            I => \N__16610\
        );

    \I__3006\ : Span12Mux_s7_h
    port map (
            O => \N__16624\,
            I => \N__16610\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__16621\,
            I => \tok.idx_1\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__16618\,
            I => \tok.idx_1\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__16615\,
            I => \tok.idx_1\
        );

    \I__3002\ : Odrv12
    port map (
            O => \N__16610\,
            I => \tok.idx_1\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__16601\,
            I => \rd_15__N_301_cascade_\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__2999\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16589\
        );

    \I__2998\ : InMux
    port map (
            O => \N__16594\,
            I => \N__16589\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__16589\,
            I => \tok.n797\
        );

    \I__2996\ : InMux
    port map (
            O => \N__16586\,
            I => \N__16579\
        );

    \I__2995\ : InMux
    port map (
            O => \N__16585\,
            I => \N__16579\
        );

    \I__2994\ : InMux
    port map (
            O => \N__16584\,
            I => \N__16576\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__16579\,
            I => \N__16573\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__16576\,
            I => \N__16570\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__16573\,
            I => \tok.n2585\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__16570\,
            I => \tok.n2585\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__16565\,
            I => \A_stk_delta_1_cascade_\
        );

    \I__2988\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16556\
        );

    \I__2987\ : InMux
    port map (
            O => \N__16561\,
            I => \N__16556\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__16556\,
            I => \tok.A_stk.tail_78\
        );

    \I__2985\ : InMux
    port map (
            O => \N__16553\,
            I => \N__16547\
        );

    \I__2984\ : InMux
    port map (
            O => \N__16552\,
            I => \N__16547\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__16547\,
            I => \tok.A_stk.tail_62\
        );

    \I__2982\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16538\
        );

    \I__2981\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16538\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__16538\,
            I => \tok.A_stk.tail_46\
        );

    \I__2979\ : InMux
    port map (
            O => \N__16535\,
            I => \N__16529\
        );

    \I__2978\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16529\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__16529\,
            I => \tok.A_stk.tail_30\
        );

    \I__2976\ : InMux
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__2974\ : Span4Mux_s2_v
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__2973\ : Span4Mux_h
    port map (
            O => \N__16517\,
            I => \N__16513\
        );

    \I__2972\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16510\
        );

    \I__2971\ : Odrv4
    port map (
            O => \N__16513\,
            I => tail_127
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__16510\,
            I => tail_127
        );

    \I__2969\ : InMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__16502\,
            I => \tok.n33_adj_814\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__16499\,
            I => \N__16494\
        );

    \I__2966\ : InMux
    port map (
            O => \N__16498\,
            I => \N__16489\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__16497\,
            I => \N__16485\
        );

    \I__2964\ : InMux
    port map (
            O => \N__16494\,
            I => \N__16481\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__16493\,
            I => \N__16477\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__16492\,
            I => \N__16473\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__16489\,
            I => \N__16470\
        );

    \I__2960\ : InMux
    port map (
            O => \N__16488\,
            I => \N__16463\
        );

    \I__2959\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16463\
        );

    \I__2958\ : InMux
    port map (
            O => \N__16484\,
            I => \N__16463\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__16481\,
            I => \N__16460\
        );

    \I__2956\ : InMux
    port map (
            O => \N__16480\,
            I => \N__16451\
        );

    \I__2955\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16451\
        );

    \I__2954\ : InMux
    port map (
            O => \N__16476\,
            I => \N__16451\
        );

    \I__2953\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16451\
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__16470\,
            I => \tok.n62\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__16463\,
            I => \tok.n62\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__16460\,
            I => \tok.n62\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__16451\,
            I => \tok.n62\
        );

    \I__2948\ : InMux
    port map (
            O => \N__16442\,
            I => \N__16439\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__16439\,
            I => \N__16436\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__16436\,
            I => \N__16429\
        );

    \I__2945\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16422\
        );

    \I__2944\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16422\
        );

    \I__2943\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16422\
        );

    \I__2942\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16419\
        );

    \I__2941\ : Odrv4
    port map (
            O => \N__16429\,
            I => \tok.n1_adj_715\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__16422\,
            I => \tok.n1_adj_715\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__16419\,
            I => \tok.n1_adj_715\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__16412\,
            I => \tok.depth_0_cascade_\
        );

    \I__2937\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__2935\ : Odrv12
    port map (
            O => \N__16403\,
            I => \tok.n5408\
        );

    \I__2934\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16397\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__16397\,
            I => \tok.n33_adj_816\
        );

    \I__2932\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16391\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__16391\,
            I => \N__16387\
        );

    \I__2930\ : InMux
    port map (
            O => \N__16390\,
            I => \N__16384\
        );

    \I__2929\ : Span4Mux_h
    port map (
            O => \N__16387\,
            I => \N__16377\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__16384\,
            I => \N__16377\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__16383\,
            I => \N__16374\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__16382\,
            I => \N__16371\
        );

    \I__2925\ : Span4Mux_v
    port map (
            O => \N__16377\,
            I => \N__16366\
        );

    \I__2924\ : InMux
    port map (
            O => \N__16374\,
            I => \N__16361\
        );

    \I__2923\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16361\
        );

    \I__2922\ : InMux
    port map (
            O => \N__16370\,
            I => \N__16358\
        );

    \I__2921\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16354\
        );

    \I__2920\ : Span4Mux_s3_h
    port map (
            O => \N__16366\,
            I => \N__16348\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__16361\,
            I => \N__16348\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__16358\,
            I => \N__16345\
        );

    \I__2917\ : InMux
    port map (
            O => \N__16357\,
            I => \N__16342\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__16354\,
            I => \N__16339\
        );

    \I__2915\ : InMux
    port map (
            O => \N__16353\,
            I => \N__16336\
        );

    \I__2914\ : Span4Mux_v
    port map (
            O => \N__16348\,
            I => \N__16333\
        );

    \I__2913\ : Span4Mux_h
    port map (
            O => \N__16345\,
            I => \N__16330\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__16342\,
            I => \N__16327\
        );

    \I__2911\ : Odrv12
    port map (
            O => \N__16339\,
            I => \tok.n820\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__16336\,
            I => \tok.n820\
        );

    \I__2909\ : Odrv4
    port map (
            O => \N__16333\,
            I => \tok.n820\
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__16330\,
            I => \tok.n820\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__16327\,
            I => \tok.n820\
        );

    \I__2906\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16313\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__16313\,
            I => \N__16306\
        );

    \I__2904\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16303\
        );

    \I__2903\ : InMux
    port map (
            O => \N__16311\,
            I => \N__16298\
        );

    \I__2902\ : InMux
    port map (
            O => \N__16310\,
            I => \N__16298\
        );

    \I__2901\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16295\
        );

    \I__2900\ : Span4Mux_v
    port map (
            O => \N__16306\,
            I => \N__16290\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__16303\,
            I => \N__16285\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__16298\,
            I => \N__16285\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__16295\,
            I => \N__16282\
        );

    \I__2896\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16278\
        );

    \I__2895\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16275\
        );

    \I__2894\ : Span4Mux_v
    port map (
            O => \N__16290\,
            I => \N__16268\
        );

    \I__2893\ : Span4Mux_v
    port map (
            O => \N__16285\,
            I => \N__16268\
        );

    \I__2892\ : Span4Mux_v
    port map (
            O => \N__16282\,
            I => \N__16268\
        );

    \I__2891\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16265\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__16278\,
            I => \tok.n5298\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__16275\,
            I => \tok.n5298\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__16268\,
            I => \tok.n5298\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__16265\,
            I => \tok.n5298\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__16256\,
            I => \tok.n13_adj_673_cascade_\
        );

    \I__2885\ : InMux
    port map (
            O => \N__16253\,
            I => \N__16248\
        );

    \I__2884\ : InMux
    port map (
            O => \N__16252\,
            I => \N__16243\
        );

    \I__2883\ : InMux
    port map (
            O => \N__16251\,
            I => \N__16243\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__16248\,
            I => \N__16239\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__16243\,
            I => \N__16236\
        );

    \I__2880\ : InMux
    port map (
            O => \N__16242\,
            I => \N__16233\
        );

    \I__2879\ : Span4Mux_h
    port map (
            O => \N__16239\,
            I => \N__16228\
        );

    \I__2878\ : Span4Mux_s3_v
    port map (
            O => \N__16236\,
            I => \N__16228\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__16233\,
            I => \tok.tc_plus_1_4\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__16228\,
            I => \tok.tc_plus_1_4\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__16223\,
            I => \n10_adj_870_cascade_\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__16220\,
            I => \N__16217\
        );

    \I__2873\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16214\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__16214\,
            I => \N__16211\
        );

    \I__2871\ : Span4Mux_h
    port map (
            O => \N__16211\,
            I => \N__16208\
        );

    \I__2870\ : Odrv4
    port map (
            O => \N__16208\,
            I => \tok.tc_4\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__16205\,
            I => \N__16198\
        );

    \I__2868\ : InMux
    port map (
            O => \N__16204\,
            I => \N__16191\
        );

    \I__2867\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16186\
        );

    \I__2866\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16186\
        );

    \I__2865\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16173\
        );

    \I__2864\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16173\
        );

    \I__2863\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16173\
        );

    \I__2862\ : InMux
    port map (
            O => \N__16196\,
            I => \N__16173\
        );

    \I__2861\ : InMux
    port map (
            O => \N__16195\,
            I => \N__16173\
        );

    \I__2860\ : InMux
    port map (
            O => \N__16194\,
            I => \N__16173\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__16191\,
            I => \N__16168\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__16186\,
            I => \N__16165\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__16173\,
            I => \N__16159\
        );

    \I__2856\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16154\
        );

    \I__2855\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16154\
        );

    \I__2854\ : Span4Mux_v
    port map (
            O => \N__16168\,
            I => \N__16149\
        );

    \I__2853\ : Span4Mux_h
    port map (
            O => \N__16165\,
            I => \N__16149\
        );

    \I__2852\ : InMux
    port map (
            O => \N__16164\,
            I => \N__16144\
        );

    \I__2851\ : InMux
    port map (
            O => \N__16163\,
            I => \N__16144\
        );

    \I__2850\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16141\
        );

    \I__2849\ : Span4Mux_h
    port map (
            O => \N__16159\,
            I => \N__16136\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__16154\,
            I => \N__16136\
        );

    \I__2847\ : Sp12to4
    port map (
            O => \N__16149\,
            I => \N__16127\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__16144\,
            I => \N__16127\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__16141\,
            I => \N__16127\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__16136\,
            I => \N__16124\
        );

    \I__2843\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16119\
        );

    \I__2842\ : InMux
    port map (
            O => \N__16134\,
            I => \N__16119\
        );

    \I__2841\ : Odrv12
    port map (
            O => \N__16127\,
            I => \stall_\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__16124\,
            I => \stall_\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__16119\,
            I => \stall_\
        );

    \I__2838\ : InMux
    port map (
            O => \N__16112\,
            I => \N__16109\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__16109\,
            I => n10_adj_870
        );

    \I__2836\ : InMux
    port map (
            O => \N__16106\,
            I => \N__16101\
        );

    \I__2835\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16098\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__16104\,
            I => \N__16095\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__16101\,
            I => \N__16091\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__16098\,
            I => \N__16088\
        );

    \I__2831\ : InMux
    port map (
            O => \N__16095\,
            I => \N__16083\
        );

    \I__2830\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16083\
        );

    \I__2829\ : Span4Mux_v
    port map (
            O => \N__16091\,
            I => \N__16080\
        );

    \I__2828\ : Odrv12
    port map (
            O => \N__16088\,
            I => tc_4
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__16083\,
            I => tc_4
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__16080\,
            I => tc_4
        );

    \I__2825\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16068\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__16072\,
            I => \N__16064\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__16071\,
            I => \N__16061\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__16068\,
            I => \N__16058\
        );

    \I__2821\ : InMux
    port map (
            O => \N__16067\,
            I => \N__16053\
        );

    \I__2820\ : InMux
    port map (
            O => \N__16064\,
            I => \N__16053\
        );

    \I__2819\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16050\
        );

    \I__2818\ : Span4Mux_s2_v
    port map (
            O => \N__16058\,
            I => \N__16047\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__16053\,
            I => \N__16044\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__16050\,
            I => \tok.c_stk_r_4\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__16047\,
            I => \tok.c_stk_r_4\
        );

    \I__2814\ : Odrv12
    port map (
            O => \N__16044\,
            I => \tok.c_stk_r_4\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__16037\,
            I => \tok.n83_adj_665_cascade_\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__16034\,
            I => \N__16031\
        );

    \I__2811\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16028\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__16028\,
            I => \tok.n5487\
        );

    \I__2809\ : InMux
    port map (
            O => \N__16025\,
            I => \N__16021\
        );

    \I__2808\ : InMux
    port map (
            O => \N__16024\,
            I => \N__16018\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__16021\,
            I => \tok.A_stk.tail_94\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__16018\,
            I => \tok.A_stk.tail_94\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__16013\,
            I => \N__16010\
        );

    \I__2804\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16007\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__16007\,
            I => \tok.n5423\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__16004\,
            I => \N__16001\
        );

    \I__2801\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15998\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__15998\,
            I => \tok.n42_adj_751\
        );

    \I__2799\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15992\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__15992\,
            I => \N__15987\
        );

    \I__2797\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15984\
        );

    \I__2796\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15981\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__15987\,
            I => \N__15978\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__15984\,
            I => capture_9
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__15981\,
            I => capture_9
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__15978\,
            I => capture_9
        );

    \I__2791\ : InMux
    port map (
            O => \N__15971\,
            I => \N__15968\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__15968\,
            I => \tok.n2609\
        );

    \I__2789\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15957\
        );

    \I__2788\ : InMux
    port map (
            O => \N__15964\,
            I => \N__15954\
        );

    \I__2787\ : InMux
    port map (
            O => \N__15963\,
            I => \N__15950\
        );

    \I__2786\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15947\
        );

    \I__2785\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15943\
        );

    \I__2784\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15940\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__15957\,
            I => \N__15935\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__15954\,
            I => \N__15935\
        );

    \I__2781\ : InMux
    port map (
            O => \N__15953\,
            I => \N__15932\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__15950\,
            I => \N__15929\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__15947\,
            I => \N__15926\
        );

    \I__2778\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15923\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__15943\,
            I => \N__15920\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__15940\,
            I => \N__15911\
        );

    \I__2775\ : Span4Mux_h
    port map (
            O => \N__15935\,
            I => \N__15911\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__15932\,
            I => \N__15911\
        );

    \I__2773\ : Span4Mux_h
    port map (
            O => \N__15929\,
            I => \N__15911\
        );

    \I__2772\ : Span4Mux_h
    port map (
            O => \N__15926\,
            I => \N__15908\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__15923\,
            I => \N__15905\
        );

    \I__2770\ : Span4Mux_h
    port map (
            O => \N__15920\,
            I => \N__15900\
        );

    \I__2769\ : Span4Mux_v
    port map (
            O => \N__15911\,
            I => \N__15900\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__15908\,
            I => \tok.n4_adj_712\
        );

    \I__2767\ : Odrv12
    port map (
            O => \N__15905\,
            I => \tok.n4_adj_712\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__15900\,
            I => \tok.n4_adj_712\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__15893\,
            I => \tok.ram.n5577_cascade_\
        );

    \I__2764\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15886\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__15889\,
            I => \N__15883\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__15886\,
            I => \N__15879\
        );

    \I__2761\ : InMux
    port map (
            O => \N__15883\,
            I => \N__15876\
        );

    \I__2760\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15870\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__15879\,
            I => \N__15865\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__15876\,
            I => \N__15865\
        );

    \I__2757\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15862\
        );

    \I__2756\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15857\
        );

    \I__2755\ : InMux
    port map (
            O => \N__15873\,
            I => \N__15854\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__15870\,
            I => \N__15851\
        );

    \I__2753\ : Span4Mux_v
    port map (
            O => \N__15865\,
            I => \N__15846\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__15862\,
            I => \N__15846\
        );

    \I__2751\ : InMux
    port map (
            O => \N__15861\,
            I => \N__15843\
        );

    \I__2750\ : InMux
    port map (
            O => \N__15860\,
            I => \N__15840\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__15857\,
            I => \N__15835\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__15854\,
            I => \N__15835\
        );

    \I__2747\ : Span4Mux_v
    port map (
            O => \N__15851\,
            I => \N__15830\
        );

    \I__2746\ : Span4Mux_h
    port map (
            O => \N__15846\,
            I => \N__15830\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__15843\,
            I => \tok.n101\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__15840\,
            I => \tok.n101\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__15835\,
            I => \tok.n101\
        );

    \I__2742\ : Odrv4
    port map (
            O => \N__15830\,
            I => \tok.n101\
        );

    \I__2741\ : InMux
    port map (
            O => \N__15821\,
            I => \N__15818\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__15818\,
            I => \tok.n3_adj_672\
        );

    \I__2739\ : InMux
    port map (
            O => \N__15815\,
            I => \N__15809\
        );

    \I__2738\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15809\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__15809\,
            I => \tok.n14_adj_701\
        );

    \I__2736\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15803\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__15803\,
            I => \N__15800\
        );

    \I__2734\ : Span4Mux_h
    port map (
            O => \N__15800\,
            I => \N__15797\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__15797\,
            I => \tok.n5429\
        );

    \I__2732\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15791\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__15791\,
            I => \tok.n5406\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__15788\,
            I => \tok.n5433_cascade_\
        );

    \I__2729\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15782\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__15782\,
            I => \tok.n5272\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__2726\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__15770\,
            I => \tok.n10_adj_796\
        );

    \I__2723\ : InMux
    port map (
            O => \N__15767\,
            I => \N__15761\
        );

    \I__2722\ : InMux
    port map (
            O => \N__15766\,
            I => \N__15761\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__15761\,
            I => \tok.n14_adj_807\
        );

    \I__2720\ : InMux
    port map (
            O => \N__15758\,
            I => \N__15755\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__15755\,
            I => \tok.n5175\
        );

    \I__2718\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15749\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__15749\,
            I => \N__15745\
        );

    \I__2716\ : InMux
    port map (
            O => \N__15748\,
            I => \N__15742\
        );

    \I__2715\ : Span4Mux_h
    port map (
            O => \N__15745\,
            I => \N__15737\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__15742\,
            I => \N__15737\
        );

    \I__2713\ : Span4Mux_v
    port map (
            O => \N__15737\,
            I => \N__15734\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__15734\,
            I => n10_adj_866
        );

    \I__2711\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15728\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__15728\,
            I => \N__15723\
        );

    \I__2709\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15719\
        );

    \I__2708\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15716\
        );

    \I__2707\ : Span12Mux_v
    port map (
            O => \N__15723\,
            I => \N__15713\
        );

    \I__2706\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15710\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__15719\,
            I => \N__15707\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__15716\,
            I => \N__15704\
        );

    \I__2703\ : Odrv12
    port map (
            O => \N__15713\,
            I => tc_1
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__15710\,
            I => tc_1
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__15707\,
            I => tc_1
        );

    \I__2700\ : Odrv12
    port map (
            O => \N__15704\,
            I => tc_1
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__15695\,
            I => \N__15692\
        );

    \I__2698\ : InMux
    port map (
            O => \N__15692\,
            I => \N__15689\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__15689\,
            I => \N__15686\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__15683\,
            I => \tok.tc_1\
        );

    \I__2694\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15677\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__15677\,
            I => \tok.n2_adj_808\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__15674\,
            I => \N__15668\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__15673\,
            I => \N__15664\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__15672\,
            I => \N__15660\
        );

    \I__2689\ : InMux
    port map (
            O => \N__15671\,
            I => \N__15647\
        );

    \I__2688\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15647\
        );

    \I__2687\ : InMux
    port map (
            O => \N__15667\,
            I => \N__15647\
        );

    \I__2686\ : InMux
    port map (
            O => \N__15664\,
            I => \N__15647\
        );

    \I__2685\ : InMux
    port map (
            O => \N__15663\,
            I => \N__15647\
        );

    \I__2684\ : InMux
    port map (
            O => \N__15660\,
            I => \N__15647\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__15647\,
            I => \N__15644\
        );

    \I__2682\ : Odrv12
    port map (
            O => \N__15644\,
            I => \tok.n10_adj_747\
        );

    \I__2681\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15635\
        );

    \I__2680\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15635\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__15635\,
            I => \N__15632\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__15632\,
            I => \tok.n2635\
        );

    \I__2677\ : InMux
    port map (
            O => \N__15629\,
            I => \N__15612\
        );

    \I__2676\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15612\
        );

    \I__2675\ : InMux
    port map (
            O => \N__15627\,
            I => \N__15612\
        );

    \I__2674\ : InMux
    port map (
            O => \N__15626\,
            I => \N__15595\
        );

    \I__2673\ : InMux
    port map (
            O => \N__15625\,
            I => \N__15595\
        );

    \I__2672\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15595\
        );

    \I__2671\ : InMux
    port map (
            O => \N__15623\,
            I => \N__15595\
        );

    \I__2670\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15595\
        );

    \I__2669\ : InMux
    port map (
            O => \N__15621\,
            I => \N__15595\
        );

    \I__2668\ : InMux
    port map (
            O => \N__15620\,
            I => \N__15595\
        );

    \I__2667\ : InMux
    port map (
            O => \N__15619\,
            I => \N__15595\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__15612\,
            I => \N__15591\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__15595\,
            I => \N__15586\
        );

    \I__2664\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15583\
        );

    \I__2663\ : Span4Mux_v
    port map (
            O => \N__15591\,
            I => \N__15580\
        );

    \I__2662\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15575\
        );

    \I__2661\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15575\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__15586\,
            I => \tok.n11\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__15583\,
            I => \tok.n11\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__15580\,
            I => \tok.n11\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__15575\,
            I => \tok.n11\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__15566\,
            I => \N__15563\
        );

    \I__2655\ : InMux
    port map (
            O => \N__15563\,
            I => \N__15551\
        );

    \I__2654\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15551\
        );

    \I__2653\ : InMux
    port map (
            O => \N__15561\,
            I => \N__15551\
        );

    \I__2652\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15551\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__15551\,
            I => \N__15548\
        );

    \I__2650\ : Odrv12
    port map (
            O => \N__15548\,
            I => \tok.n2697\
        );

    \I__2649\ : InMux
    port map (
            O => \N__15545\,
            I => \N__15539\
        );

    \I__2648\ : InMux
    port map (
            O => \N__15544\,
            I => \N__15536\
        );

    \I__2647\ : InMux
    port map (
            O => \N__15543\,
            I => \N__15532\
        );

    \I__2646\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15529\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__15539\,
            I => \N__15524\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__15536\,
            I => \N__15521\
        );

    \I__2643\ : InMux
    port map (
            O => \N__15535\,
            I => \N__15518\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__15532\,
            I => \N__15512\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__15529\,
            I => \N__15512\
        );

    \I__2640\ : InMux
    port map (
            O => \N__15528\,
            I => \N__15509\
        );

    \I__2639\ : InMux
    port map (
            O => \N__15527\,
            I => \N__15505\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__15524\,
            I => \N__15500\
        );

    \I__2637\ : Span4Mux_s1_h
    port map (
            O => \N__15521\,
            I => \N__15500\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__15518\,
            I => \N__15497\
        );

    \I__2635\ : InMux
    port map (
            O => \N__15517\,
            I => \N__15494\
        );

    \I__2634\ : Span4Mux_s2_h
    port map (
            O => \N__15512\,
            I => \N__15489\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__15509\,
            I => \N__15489\
        );

    \I__2632\ : InMux
    port map (
            O => \N__15508\,
            I => \N__15486\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__15505\,
            I => \N__15483\
        );

    \I__2630\ : Span4Mux_h
    port map (
            O => \N__15500\,
            I => \N__15476\
        );

    \I__2629\ : Span4Mux_h
    port map (
            O => \N__15497\,
            I => \N__15476\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__15494\,
            I => \N__15476\
        );

    \I__2627\ : Span4Mux_h
    port map (
            O => \N__15489\,
            I => \N__15471\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__15486\,
            I => \N__15471\
        );

    \I__2625\ : Odrv12
    port map (
            O => \N__15483\,
            I => \tok.n15_adj_789\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__15476\,
            I => \tok.n15_adj_789\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__15471\,
            I => \tok.n15_adj_789\
        );

    \I__2622\ : InMux
    port map (
            O => \N__15464\,
            I => \N__15461\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__15461\,
            I => \tok.n2520\
        );

    \I__2620\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15455\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__15455\,
            I => \N__15452\
        );

    \I__2618\ : Span4Mux_v
    port map (
            O => \N__15452\,
            I => \N__15447\
        );

    \I__2617\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15442\
        );

    \I__2616\ : InMux
    port map (
            O => \N__15450\,
            I => \N__15442\
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__15447\,
            I => \tok.n10_adj_803\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__15442\,
            I => \tok.n10_adj_803\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__15437\,
            I => \tok.n2520_cascade_\
        );

    \I__2612\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15425\
        );

    \I__2611\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15425\
        );

    \I__2610\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15425\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__15425\,
            I => \N__15420\
        );

    \I__2608\ : InMux
    port map (
            O => \N__15424\,
            I => \N__15412\
        );

    \I__2607\ : InMux
    port map (
            O => \N__15423\,
            I => \N__15412\
        );

    \I__2606\ : Span4Mux_h
    port map (
            O => \N__15420\,
            I => \N__15409\
        );

    \I__2605\ : InMux
    port map (
            O => \N__15419\,
            I => \N__15402\
        );

    \I__2604\ : InMux
    port map (
            O => \N__15418\,
            I => \N__15402\
        );

    \I__2603\ : InMux
    port map (
            O => \N__15417\,
            I => \N__15402\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__15412\,
            I => \tok.n9_adj_802\
        );

    \I__2601\ : Odrv4
    port map (
            O => \N__15409\,
            I => \tok.n9_adj_802\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__15402\,
            I => \tok.n9_adj_802\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__15395\,
            I => \N__15392\
        );

    \I__2598\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15388\
        );

    \I__2597\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15385\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__15388\,
            I => \N__15382\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__15385\,
            I => \N__15379\
        );

    \I__2594\ : Span4Mux_h
    port map (
            O => \N__15382\,
            I => \N__15376\
        );

    \I__2593\ : Span4Mux_h
    port map (
            O => \N__15379\,
            I => \N__15371\
        );

    \I__2592\ : Span4Mux_v
    port map (
            O => \N__15376\,
            I => \N__15371\
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__15371\,
            I => \tok.table_rd_3\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__15368\,
            I => \tok.n2661_cascade_\
        );

    \I__2589\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15362\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__15362\,
            I => \tok.n10_adj_845\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__15359\,
            I => \tok.n9_adj_847_cascade_\
        );

    \I__2586\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15350\
        );

    \I__2585\ : InMux
    port map (
            O => \N__15355\,
            I => \N__15350\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__15350\,
            I => uart_rx_data_6
        );

    \I__2583\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__15344\,
            I => \tok.n6_adj_843\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__15341\,
            I => \tok.n31_adj_844_cascade_\
        );

    \I__2580\ : InMux
    port map (
            O => \N__15338\,
            I => \N__15332\
        );

    \I__2579\ : InMux
    port map (
            O => \N__15337\,
            I => \N__15332\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__15332\,
            I => uart_rx_data_3
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__2576\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15317\
        );

    \I__2575\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15317\
        );

    \I__2574\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15317\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__15317\,
            I => capture_4
        );

    \I__2572\ : InMux
    port map (
            O => \N__15314\,
            I => \N__15308\
        );

    \I__2571\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15303\
        );

    \I__2570\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15303\
        );

    \I__2569\ : InMux
    port map (
            O => \N__15311\,
            I => \N__15300\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__15308\,
            I => \N__15295\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15295\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__15300\,
            I => \tok.tc_plus_1_6\
        );

    \I__2565\ : Odrv12
    port map (
            O => \N__15295\,
            I => \tok.tc_plus_1_6\
        );

    \I__2564\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15287\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__15287\,
            I => \N__15284\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__15284\,
            I => \N__15281\
        );

    \I__2561\ : Span4Mux_h
    port map (
            O => \N__15281\,
            I => \N__15278\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__15278\,
            I => \tok.table_wr_data_6\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__15275\,
            I => \N__15271\
        );

    \I__2558\ : InMux
    port map (
            O => \N__15274\,
            I => \N__15266\
        );

    \I__2557\ : InMux
    port map (
            O => \N__15271\,
            I => \N__15266\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__15266\,
            I => \N__15263\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__15263\,
            I => \N__15260\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__15260\,
            I => \tok.key_rd_8\
        );

    \I__2553\ : InMux
    port map (
            O => \N__15257\,
            I => \N__15254\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__15254\,
            I => \tok.n28_adj_755\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__15251\,
            I => \tok.n26_adj_756_cascade_\
        );

    \I__2550\ : InMux
    port map (
            O => \N__15248\,
            I => \N__15245\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__15245\,
            I => \tok.n27_adj_757\
        );

    \I__2548\ : InMux
    port map (
            O => \N__15242\,
            I => \N__15239\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__15239\,
            I => \tok.found_slot_N_145\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__15236\,
            I => \N__15226\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__15235\,
            I => \N__15223\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__15234\,
            I => \N__15220\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__15233\,
            I => \N__15217\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__15232\,
            I => \N__15214\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__15231\,
            I => \N__15211\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__15230\,
            I => \N__15208\
        );

    \I__2539\ : CascadeMux
    port map (
            O => \N__15229\,
            I => \N__15205\
        );

    \I__2538\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15196\
        );

    \I__2537\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15196\
        );

    \I__2536\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15196\
        );

    \I__2535\ : InMux
    port map (
            O => \N__15217\,
            I => \N__15196\
        );

    \I__2534\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15187\
        );

    \I__2533\ : InMux
    port map (
            O => \N__15211\,
            I => \N__15187\
        );

    \I__2532\ : InMux
    port map (
            O => \N__15208\,
            I => \N__15187\
        );

    \I__2531\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15187\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__15196\,
            I => \N__15180\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__15187\,
            I => \N__15180\
        );

    \I__2528\ : InMux
    port map (
            O => \N__15186\,
            I => \N__15177\
        );

    \I__2527\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15174\
        );

    \I__2526\ : Span4Mux_s2_v
    port map (
            O => \N__15180\,
            I => \N__15169\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__15177\,
            I => \N__15169\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__15174\,
            I => \tok.found_slot\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__15169\,
            I => \tok.found_slot\
        );

    \I__2522\ : SRMux
    port map (
            O => \N__15164\,
            I => \N__15160\
        );

    \I__2521\ : SRMux
    port map (
            O => \N__15163\,
            I => \N__15157\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__15160\,
            I => \N__15152\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__15157\,
            I => \N__15152\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__15152\,
            I => \N__15149\
        );

    \I__2517\ : Span4Mux_h
    port map (
            O => \N__15149\,
            I => \N__15146\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__15146\,
            I => \tok.write_slot\
        );

    \I__2515\ : InMux
    port map (
            O => \N__15143\,
            I => \N__15137\
        );

    \I__2514\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15137\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__15137\,
            I => \N__15134\
        );

    \I__2512\ : Span4Mux_h
    port map (
            O => \N__15134\,
            I => \N__15131\
        );

    \I__2511\ : Odrv4
    port map (
            O => \N__15131\,
            I => \tok.key_rd_3\
        );

    \I__2510\ : InMux
    port map (
            O => \N__15128\,
            I => \N__15122\
        );

    \I__2509\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15122\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__15122\,
            I => \N__15119\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__15119\,
            I => \N__15116\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__15116\,
            I => \tok.key_rd_5\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__15113\,
            I => \N__15110\
        );

    \I__2504\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15107\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__15107\,
            I => \tok.n20\
        );

    \I__2502\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15101\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__15101\,
            I => \tok.n18_adj_759\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__15098\,
            I => \N__15095\
        );

    \I__2499\ : InMux
    port map (
            O => \N__15095\,
            I => \N__15089\
        );

    \I__2498\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15089\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__15089\,
            I => \N__15086\
        );

    \I__2496\ : Span4Mux_h
    port map (
            O => \N__15086\,
            I => \N__15083\
        );

    \I__2495\ : Odrv4
    port map (
            O => \N__15083\,
            I => \tok.key_rd_1\
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__2493\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15071\
        );

    \I__2492\ : InMux
    port map (
            O => \N__15076\,
            I => \N__15071\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__15071\,
            I => \N__15068\
        );

    \I__2490\ : Span4Mux_h
    port map (
            O => \N__15068\,
            I => \N__15065\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__15065\,
            I => \tok.key_rd_4\
        );

    \I__2488\ : InMux
    port map (
            O => \N__15062\,
            I => \N__15059\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__15059\,
            I => \tok.n25_adj_758\
        );

    \I__2486\ : InMux
    port map (
            O => \N__15056\,
            I => \N__15050\
        );

    \I__2485\ : InMux
    port map (
            O => \N__15055\,
            I => \N__15050\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__15050\,
            I => \N__15047\
        );

    \I__2483\ : Span4Mux_h
    port map (
            O => \N__15047\,
            I => \N__15044\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__15044\,
            I => \tok.key_rd_0\
        );

    \I__2481\ : InMux
    port map (
            O => \N__15041\,
            I => \N__15035\
        );

    \I__2480\ : InMux
    port map (
            O => \N__15040\,
            I => \N__15035\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__15035\,
            I => \N__15032\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__15032\,
            I => \N__15029\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__15029\,
            I => \tok.key_rd_6\
        );

    \I__2476\ : InMux
    port map (
            O => \N__15026\,
            I => \N__15023\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__15023\,
            I => \tok.n5590\
        );

    \I__2474\ : InMux
    port map (
            O => \N__15020\,
            I => \N__15010\
        );

    \I__2473\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15010\
        );

    \I__2472\ : InMux
    port map (
            O => \N__15018\,
            I => \N__15010\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__15017\,
            I => \N__15007\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__15010\,
            I => \N__15004\
        );

    \I__2469\ : InMux
    port map (
            O => \N__15007\,
            I => \N__15001\
        );

    \I__2468\ : Span12Mux_s6_v
    port map (
            O => \N__15004\,
            I => \N__14998\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__15001\,
            I => \tok.c_stk_r_3\
        );

    \I__2466\ : Odrv12
    port map (
            O => \N__14998\,
            I => \tok.c_stk_r_3\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__14993\,
            I => \tok.ram.n5580_cascade_\
        );

    \I__2464\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14987\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__14987\,
            I => \tok.n5460\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__14984\,
            I => \tok.n3_adj_659_cascade_\
        );

    \I__2461\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14978\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__14978\,
            I => \N__14973\
        );

    \I__2459\ : InMux
    port map (
            O => \N__14977\,
            I => \N__14968\
        );

    \I__2458\ : InMux
    port map (
            O => \N__14976\,
            I => \N__14968\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__14973\,
            I => \N__14964\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__14968\,
            I => \N__14961\
        );

    \I__2455\ : InMux
    port map (
            O => \N__14967\,
            I => \N__14958\
        );

    \I__2454\ : Span4Mux_h
    port map (
            O => \N__14964\,
            I => \N__14953\
        );

    \I__2453\ : Span4Mux_h
    port map (
            O => \N__14961\,
            I => \N__14953\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__14958\,
            I => \tok.tc_plus_1_3\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__14953\,
            I => \tok.tc_plus_1_3\
        );

    \I__2450\ : CascadeMux
    port map (
            O => \N__14948\,
            I => \tok.n13_adj_660_cascade_\
        );

    \I__2449\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14939\
        );

    \I__2448\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14939\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__14939\,
            I => \N__14936\
        );

    \I__2446\ : Span4Mux_h
    port map (
            O => \N__14936\,
            I => \N__14933\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__14933\,
            I => n92_adj_867
        );

    \I__2444\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14927\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__2442\ : Span4Mux_v
    port map (
            O => \N__14924\,
            I => \N__14920\
        );

    \I__2441\ : InMux
    port map (
            O => \N__14923\,
            I => \N__14917\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__14920\,
            I => \tok.n17_adj_777\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__14917\,
            I => \tok.n17_adj_777\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__14912\,
            I => \tok.n4_adj_778_cascade_\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__14909\,
            I => \tok.n26_adj_760_cascade_\
        );

    \I__2436\ : InMux
    port map (
            O => \N__14906\,
            I => \N__14903\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__14903\,
            I => \tok.n30_adj_761\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__14900\,
            I => \tok.n5587_cascade_\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__14897\,
            I => \tok.n5_cascade_\
        );

    \I__2432\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__14891\,
            I => \tok.n5\
        );

    \I__2430\ : InMux
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__14885\,
            I => \tok.n33\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__14882\,
            I => \tok.n27_cascade_\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__14879\,
            I => \N__14876\
        );

    \I__2426\ : CascadeBuf
    port map (
            O => \N__14876\,
            I => \N__14872\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__14875\,
            I => \N__14869\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__14872\,
            I => \N__14866\
        );

    \I__2423\ : CascadeBuf
    port map (
            O => \N__14869\,
            I => \N__14863\
        );

    \I__2422\ : InMux
    port map (
            O => \N__14866\,
            I => \N__14860\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__14863\,
            I => \N__14857\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__14860\,
            I => \N__14854\
        );

    \I__2419\ : InMux
    port map (
            O => \N__14857\,
            I => \N__14851\
        );

    \I__2418\ : Span4Mux_h
    port map (
            O => \N__14854\,
            I => \N__14845\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__14851\,
            I => \N__14842\
        );

    \I__2416\ : InMux
    port map (
            O => \N__14850\,
            I => \N__14839\
        );

    \I__2415\ : InMux
    port map (
            O => \N__14849\,
            I => \N__14836\
        );

    \I__2414\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14833\
        );

    \I__2413\ : Span4Mux_v
    port map (
            O => \N__14845\,
            I => \N__14830\
        );

    \I__2412\ : Span12Mux_s6_h
    port map (
            O => \N__14842\,
            I => \N__14827\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__14839\,
            I => \tok.idx_0\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__14836\,
            I => \tok.idx_0\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__14833\,
            I => \tok.idx_0\
        );

    \I__2408\ : Odrv4
    port map (
            O => \N__14830\,
            I => \tok.idx_0\
        );

    \I__2407\ : Odrv12
    port map (
            O => \N__14827\,
            I => \tok.idx_0\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__14816\,
            I => \tok.n83_adj_652_cascade_\
        );

    \I__2405\ : InMux
    port map (
            O => \N__14813\,
            I => \bfn_6_3_0_\
        );

    \I__2404\ : InMux
    port map (
            O => \N__14810\,
            I => \tok.n4747\
        );

    \I__2403\ : InMux
    port map (
            O => \N__14807\,
            I => \tok.n4748\
        );

    \I__2402\ : InMux
    port map (
            O => \N__14804\,
            I => \tok.n4749\
        );

    \I__2401\ : CascadeMux
    port map (
            O => \N__14801\,
            I => \N__14798\
        );

    \I__2400\ : CascadeBuf
    port map (
            O => \N__14798\,
            I => \N__14794\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__14797\,
            I => \N__14791\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__14794\,
            I => \N__14788\
        );

    \I__2397\ : CascadeBuf
    port map (
            O => \N__14791\,
            I => \N__14785\
        );

    \I__2396\ : InMux
    port map (
            O => \N__14788\,
            I => \N__14782\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__14785\,
            I => \N__14779\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__14782\,
            I => \N__14775\
        );

    \I__2393\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14772\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__14778\,
            I => \N__14769\
        );

    \I__2391\ : Span4Mux_h
    port map (
            O => \N__14775\,
            I => \N__14764\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__14772\,
            I => \N__14761\
        );

    \I__2389\ : InMux
    port map (
            O => \N__14769\,
            I => \N__14758\
        );

    \I__2388\ : InMux
    port map (
            O => \N__14768\,
            I => \N__14755\
        );

    \I__2387\ : InMux
    port map (
            O => \N__14767\,
            I => \N__14752\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__14764\,
            I => \N__14749\
        );

    \I__2385\ : Span12Mux_s5_h
    port map (
            O => \N__14761\,
            I => \N__14746\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__14758\,
            I => \tok.idx_4\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__14755\,
            I => \tok.idx_4\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__14752\,
            I => \tok.idx_4\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__14749\,
            I => \tok.idx_4\
        );

    \I__2380\ : Odrv12
    port map (
            O => \N__14746\,
            I => \tok.idx_4\
        );

    \I__2379\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__14732\,
            I => \tok.n33_adj_819\
        );

    \I__2377\ : InMux
    port map (
            O => \N__14729\,
            I => \tok.n4750\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__14726\,
            I => \N__14723\
        );

    \I__2375\ : CascadeBuf
    port map (
            O => \N__14723\,
            I => \N__14719\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__14722\,
            I => \N__14716\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__14719\,
            I => \N__14713\
        );

    \I__2372\ : CascadeBuf
    port map (
            O => \N__14716\,
            I => \N__14710\
        );

    \I__2371\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14707\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__14710\,
            I => \N__14704\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__14707\,
            I => \N__14701\
        );

    \I__2368\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14698\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__14701\,
            I => \N__14692\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__14698\,
            I => \N__14689\
        );

    \I__2365\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14686\
        );

    \I__2364\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14683\
        );

    \I__2363\ : InMux
    port map (
            O => \N__14695\,
            I => \N__14680\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__14692\,
            I => \N__14677\
        );

    \I__2361\ : Span4Mux_h
    port map (
            O => \N__14689\,
            I => \N__14674\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__14686\,
            I => \N__14665\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__14683\,
            I => \N__14665\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__14680\,
            I => \N__14665\
        );

    \I__2357\ : Span4Mux_s2_v
    port map (
            O => \N__14677\,
            I => \N__14665\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__14674\,
            I => \N__14662\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__14665\,
            I => \tok.idx_5\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__14662\,
            I => \tok.idx_5\
        );

    \I__2353\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14654\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__14654\,
            I => \tok.n33_adj_811\
        );

    \I__2351\ : InMux
    port map (
            O => \N__14651\,
            I => \tok.n4751\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__14648\,
            I => \N__14644\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__14647\,
            I => \N__14641\
        );

    \I__2348\ : CascadeBuf
    port map (
            O => \N__14644\,
            I => \N__14638\
        );

    \I__2347\ : CascadeBuf
    port map (
            O => \N__14641\,
            I => \N__14635\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__14638\,
            I => \N__14632\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__14635\,
            I => \N__14629\
        );

    \I__2344\ : InMux
    port map (
            O => \N__14632\,
            I => \N__14626\
        );

    \I__2343\ : InMux
    port map (
            O => \N__14629\,
            I => \N__14623\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__14626\,
            I => \N__14619\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__14623\,
            I => \N__14616\
        );

    \I__2340\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14611\
        );

    \I__2339\ : Span4Mux_v
    port map (
            O => \N__14619\,
            I => \N__14608\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__14616\,
            I => \N__14605\
        );

    \I__2337\ : InMux
    port map (
            O => \N__14615\,
            I => \N__14602\
        );

    \I__2336\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14599\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__14611\,
            I => \N__14594\
        );

    \I__2334\ : Span4Mux_v
    port map (
            O => \N__14608\,
            I => \N__14594\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__14605\,
            I => \N__14591\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__14602\,
            I => \tok.idx_6\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__14599\,
            I => \tok.idx_6\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__14594\,
            I => \tok.idx_6\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__14591\,
            I => \tok.idx_6\
        );

    \I__2328\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14579\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__14579\,
            I => \tok.n33_adj_804\
        );

    \I__2326\ : InMux
    port map (
            O => \N__14576\,
            I => \tok.n4752\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__14573\,
            I => \N__14569\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__14572\,
            I => \N__14566\
        );

    \I__2323\ : CascadeBuf
    port map (
            O => \N__14569\,
            I => \N__14563\
        );

    \I__2322\ : CascadeBuf
    port map (
            O => \N__14566\,
            I => \N__14560\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__14563\,
            I => \N__14557\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__14560\,
            I => \N__14554\
        );

    \I__2319\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14549\
        );

    \I__2318\ : InMux
    port map (
            O => \N__14554\,
            I => \N__14546\
        );

    \I__2317\ : InMux
    port map (
            O => \N__14553\,
            I => \N__14542\
        );

    \I__2316\ : InMux
    port map (
            O => \N__14552\,
            I => \N__14539\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__14549\,
            I => \N__14534\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__14546\,
            I => \N__14534\
        );

    \I__2313\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14531\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__14542\,
            I => \N__14526\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__14539\,
            I => \N__14526\
        );

    \I__2310\ : Span12Mux_s11_v
    port map (
            O => \N__14534\,
            I => \N__14523\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__14531\,
            I => \tok.idx_7\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__14526\,
            I => \tok.idx_7\
        );

    \I__2307\ : Odrv12
    port map (
            O => \N__14523\,
            I => \tok.idx_7\
        );

    \I__2306\ : InMux
    port map (
            O => \N__14516\,
            I => \tok.n4753\
        );

    \I__2305\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14510\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__14510\,
            I => \tok.n33_adj_801\
        );

    \I__2303\ : InMux
    port map (
            O => \N__14507\,
            I => \N__14504\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__14504\,
            I => \N__14501\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__14501\,
            I => reset_c
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__14498\,
            I => \N__14495\
        );

    \I__2299\ : InMux
    port map (
            O => \N__14495\,
            I => \N__14489\
        );

    \I__2298\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14489\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__14489\,
            I => \tok.A_stk.tail_16\
        );

    \I__2296\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14480\
        );

    \I__2295\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14480\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__14480\,
            I => \tok.A_stk.tail_32\
        );

    \I__2293\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14471\
        );

    \I__2292\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14471\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__14471\,
            I => \tok.A_stk.tail_48\
        );

    \I__2290\ : InMux
    port map (
            O => \N__14468\,
            I => \N__14462\
        );

    \I__2289\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14462\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__14462\,
            I => \tok.A_stk.tail_64\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__14459\,
            I => \N__14455\
        );

    \I__2286\ : InMux
    port map (
            O => \N__14458\,
            I => \N__14452\
        );

    \I__2285\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14449\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__14452\,
            I => \N__14444\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__14449\,
            I => \N__14444\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__14444\,
            I => tail_112
        );

    \I__2281\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14435\
        );

    \I__2280\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14435\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__14435\,
            I => \tok.A_stk.tail_80\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__14432\,
            I => \N__14428\
        );

    \I__2277\ : InMux
    port map (
            O => \N__14431\,
            I => \N__14425\
        );

    \I__2276\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14422\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__14425\,
            I => tail_96
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__14422\,
            I => tail_96
        );

    \I__2273\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14411\
        );

    \I__2272\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14411\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__14411\,
            I => \tok.A_stk.tail_0\
        );

    \I__2270\ : InMux
    port map (
            O => \N__14408\,
            I => \N__14405\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__14405\,
            I => \N__14402\
        );

    \I__2268\ : Span4Mux_h
    port map (
            O => \N__14402\,
            I => \N__14398\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__14401\,
            I => \N__14395\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__14398\,
            I => \N__14392\
        );

    \I__2265\ : InMux
    port map (
            O => \N__14395\,
            I => \N__14389\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__14392\,
            I => \N__14386\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__14389\,
            I => sender_9
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__14386\,
            I => sender_9
        );

    \I__2261\ : SRMux
    port map (
            O => \N__14381\,
            I => \N__14378\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__14378\,
            I => \N__14375\
        );

    \I__2259\ : Span4Mux_s3_h
    port map (
            O => \N__14375\,
            I => \N__14362\
        );

    \I__2258\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14357\
        );

    \I__2257\ : InMux
    port map (
            O => \N__14373\,
            I => \N__14357\
        );

    \I__2256\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14342\
        );

    \I__2255\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14342\
        );

    \I__2254\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14342\
        );

    \I__2253\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14342\
        );

    \I__2252\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14342\
        );

    \I__2251\ : InMux
    port map (
            O => \N__14367\,
            I => \N__14342\
        );

    \I__2250\ : InMux
    port map (
            O => \N__14366\,
            I => \N__14342\
        );

    \I__2249\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14339\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__14362\,
            I => \N__14336\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__14357\,
            I => \N__14333\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14329\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__14339\,
            I => \N__14326\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__14336\,
            I => \N__14321\
        );

    \I__2243\ : Span4Mux_v
    port map (
            O => \N__14333\,
            I => \N__14321\
        );

    \I__2242\ : InMux
    port map (
            O => \N__14332\,
            I => \N__14318\
        );

    \I__2241\ : Span4Mux_v
    port map (
            O => \N__14329\,
            I => \N__14313\
        );

    \I__2240\ : Span4Mux_h
    port map (
            O => \N__14326\,
            I => \N__14313\
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__14321\,
            I => n23
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__14318\,
            I => n23
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__14313\,
            I => n23
        );

    \I__2236\ : InMux
    port map (
            O => \N__14306\,
            I => \N__14303\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__14303\,
            I => \tok.uart.sender_8\
        );

    \I__2234\ : CEMux
    port map (
            O => \N__14300\,
            I => \N__14297\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__14297\,
            I => \N__14294\
        );

    \I__2232\ : Span4Mux_h
    port map (
            O => \N__14294\,
            I => \N__14290\
        );

    \I__2231\ : CEMux
    port map (
            O => \N__14293\,
            I => \N__14287\
        );

    \I__2230\ : Span4Mux_v
    port map (
            O => \N__14290\,
            I => \N__14284\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__14287\,
            I => \N__14281\
        );

    \I__2228\ : Span4Mux_s2_h
    port map (
            O => \N__14284\,
            I => \N__14278\
        );

    \I__2227\ : Span12Mux_s4_v
    port map (
            O => \N__14281\,
            I => \N__14275\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__14278\,
            I => \tok.uart.n1017\
        );

    \I__2225\ : Odrv12
    port map (
            O => \N__14275\,
            I => \tok.uart.n1017\
        );

    \I__2224\ : InMux
    port map (
            O => \N__14270\,
            I => \N__14266\
        );

    \I__2223\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14261\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__14266\,
            I => \N__14257\
        );

    \I__2221\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14252\
        );

    \I__2220\ : InMux
    port map (
            O => \N__14264\,
            I => \N__14248\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__14261\,
            I => \N__14245\
        );

    \I__2218\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14242\
        );

    \I__2217\ : Span4Mux_s3_v
    port map (
            O => \N__14257\,
            I => \N__14239\
        );

    \I__2216\ : InMux
    port map (
            O => \N__14256\,
            I => \N__14236\
        );

    \I__2215\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14233\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__14252\,
            I => \N__14230\
        );

    \I__2213\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14227\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__14248\,
            I => \N__14220\
        );

    \I__2211\ : Span4Mux_h
    port map (
            O => \N__14245\,
            I => \N__14220\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__14242\,
            I => \N__14220\
        );

    \I__2209\ : Span4Mux_h
    port map (
            O => \N__14239\,
            I => \N__14213\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__14236\,
            I => \N__14213\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__14233\,
            I => \N__14213\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__14230\,
            I => \tok.C_stk.n602\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__14227\,
            I => \tok.C_stk.n602\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__14220\,
            I => \tok.C_stk.n602\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__14213\,
            I => \tok.C_stk.n602\
        );

    \I__2202\ : InMux
    port map (
            O => \N__14204\,
            I => \N__14201\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__14201\,
            I => \N__14198\
        );

    \I__2200\ : IoSpan4Mux
    port map (
            O => \N__14198\,
            I => \N__14192\
        );

    \I__2199\ : InMux
    port map (
            O => \N__14197\,
            I => \N__14189\
        );

    \I__2198\ : InMux
    port map (
            O => \N__14196\,
            I => \N__14182\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__14195\,
            I => \N__14179\
        );

    \I__2196\ : Span4Mux_s3_v
    port map (
            O => \N__14192\,
            I => \N__14174\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__14189\,
            I => \N__14174\
        );

    \I__2194\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14171\
        );

    \I__2193\ : InMux
    port map (
            O => \N__14187\,
            I => \N__14168\
        );

    \I__2192\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14165\
        );

    \I__2191\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14161\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__14182\,
            I => \N__14158\
        );

    \I__2189\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14155\
        );

    \I__2188\ : Span4Mux_v
    port map (
            O => \N__14174\,
            I => \N__14146\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__14171\,
            I => \N__14146\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__14168\,
            I => \N__14146\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__14165\,
            I => \N__14146\
        );

    \I__2184\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14143\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__14161\,
            I => \N__14140\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__14158\,
            I => \N__14135\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__14155\,
            I => \N__14135\
        );

    \I__2180\ : Span4Mux_h
    port map (
            O => \N__14146\,
            I => \N__14132\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__14143\,
            I => \N__14129\
        );

    \I__2178\ : Span4Mux_v
    port map (
            O => \N__14140\,
            I => \N__14124\
        );

    \I__2177\ : Span4Mux_h
    port map (
            O => \N__14135\,
            I => \N__14124\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__14132\,
            I => \tok.n241\
        );

    \I__2175\ : Odrv12
    port map (
            O => \N__14129\,
            I => \tok.n241\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__14124\,
            I => \tok.n241\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__14117\,
            I => \tok.C_stk.n5438_cascade_\
        );

    \I__2172\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14109\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__14113\,
            I => \N__14106\
        );

    \I__2170\ : InMux
    port map (
            O => \N__14112\,
            I => \N__14102\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__14109\,
            I => \N__14099\
        );

    \I__2168\ : InMux
    port map (
            O => \N__14106\,
            I => \N__14094\
        );

    \I__2167\ : InMux
    port map (
            O => \N__14105\,
            I => \N__14094\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__14102\,
            I => \N__14091\
        );

    \I__2165\ : Odrv12
    port map (
            O => \N__14099\,
            I => tc_6
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__14094\,
            I => tc_6
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__14091\,
            I => tc_6
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__14084\,
            I => \N__14080\
        );

    \I__2161\ : InMux
    port map (
            O => \N__14083\,
            I => \N__14076\
        );

    \I__2160\ : InMux
    port map (
            O => \N__14080\,
            I => \N__14071\
        );

    \I__2159\ : InMux
    port map (
            O => \N__14079\,
            I => \N__14071\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__14076\,
            I => \N__14065\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__14071\,
            I => \N__14065\
        );

    \I__2156\ : InMux
    port map (
            O => \N__14070\,
            I => \N__14062\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__14065\,
            I => \N__14059\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__14062\,
            I => \tok.c_stk_r_6\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__14059\,
            I => \tok.c_stk_r_6\
        );

    \I__2152\ : InMux
    port map (
            O => \N__14054\,
            I => \N__14048\
        );

    \I__2151\ : InMux
    port map (
            O => \N__14053\,
            I => \N__14048\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__14048\,
            I => \tok.C_stk.tail_6\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__14045\,
            I => \N__14041\
        );

    \I__2148\ : InMux
    port map (
            O => \N__14044\,
            I => \N__13991\
        );

    \I__2147\ : InMux
    port map (
            O => \N__14041\,
            I => \N__13988\
        );

    \I__2146\ : InMux
    port map (
            O => \N__14040\,
            I => \N__13983\
        );

    \I__2145\ : InMux
    port map (
            O => \N__14039\,
            I => \N__13983\
        );

    \I__2144\ : InMux
    port map (
            O => \N__14038\,
            I => \N__13980\
        );

    \I__2143\ : InMux
    port map (
            O => \N__14037\,
            I => \N__13963\
        );

    \I__2142\ : InMux
    port map (
            O => \N__14036\,
            I => \N__13963\
        );

    \I__2141\ : InMux
    port map (
            O => \N__14035\,
            I => \N__13963\
        );

    \I__2140\ : InMux
    port map (
            O => \N__14034\,
            I => \N__13963\
        );

    \I__2139\ : InMux
    port map (
            O => \N__14033\,
            I => \N__13963\
        );

    \I__2138\ : InMux
    port map (
            O => \N__14032\,
            I => \N__13963\
        );

    \I__2137\ : InMux
    port map (
            O => \N__14031\,
            I => \N__13950\
        );

    \I__2136\ : InMux
    port map (
            O => \N__14030\,
            I => \N__13950\
        );

    \I__2135\ : InMux
    port map (
            O => \N__14029\,
            I => \N__13950\
        );

    \I__2134\ : InMux
    port map (
            O => \N__14028\,
            I => \N__13950\
        );

    \I__2133\ : InMux
    port map (
            O => \N__14027\,
            I => \N__13950\
        );

    \I__2132\ : InMux
    port map (
            O => \N__14026\,
            I => \N__13950\
        );

    \I__2131\ : InMux
    port map (
            O => \N__14025\,
            I => \N__13943\
        );

    \I__2130\ : InMux
    port map (
            O => \N__14024\,
            I => \N__13943\
        );

    \I__2129\ : InMux
    port map (
            O => \N__14023\,
            I => \N__13943\
        );

    \I__2128\ : InMux
    port map (
            O => \N__14022\,
            I => \N__13930\
        );

    \I__2127\ : InMux
    port map (
            O => \N__14021\,
            I => \N__13930\
        );

    \I__2126\ : InMux
    port map (
            O => \N__14020\,
            I => \N__13930\
        );

    \I__2125\ : InMux
    port map (
            O => \N__14019\,
            I => \N__13930\
        );

    \I__2124\ : InMux
    port map (
            O => \N__14018\,
            I => \N__13930\
        );

    \I__2123\ : InMux
    port map (
            O => \N__14017\,
            I => \N__13930\
        );

    \I__2122\ : InMux
    port map (
            O => \N__14016\,
            I => \N__13921\
        );

    \I__2121\ : InMux
    port map (
            O => \N__14015\,
            I => \N__13921\
        );

    \I__2120\ : InMux
    port map (
            O => \N__14014\,
            I => \N__13921\
        );

    \I__2119\ : InMux
    port map (
            O => \N__14013\,
            I => \N__13921\
        );

    \I__2118\ : InMux
    port map (
            O => \N__14012\,
            I => \N__13908\
        );

    \I__2117\ : InMux
    port map (
            O => \N__14011\,
            I => \N__13908\
        );

    \I__2116\ : InMux
    port map (
            O => \N__14010\,
            I => \N__13908\
        );

    \I__2115\ : InMux
    port map (
            O => \N__14009\,
            I => \N__13908\
        );

    \I__2114\ : InMux
    port map (
            O => \N__14008\,
            I => \N__13908\
        );

    \I__2113\ : InMux
    port map (
            O => \N__14007\,
            I => \N__13908\
        );

    \I__2112\ : InMux
    port map (
            O => \N__14006\,
            I => \N__13893\
        );

    \I__2111\ : InMux
    port map (
            O => \N__14005\,
            I => \N__13880\
        );

    \I__2110\ : InMux
    port map (
            O => \N__14004\,
            I => \N__13880\
        );

    \I__2109\ : InMux
    port map (
            O => \N__14003\,
            I => \N__13880\
        );

    \I__2108\ : InMux
    port map (
            O => \N__14002\,
            I => \N__13880\
        );

    \I__2107\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13880\
        );

    \I__2106\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13880\
        );

    \I__2105\ : InMux
    port map (
            O => \N__13999\,
            I => \N__13867\
        );

    \I__2104\ : InMux
    port map (
            O => \N__13998\,
            I => \N__13867\
        );

    \I__2103\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13867\
        );

    \I__2102\ : InMux
    port map (
            O => \N__13996\,
            I => \N__13867\
        );

    \I__2101\ : InMux
    port map (
            O => \N__13995\,
            I => \N__13867\
        );

    \I__2100\ : InMux
    port map (
            O => \N__13994\,
            I => \N__13867\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__13991\,
            I => \N__13864\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__13988\,
            I => \N__13859\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__13983\,
            I => \N__13859\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__13980\,
            I => \N__13856\
        );

    \I__2095\ : InMux
    port map (
            O => \N__13979\,
            I => \N__13847\
        );

    \I__2094\ : InMux
    port map (
            O => \N__13978\,
            I => \N__13847\
        );

    \I__2093\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13847\
        );

    \I__2092\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13847\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__13963\,
            I => \N__13842\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__13950\,
            I => \N__13842\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__13943\,
            I => \N__13839\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__13930\,
            I => \N__13836\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__13921\,
            I => \N__13833\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__13908\,
            I => \N__13830\
        );

    \I__2085\ : InMux
    port map (
            O => \N__13907\,
            I => \N__13817\
        );

    \I__2084\ : InMux
    port map (
            O => \N__13906\,
            I => \N__13817\
        );

    \I__2083\ : InMux
    port map (
            O => \N__13905\,
            I => \N__13817\
        );

    \I__2082\ : InMux
    port map (
            O => \N__13904\,
            I => \N__13817\
        );

    \I__2081\ : InMux
    port map (
            O => \N__13903\,
            I => \N__13817\
        );

    \I__2080\ : InMux
    port map (
            O => \N__13902\,
            I => \N__13817\
        );

    \I__2079\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13804\
        );

    \I__2078\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13804\
        );

    \I__2077\ : InMux
    port map (
            O => \N__13899\,
            I => \N__13804\
        );

    \I__2076\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13804\
        );

    \I__2075\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13804\
        );

    \I__2074\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13804\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__13893\,
            I => \N__13801\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__13880\,
            I => \N__13794\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__13867\,
            I => \N__13794\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__13864\,
            I => \N__13794\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__13859\,
            I => \N__13785\
        );

    \I__2068\ : Span4Mux_s1_h
    port map (
            O => \N__13856\,
            I => \N__13785\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__13847\,
            I => \N__13785\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__13842\,
            I => \N__13785\
        );

    \I__2065\ : Span4Mux_h
    port map (
            O => \N__13839\,
            I => \N__13778\
        );

    \I__2064\ : Span4Mux_h
    port map (
            O => \N__13836\,
            I => \N__13778\
        );

    \I__2063\ : Span4Mux_h
    port map (
            O => \N__13833\,
            I => \N__13778\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__13830\,
            I => \N__13773\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__13817\,
            I => \N__13773\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__13804\,
            I => \N__13770\
        );

    \I__2059\ : Span4Mux_v
    port map (
            O => \N__13801\,
            I => \N__13765\
        );

    \I__2058\ : Span4Mux_v
    port map (
            O => \N__13794\,
            I => \N__13765\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__13785\,
            I => \N__13762\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__13778\,
            I => \N__13757\
        );

    \I__2055\ : Span4Mux_h
    port map (
            O => \N__13773\,
            I => \N__13757\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__13770\,
            I => \tok.n2515\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__13765\,
            I => \tok.n2515\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__13762\,
            I => \tok.n2515\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__13757\,
            I => \tok.n2515\
        );

    \I__2050\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13742\
        );

    \I__2049\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13742\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__13742\,
            I => \tok.tail_14\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__13739\,
            I => \N__13736\
        );

    \I__2046\ : InMux
    port map (
            O => \N__13736\,
            I => \N__13733\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__13733\,
            I => \N__13729\
        );

    \I__2044\ : InMux
    port map (
            O => \N__13732\,
            I => \N__13726\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__13729\,
            I => \tok.tail_30\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__13726\,
            I => \tok.tail_30\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__13721\,
            I => \N__13717\
        );

    \I__2040\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13708\
        );

    \I__2039\ : InMux
    port map (
            O => \N__13717\,
            I => \N__13703\
        );

    \I__2038\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13703\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__13715\,
            I => \N__13700\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__13714\,
            I => \N__13697\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__13713\,
            I => \N__13678\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__13712\,
            I => \N__13675\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__13711\,
            I => \N__13672\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__13708\,
            I => \N__13658\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__13703\,
            I => \N__13658\
        );

    \I__2030\ : InMux
    port map (
            O => \N__13700\,
            I => \N__13649\
        );

    \I__2029\ : InMux
    port map (
            O => \N__13697\,
            I => \N__13649\
        );

    \I__2028\ : InMux
    port map (
            O => \N__13696\,
            I => \N__13649\
        );

    \I__2027\ : InMux
    port map (
            O => \N__13695\,
            I => \N__13649\
        );

    \I__2026\ : InMux
    port map (
            O => \N__13694\,
            I => \N__13639\
        );

    \I__2025\ : InMux
    port map (
            O => \N__13693\,
            I => \N__13636\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__13692\,
            I => \N__13628\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__13691\,
            I => \N__13624\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__13690\,
            I => \N__13619\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__13689\,
            I => \N__13616\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__13688\,
            I => \N__13613\
        );

    \I__2019\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13590\
        );

    \I__2018\ : InMux
    port map (
            O => \N__13686\,
            I => \N__13590\
        );

    \I__2017\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13590\
        );

    \I__2016\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13590\
        );

    \I__2015\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13583\
        );

    \I__2014\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13583\
        );

    \I__2013\ : InMux
    port map (
            O => \N__13681\,
            I => \N__13583\
        );

    \I__2012\ : InMux
    port map (
            O => \N__13678\,
            I => \N__13570\
        );

    \I__2011\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13570\
        );

    \I__2010\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13570\
        );

    \I__2009\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13570\
        );

    \I__2008\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13570\
        );

    \I__2007\ : InMux
    port map (
            O => \N__13669\,
            I => \N__13570\
        );

    \I__2006\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13557\
        );

    \I__2005\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13557\
        );

    \I__2004\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13557\
        );

    \I__2003\ : InMux
    port map (
            O => \N__13665\,
            I => \N__13557\
        );

    \I__2002\ : InMux
    port map (
            O => \N__13664\,
            I => \N__13557\
        );

    \I__2001\ : InMux
    port map (
            O => \N__13663\,
            I => \N__13557\
        );

    \I__2000\ : Span4Mux_h
    port map (
            O => \N__13658\,
            I => \N__13552\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__13649\,
            I => \N__13552\
        );

    \I__1998\ : InMux
    port map (
            O => \N__13648\,
            I => \N__13546\
        );

    \I__1997\ : InMux
    port map (
            O => \N__13647\,
            I => \N__13533\
        );

    \I__1996\ : InMux
    port map (
            O => \N__13646\,
            I => \N__13533\
        );

    \I__1995\ : InMux
    port map (
            O => \N__13645\,
            I => \N__13533\
        );

    \I__1994\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13533\
        );

    \I__1993\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13533\
        );

    \I__1992\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13533\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__13639\,
            I => \N__13530\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__13636\,
            I => \N__13527\
        );

    \I__1989\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13520\
        );

    \I__1988\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13520\
        );

    \I__1987\ : InMux
    port map (
            O => \N__13633\,
            I => \N__13520\
        );

    \I__1986\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13515\
        );

    \I__1985\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13515\
        );

    \I__1984\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13512\
        );

    \I__1983\ : InMux
    port map (
            O => \N__13627\,
            I => \N__13503\
        );

    \I__1982\ : InMux
    port map (
            O => \N__13624\,
            I => \N__13503\
        );

    \I__1981\ : InMux
    port map (
            O => \N__13623\,
            I => \N__13503\
        );

    \I__1980\ : InMux
    port map (
            O => \N__13622\,
            I => \N__13503\
        );

    \I__1979\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13492\
        );

    \I__1978\ : InMux
    port map (
            O => \N__13616\,
            I => \N__13492\
        );

    \I__1977\ : InMux
    port map (
            O => \N__13613\,
            I => \N__13492\
        );

    \I__1976\ : InMux
    port map (
            O => \N__13612\,
            I => \N__13492\
        );

    \I__1975\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13492\
        );

    \I__1974\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13479\
        );

    \I__1973\ : InMux
    port map (
            O => \N__13609\,
            I => \N__13479\
        );

    \I__1972\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13479\
        );

    \I__1971\ : InMux
    port map (
            O => \N__13607\,
            I => \N__13479\
        );

    \I__1970\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13479\
        );

    \I__1969\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13479\
        );

    \I__1968\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13466\
        );

    \I__1967\ : InMux
    port map (
            O => \N__13603\,
            I => \N__13466\
        );

    \I__1966\ : InMux
    port map (
            O => \N__13602\,
            I => \N__13466\
        );

    \I__1965\ : InMux
    port map (
            O => \N__13601\,
            I => \N__13466\
        );

    \I__1964\ : InMux
    port map (
            O => \N__13600\,
            I => \N__13466\
        );

    \I__1963\ : InMux
    port map (
            O => \N__13599\,
            I => \N__13466\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13463\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__13583\,
            I => \N__13454\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__13570\,
            I => \N__13454\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__13557\,
            I => \N__13454\
        );

    \I__1958\ : Span4Mux_h
    port map (
            O => \N__13552\,
            I => \N__13454\
        );

    \I__1957\ : InMux
    port map (
            O => \N__13551\,
            I => \N__13447\
        );

    \I__1956\ : InMux
    port map (
            O => \N__13550\,
            I => \N__13447\
        );

    \I__1955\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13447\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__13546\,
            I => \N__13444\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__13533\,
            I => \N__13439\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__13530\,
            I => \N__13439\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__13527\,
            I => \N__13436\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__13520\,
            I => \N__13415\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__13515\,
            I => \N__13415\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__13512\,
            I => \N__13415\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__13503\,
            I => \N__13415\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__13492\,
            I => \N__13415\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__13479\,
            I => \N__13415\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__13466\,
            I => \N__13415\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__13463\,
            I => \N__13415\
        );

    \I__1942\ : Span4Mux_v
    port map (
            O => \N__13454\,
            I => \N__13415\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__13447\,
            I => \N__13415\
        );

    \I__1940\ : Span4Mux_h
    port map (
            O => \N__13444\,
            I => \N__13412\
        );

    \I__1939\ : Span4Mux_h
    port map (
            O => \N__13439\,
            I => \N__13407\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__13436\,
            I => \N__13407\
        );

    \I__1937\ : Span4Mux_v
    port map (
            O => \N__13415\,
            I => \N__13404\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__13412\,
            I => \tok.n29_adj_787\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__13407\,
            I => \tok.n29_adj_787\
        );

    \I__1934\ : Odrv4
    port map (
            O => \N__13404\,
            I => \tok.n29_adj_787\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__13397\,
            I => \N__13393\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__13396\,
            I => \N__13390\
        );

    \I__1931\ : InMux
    port map (
            O => \N__13393\,
            I => \N__13387\
        );

    \I__1930\ : InMux
    port map (
            O => \N__13390\,
            I => \N__13384\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__13387\,
            I => \N__13381\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__13384\,
            I => \tok.C_stk.tail_22\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__13381\,
            I => \tok.C_stk.tail_22\
        );

    \I__1926\ : CEMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__13373\,
            I => \N__13367\
        );

    \I__1924\ : CEMux
    port map (
            O => \N__13372\,
            I => \N__13364\
        );

    \I__1923\ : CEMux
    port map (
            O => \N__13371\,
            I => \N__13357\
        );

    \I__1922\ : CEMux
    port map (
            O => \N__13370\,
            I => \N__13354\
        );

    \I__1921\ : Span4Mux_v
    port map (
            O => \N__13367\,
            I => \N__13349\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__13364\,
            I => \N__13349\
        );

    \I__1919\ : CEMux
    port map (
            O => \N__13363\,
            I => \N__13346\
        );

    \I__1918\ : CEMux
    port map (
            O => \N__13362\,
            I => \N__13342\
        );

    \I__1917\ : CEMux
    port map (
            O => \N__13361\,
            I => \N__13339\
        );

    \I__1916\ : CEMux
    port map (
            O => \N__13360\,
            I => \N__13336\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__13357\,
            I => \N__13331\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__13354\,
            I => \N__13331\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__13349\,
            I => \N__13325\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__13346\,
            I => \N__13322\
        );

    \I__1911\ : CEMux
    port map (
            O => \N__13345\,
            I => \N__13319\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__13342\,
            I => \N__13316\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__13339\,
            I => \N__13313\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__13336\,
            I => \N__13310\
        );

    \I__1907\ : Span4Mux_v
    port map (
            O => \N__13331\,
            I => \N__13307\
        );

    \I__1906\ : CEMux
    port map (
            O => \N__13330\,
            I => \N__13304\
        );

    \I__1905\ : CEMux
    port map (
            O => \N__13329\,
            I => \N__13301\
        );

    \I__1904\ : CEMux
    port map (
            O => \N__13328\,
            I => \N__13298\
        );

    \I__1903\ : Span4Mux_s2_h
    port map (
            O => \N__13325\,
            I => \N__13295\
        );

    \I__1902\ : Span4Mux_h
    port map (
            O => \N__13322\,
            I => \N__13290\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__13319\,
            I => \N__13290\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__13316\,
            I => \N__13285\
        );

    \I__1899\ : Span4Mux_v
    port map (
            O => \N__13313\,
            I => \N__13285\
        );

    \I__1898\ : Span4Mux_v
    port map (
            O => \N__13310\,
            I => \N__13276\
        );

    \I__1897\ : Span4Mux_v
    port map (
            O => \N__13307\,
            I => \N__13276\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__13304\,
            I => \N__13276\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__13301\,
            I => \N__13276\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__13298\,
            I => \N__13273\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__13295\,
            I => \tok.C_stk_delta_0\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__13290\,
            I => \tok.C_stk_delta_0\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__13285\,
            I => \tok.C_stk_delta_0\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__13276\,
            I => \tok.C_stk_delta_0\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__13273\,
            I => \tok.C_stk_delta_0\
        );

    \I__1888\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13256\
        );

    \I__1887\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13256\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__13256\,
            I => uart_rx_data_4
        );

    \I__1885\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13250\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__13250\,
            I => \N__13247\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__13247\,
            I => \tok.n12_adj_826\
        );

    \I__1882\ : InMux
    port map (
            O => \N__13244\,
            I => \N__13241\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__13241\,
            I => \N__13238\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__13238\,
            I => \N__13234\
        );

    \I__1879\ : InMux
    port map (
            O => \N__13237\,
            I => \N__13231\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__13234\,
            I => \tok.n11_adj_788\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__13231\,
            I => \tok.n11_adj_788\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__13226\,
            I => \N__13223\
        );

    \I__1875\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13220\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__13220\,
            I => \N__13217\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__13217\,
            I => \N__13214\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__13214\,
            I => \N__13211\
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__13211\,
            I => sender_2
        );

    \I__1870\ : InMux
    port map (
            O => \N__13208\,
            I => \N__13205\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__13205\,
            I => \tok.uart.sender_3\
        );

    \I__1868\ : InMux
    port map (
            O => \N__13202\,
            I => \N__13199\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__13199\,
            I => \tok.uart.sender_4\
        );

    \I__1866\ : InMux
    port map (
            O => \N__13196\,
            I => \N__13193\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__13193\,
            I => \tok.uart.sender_5\
        );

    \I__1864\ : InMux
    port map (
            O => \N__13190\,
            I => \N__13187\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__13187\,
            I => \tok.uart.sender_6\
        );

    \I__1862\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13181\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__13181\,
            I => \tok.uart.sender_7\
        );

    \I__1860\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13175\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13172\
        );

    \I__1858\ : Span4Mux_h
    port map (
            O => \N__13172\,
            I => \N__13169\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__13169\,
            I => \tok.n5391\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__13166\,
            I => \tok.n14_adj_688_cascade_\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__13163\,
            I => \tok.n2735_cascade_\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__13160\,
            I => \tok.n1_adj_850_cascade_\
        );

    \I__1853\ : InMux
    port map (
            O => \N__13157\,
            I => \N__13154\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__13154\,
            I => \tok.n26_adj_750\
        );

    \I__1851\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13148\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__13148\,
            I => \tok.n5380\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__13145\,
            I => \N__13142\
        );

    \I__1848\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13139\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__13139\,
            I => \tok.n8_adj_805\
        );

    \I__1846\ : InMux
    port map (
            O => \N__13136\,
            I => \N__13133\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__13133\,
            I => \N__13130\
        );

    \I__1844\ : Span4Mux_v
    port map (
            O => \N__13130\,
            I => \N__13125\
        );

    \I__1843\ : InMux
    port map (
            O => \N__13129\,
            I => \N__13122\
        );

    \I__1842\ : InMux
    port map (
            O => \N__13128\,
            I => \N__13119\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__13125\,
            I => \tok.n11_adj_793\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__13122\,
            I => \tok.n11_adj_793\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__13119\,
            I => \tok.n11_adj_793\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__13112\,
            I => \tok.n5271_cascade_\
        );

    \I__1837\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13106\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__13106\,
            I => \tok.n5318\
        );

    \I__1835\ : InMux
    port map (
            O => \N__13103\,
            I => \N__13100\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__13100\,
            I => \tok.n11_adj_694\
        );

    \I__1833\ : InMux
    port map (
            O => \N__13097\,
            I => \N__13094\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__13094\,
            I => \tok.n15_adj_695\
        );

    \I__1831\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13087\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__13090\,
            I => \N__13083\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__13087\,
            I => \N__13080\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__13086\,
            I => \N__13077\
        );

    \I__1827\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13073\
        );

    \I__1826\ : Span4Mux_s2_h
    port map (
            O => \N__13080\,
            I => \N__13070\
        );

    \I__1825\ : InMux
    port map (
            O => \N__13077\,
            I => \N__13065\
        );

    \I__1824\ : InMux
    port map (
            O => \N__13076\,
            I => \N__13065\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__13073\,
            I => \N__13062\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__13070\,
            I => tc_3
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__13065\,
            I => tc_3
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__13062\,
            I => tc_3
        );

    \I__1819\ : InMux
    port map (
            O => \N__13055\,
            I => \tok.n4756\
        );

    \I__1818\ : InMux
    port map (
            O => \N__13052\,
            I => \tok.n4757\
        );

    \I__1817\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13045\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__13048\,
            I => \N__13042\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__13045\,
            I => \N__13037\
        );

    \I__1814\ : InMux
    port map (
            O => \N__13042\,
            I => \N__13032\
        );

    \I__1813\ : InMux
    port map (
            O => \N__13041\,
            I => \N__13032\
        );

    \I__1812\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13029\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__13037\,
            I => tc_5
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__13032\,
            I => tc_5
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__13029\,
            I => tc_5
        );

    \I__1808\ : InMux
    port map (
            O => \N__13022\,
            I => \N__13019\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__13019\,
            I => \N__13015\
        );

    \I__1806\ : InMux
    port map (
            O => \N__13018\,
            I => \N__13010\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__13015\,
            I => \N__13007\
        );

    \I__1804\ : InMux
    port map (
            O => \N__13014\,
            I => \N__13002\
        );

    \I__1803\ : InMux
    port map (
            O => \N__13013\,
            I => \N__13002\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__13010\,
            I => \tok.tc_plus_1_5\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__13007\,
            I => \tok.tc_plus_1_5\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__13002\,
            I => \tok.tc_plus_1_5\
        );

    \I__1799\ : InMux
    port map (
            O => \N__12995\,
            I => \tok.n4758\
        );

    \I__1798\ : InMux
    port map (
            O => \N__12992\,
            I => \tok.n4759\
        );

    \I__1797\ : InMux
    port map (
            O => \N__12989\,
            I => \N__12984\
        );

    \I__1796\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12978\
        );

    \I__1795\ : InMux
    port map (
            O => \N__12987\,
            I => \N__12978\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__12984\,
            I => \N__12975\
        );

    \I__1793\ : InMux
    port map (
            O => \N__12983\,
            I => \N__12972\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__12978\,
            I => \N__12967\
        );

    \I__1791\ : Span4Mux_h
    port map (
            O => \N__12975\,
            I => \N__12967\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__12972\,
            I => tc_7
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__12967\,
            I => tc_7
        );

    \I__1788\ : InMux
    port map (
            O => \N__12962\,
            I => \tok.n4760\
        );

    \I__1787\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12954\
        );

    \I__1786\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12949\
        );

    \I__1785\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12949\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__12954\,
            I => \N__12943\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__12949\,
            I => \N__12943\
        );

    \I__1782\ : InMux
    port map (
            O => \N__12948\,
            I => \N__12940\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__12943\,
            I => \N__12937\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__12940\,
            I => \tok.tc_plus_1_7\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__12937\,
            I => \tok.tc_plus_1_7\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__12932\,
            I => \N__12929\
        );

    \I__1777\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12920\
        );

    \I__1776\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12907\
        );

    \I__1775\ : InMux
    port map (
            O => \N__12927\,
            I => \N__12907\
        );

    \I__1774\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12907\
        );

    \I__1773\ : InMux
    port map (
            O => \N__12925\,
            I => \N__12907\
        );

    \I__1772\ : InMux
    port map (
            O => \N__12924\,
            I => \N__12907\
        );

    \I__1771\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12907\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__12920\,
            I => \N__12904\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__12907\,
            I => \N__12901\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__12904\,
            I => \N__12898\
        );

    \I__1767\ : Odrv12
    port map (
            O => \N__12901\,
            I => \tok.n9_adj_798\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__12898\,
            I => \tok.n9_adj_798\
        );

    \I__1765\ : InMux
    port map (
            O => \N__12893\,
            I => \N__12890\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__12890\,
            I => \tok.n5293\
        );

    \I__1763\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12881\
        );

    \I__1762\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12881\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__12881\,
            I => \N__12878\
        );

    \I__1760\ : Span4Mux_v
    port map (
            O => \N__12878\,
            I => \N__12875\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__12875\,
            I => \tok.key_rd_7\
        );

    \I__1758\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12866\
        );

    \I__1757\ : InMux
    port map (
            O => \N__12871\,
            I => \N__12866\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__12866\,
            I => \N__12863\
        );

    \I__1755\ : Span4Mux_h
    port map (
            O => \N__12863\,
            I => \N__12860\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__12860\,
            I => \tok.key_rd_2\
        );

    \I__1753\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12854\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__12854\,
            I => \tok.n22_adj_721\
        );

    \I__1751\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12848\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__12848\,
            I => \tok.n23_adj_731\
        );

    \I__1749\ : InMux
    port map (
            O => \N__12845\,
            I => \N__12842\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__12842\,
            I => \tok.n24_adj_651\
        );

    \I__1747\ : InMux
    port map (
            O => \N__12839\,
            I => \N__12833\
        );

    \I__1746\ : InMux
    port map (
            O => \N__12838\,
            I => \N__12833\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__12833\,
            I => \N__12830\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__12830\,
            I => \tok.key_rd_14\
        );

    \I__1743\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12821\
        );

    \I__1742\ : InMux
    port map (
            O => \N__12826\,
            I => \N__12821\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__12821\,
            I => \N__12818\
        );

    \I__1740\ : Span4Mux_h
    port map (
            O => \N__12818\,
            I => \N__12815\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__12815\,
            I => \tok.key_rd_15\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__12812\,
            I => \N__12809\
        );

    \I__1737\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12803\
        );

    \I__1736\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12803\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__12803\,
            I => \N__12800\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__12800\,
            I => \tok.key_rd_9\
        );

    \I__1733\ : InMux
    port map (
            O => \N__12797\,
            I => \N__12791\
        );

    \I__1732\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12791\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__12791\,
            I => \N__12788\
        );

    \I__1730\ : Odrv4
    port map (
            O => \N__12788\,
            I => \tok.key_rd_11\
        );

    \I__1729\ : InMux
    port map (
            O => \N__12785\,
            I => \N__12781\
        );

    \I__1728\ : InMux
    port map (
            O => \N__12784\,
            I => \N__12776\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__12781\,
            I => \N__12773\
        );

    \I__1726\ : InMux
    port map (
            O => \N__12780\,
            I => \N__12768\
        );

    \I__1725\ : InMux
    port map (
            O => \N__12779\,
            I => \N__12768\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__12776\,
            I => \N__12765\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__12773\,
            I => tc_0
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__12768\,
            I => tc_0
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__12765\,
            I => tc_0
        );

    \I__1720\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12753\
        );

    \I__1719\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12749\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__12756\,
            I => \N__12746\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__12753\,
            I => \N__12743\
        );

    \I__1716\ : InMux
    port map (
            O => \N__12752\,
            I => \N__12740\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__12749\,
            I => \N__12737\
        );

    \I__1714\ : InMux
    port map (
            O => \N__12746\,
            I => \N__12734\
        );

    \I__1713\ : Span12Mux_s1_h
    port map (
            O => \N__12743\,
            I => \N__12729\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__12740\,
            I => \N__12729\
        );

    \I__1711\ : Span4Mux_h
    port map (
            O => \N__12737\,
            I => \N__12726\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__12734\,
            I => \tok.tc_plus_1_0\
        );

    \I__1709\ : Odrv12
    port map (
            O => \N__12729\,
            I => \tok.tc_plus_1_0\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__12726\,
            I => \tok.tc_plus_1_0\
        );

    \I__1707\ : InMux
    port map (
            O => \N__12719\,
            I => \bfn_5_8_0_\
        );

    \I__1706\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12713\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__12713\,
            I => \N__12707\
        );

    \I__1704\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12702\
        );

    \I__1703\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12702\
        );

    \I__1702\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12699\
        );

    \I__1701\ : Span4Mux_h
    port map (
            O => \N__12707\,
            I => \N__12696\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__12702\,
            I => \N__12693\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__12699\,
            I => \tok.tc_plus_1_1\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__12696\,
            I => \tok.tc_plus_1_1\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__12693\,
            I => \tok.tc_plus_1_1\
        );

    \I__1696\ : InMux
    port map (
            O => \N__12686\,
            I => \tok.n4754\
        );

    \I__1695\ : InMux
    port map (
            O => \N__12683\,
            I => \N__12677\
        );

    \I__1694\ : InMux
    port map (
            O => \N__12682\,
            I => \N__12674\
        );

    \I__1693\ : InMux
    port map (
            O => \N__12681\,
            I => \N__12669\
        );

    \I__1692\ : InMux
    port map (
            O => \N__12680\,
            I => \N__12669\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__12677\,
            I => \N__12666\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__12674\,
            I => tc_2
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__12669\,
            I => tc_2
        );

    \I__1688\ : Odrv12
    port map (
            O => \N__12666\,
            I => tc_2
        );

    \I__1687\ : InMux
    port map (
            O => \N__12659\,
            I => \N__12655\
        );

    \I__1686\ : InMux
    port map (
            O => \N__12658\,
            I => \N__12651\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__12655\,
            I => \N__12647\
        );

    \I__1684\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12644\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__12651\,
            I => \N__12641\
        );

    \I__1682\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12638\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__12647\,
            I => \N__12633\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__12644\,
            I => \N__12633\
        );

    \I__1679\ : Span4Mux_h
    port map (
            O => \N__12641\,
            I => \N__12630\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__12638\,
            I => \tok.tc_plus_1_2\
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__12633\,
            I => \tok.tc_plus_1_2\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__12630\,
            I => \tok.tc_plus_1_2\
        );

    \I__1675\ : InMux
    port map (
            O => \N__12623\,
            I => \tok.n4755\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__12620\,
            I => \tok.n83_adj_848_cascade_\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__12617\,
            I => \N__12613\
        );

    \I__1672\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12606\
        );

    \I__1671\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12606\
        );

    \I__1670\ : InMux
    port map (
            O => \N__12612\,
            I => \N__12603\
        );

    \I__1669\ : InMux
    port map (
            O => \N__12611\,
            I => \N__12600\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__12606\,
            I => \N__12595\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__12603\,
            I => \N__12595\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__12600\,
            I => \tok.c_stk_r_1\
        );

    \I__1665\ : Odrv12
    port map (
            O => \N__12595\,
            I => \tok.c_stk_r_1\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__12590\,
            I => \tok.ram.n5594_cascade_\
        );

    \I__1663\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12584\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__12584\,
            I => \tok.n5610\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__12581\,
            I => \tok.n3_cascade_\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__12578\,
            I => \tok.n13_cascade_\
        );

    \I__1659\ : InMux
    port map (
            O => \N__12575\,
            I => \N__12572\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__12572\,
            I => \N__12569\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__12569\,
            I => \N__12566\
        );

    \I__1656\ : Span4Mux_s3_h
    port map (
            O => \N__12566\,
            I => \N__12563\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__12563\,
            I => \tok.uart.n5\
        );

    \I__1654\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12554\
        );

    \I__1653\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12554\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__12554\,
            I => \N__12551\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__12551\,
            I => \tok.key_rd_10\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__12548\,
            I => \N__12545\
        );

    \I__1649\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12539\
        );

    \I__1648\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12539\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__12539\,
            I => \N__12536\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__12536\,
            I => \tok.key_rd_12\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__12533\,
            I => \tok.n21_adj_733_cascade_\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__12530\,
            I => \tok.n13_adj_691_cascade_\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__12527\,
            I => \n10_adj_871_cascade_\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__12524\,
            I => \N__12521\
        );

    \I__1641\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12518\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__12518\,
            I => \N__12515\
        );

    \I__1639\ : Span4Mux_h
    port map (
            O => \N__12515\,
            I => \N__12512\
        );

    \I__1638\ : Sp12to4
    port map (
            O => \N__12512\,
            I => \N__12509\
        );

    \I__1637\ : Odrv12
    port map (
            O => \N__12509\,
            I => \tok.tc_6\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__12506\,
            I => \tok.ram.n5605_cascade_\
        );

    \I__1635\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12500\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__12500\,
            I => \tok.n3_adj_690\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__12497\,
            I => \tok.n83_adj_687_cascade_\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__12494\,
            I => \N__12491\
        );

    \I__1631\ : InMux
    port map (
            O => \N__12491\,
            I => \N__12488\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__12488\,
            I => \tok.n5505\
        );

    \I__1629\ : InMux
    port map (
            O => \N__12485\,
            I => \N__12482\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__12482\,
            I => n10_adj_871
        );

    \I__1627\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12476\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__12476\,
            I => \tok.n27_adj_825\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__12473\,
            I => \tok.n5285_cascade_\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__12470\,
            I => \tok.n1_adj_715_cascade_\
        );

    \I__1623\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12455\
        );

    \I__1622\ : InMux
    port map (
            O => \N__12466\,
            I => \N__12455\
        );

    \I__1621\ : InMux
    port map (
            O => \N__12465\,
            I => \N__12455\
        );

    \I__1620\ : InMux
    port map (
            O => \N__12464\,
            I => \N__12455\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__12455\,
            I => \tok.n190\
        );

    \I__1618\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12447\
        );

    \I__1617\ : InMux
    port map (
            O => \N__12451\,
            I => \N__12441\
        );

    \I__1616\ : InMux
    port map (
            O => \N__12450\,
            I => \N__12441\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__12447\,
            I => \N__12438\
        );

    \I__1614\ : InMux
    port map (
            O => \N__12446\,
            I => \N__12435\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__12441\,
            I => \N__12432\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__12438\,
            I => \tok.n890\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__12435\,
            I => \tok.n890\
        );

    \I__1610\ : Odrv4
    port map (
            O => \N__12432\,
            I => \tok.n890\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__12425\,
            I => \tok.n10_adj_763_cascade_\
        );

    \I__1608\ : InMux
    port map (
            O => \N__12422\,
            I => \N__12416\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__12421\,
            I => \N__12412\
        );

    \I__1606\ : InMux
    port map (
            O => \N__12420\,
            I => \N__12409\
        );

    \I__1605\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12406\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__12416\,
            I => \N__12403\
        );

    \I__1603\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12398\
        );

    \I__1602\ : InMux
    port map (
            O => \N__12412\,
            I => \N__12398\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__12409\,
            I => \tok.n5338\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__12406\,
            I => \tok.n5338\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__12403\,
            I => \tok.n5338\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__12398\,
            I => \tok.n5338\
        );

    \I__1597\ : InMux
    port map (
            O => \N__12389\,
            I => \N__12383\
        );

    \I__1596\ : InMux
    port map (
            O => \N__12388\,
            I => \N__12383\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__12383\,
            I => \tok.n5340\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__12380\,
            I => \N__12374\
        );

    \I__1593\ : InMux
    port map (
            O => \N__12379\,
            I => \N__12371\
        );

    \I__1592\ : InMux
    port map (
            O => \N__12378\,
            I => \N__12364\
        );

    \I__1591\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12364\
        );

    \I__1590\ : InMux
    port map (
            O => \N__12374\,
            I => \N__12364\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__12371\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__12364\,
            I => \tok.A_stk_delta_1__N_4\
        );

    \I__1587\ : InMux
    port map (
            O => \N__12359\,
            I => \N__12348\
        );

    \I__1586\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12348\
        );

    \I__1585\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12345\
        );

    \I__1584\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12336\
        );

    \I__1583\ : InMux
    port map (
            O => \N__12355\,
            I => \N__12336\
        );

    \I__1582\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12336\
        );

    \I__1581\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12336\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__12348\,
            I => \tok.n61\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__12345\,
            I => \tok.n61\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__12336\,
            I => \tok.n61\
        );

    \I__1577\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12317\
        );

    \I__1576\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12317\
        );

    \I__1575\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12317\
        );

    \I__1574\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12317\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__12317\,
            I => \tok.n4_adj_813\
        );

    \I__1572\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12310\
        );

    \I__1571\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12307\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__12310\,
            I => tail_97
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__12307\,
            I => tail_97
        );

    \I__1568\ : InMux
    port map (
            O => \N__12302\,
            I => \N__12299\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__12299\,
            I => \N__12295\
        );

    \I__1566\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12292\
        );

    \I__1565\ : Odrv12
    port map (
            O => \N__12295\,
            I => tail_113
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__12292\,
            I => tail_113
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__12287\,
            I => \tok.n27_adj_828_cascade_\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__12284\,
            I => \tok.n27_adj_831_cascade_\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__12281\,
            I => \tok.n27_adj_833_cascade_\
        );

    \I__1560\ : InMux
    port map (
            O => \N__12278\,
            I => \N__12275\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__12275\,
            I => \N__12272\
        );

    \I__1558\ : Odrv12
    port map (
            O => \N__12272\,
            I => \tok.n7_adj_785\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__12269\,
            I => \tok.n14_adj_644_cascade_\
        );

    \I__1556\ : InMux
    port map (
            O => \N__12266\,
            I => \N__12263\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__12263\,
            I => \N__12260\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__12260\,
            I => \tok.table_wr_data_11\
        );

    \I__1553\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12254\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__12254\,
            I => \tok.table_wr_data_10\
        );

    \I__1551\ : InMux
    port map (
            O => \N__12251\,
            I => \N__12248\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__12248\,
            I => \tok.table_wr_data_9\
        );

    \I__1549\ : InMux
    port map (
            O => \N__12245\,
            I => \N__12242\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__12242\,
            I => \tok.table_wr_data_8\
        );

    \I__1547\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12236\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__12236\,
            I => \tok.table_wr_data_0\
        );

    \I__1545\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12230\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__12230\,
            I => \N__12227\
        );

    \I__1543\ : Odrv12
    port map (
            O => \N__12227\,
            I => \tok.n8_adj_790\
        );

    \I__1542\ : InMux
    port map (
            O => \N__12224\,
            I => \N__12221\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__12221\,
            I => \N__12218\
        );

    \I__1540\ : Span12Mux_s4_h
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__12215\,
            I => \tok.table_wr_data_15\
        );

    \I__1538\ : InMux
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__12209\,
            I => \tok.table_wr_data_14\
        );

    \I__1536\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12203\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__12203\,
            I => \N__12200\
        );

    \I__1534\ : Span4Mux_v
    port map (
            O => \N__12200\,
            I => \N__12197\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__12197\,
            I => \tok.table_wr_data_3\
        );

    \I__1532\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12191\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__12191\,
            I => \N__12188\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__12188\,
            I => \N__12185\
        );

    \I__1529\ : Span4Mux_h
    port map (
            O => \N__12185\,
            I => \N__12182\
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__12182\,
            I => \tok.table_wr_data_2\
        );

    \I__1527\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12176\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__12176\,
            I => \N__12173\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__12173\,
            I => \tok.table_wr_data_1\
        );

    \I__1524\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12167\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__12167\,
            I => \N__12164\
        );

    \I__1522\ : Odrv4
    port map (
            O => \N__12164\,
            I => \tok.table_wr_data_5\
        );

    \I__1521\ : InMux
    port map (
            O => \N__12161\,
            I => \N__12158\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__12158\,
            I => \N__12155\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__12155\,
            I => \tok.table_wr_data_7\
        );

    \I__1518\ : InMux
    port map (
            O => \N__12152\,
            I => \N__12149\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__12149\,
            I => \N__12146\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__12146\,
            I => \tok.table_wr_data_13\
        );

    \I__1515\ : InMux
    port map (
            O => \N__12143\,
            I => \N__12140\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__12140\,
            I => \tok.table_wr_data_12\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__12137\,
            I => \tok.ram.n5608_cascade_\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__12134\,
            I => \N__12129\
        );

    \I__1511\ : InMux
    port map (
            O => \N__12133\,
            I => \N__12121\
        );

    \I__1510\ : InMux
    port map (
            O => \N__12132\,
            I => \N__12121\
        );

    \I__1509\ : InMux
    port map (
            O => \N__12129\,
            I => \N__12121\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__12128\,
            I => \N__12118\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__12121\,
            I => \N__12115\
        );

    \I__1506\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12112\
        );

    \I__1505\ : Span4Mux_h
    port map (
            O => \N__12115\,
            I => \N__12109\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__12112\,
            I => \tok.c_stk_r_5\
        );

    \I__1503\ : Odrv4
    port map (
            O => \N__12109\,
            I => \tok.c_stk_r_5\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__12104\,
            I => \tok.n83_adj_678_cascade_\
        );

    \I__1501\ : InMux
    port map (
            O => \N__12101\,
            I => \N__12098\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__12098\,
            I => \tok.n3_adj_683\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__12095\,
            I => \tok.n5483_cascade_\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__12092\,
            I => \tok.n5_adj_684_cascade_\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__12089\,
            I => \n92_adj_868_cascade_\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__12086\,
            I => \N__12083\
        );

    \I__1495\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12080\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__12080\,
            I => \N__12077\
        );

    \I__1493\ : Span4Mux_v
    port map (
            O => \N__12077\,
            I => \N__12074\
        );

    \I__1492\ : Odrv4
    port map (
            O => \N__12074\,
            I => \tok.tc_5\
        );

    \I__1491\ : InMux
    port map (
            O => \N__12071\,
            I => \N__12068\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__12068\,
            I => n92_adj_868
        );

    \I__1489\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12062\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__12062\,
            I => \N__12059\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__12059\,
            I => \tok.table_wr_data_4\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__12056\,
            I => \N__12052\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__12055\,
            I => \N__12049\
        );

    \I__1484\ : InMux
    port map (
            O => \N__12052\,
            I => \N__12041\
        );

    \I__1483\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12041\
        );

    \I__1482\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12041\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__12041\,
            I => \N__12036\
        );

    \I__1480\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12031\
        );

    \I__1479\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12031\
        );

    \I__1478\ : Span4Mux_h
    port map (
            O => \N__12036\,
            I => \N__12028\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__12031\,
            I => \tok.uart.sentbits_0\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__12028\,
            I => \tok.uart.sentbits_0\
        );

    \I__1475\ : InMux
    port map (
            O => \N__12023\,
            I => \N__12014\
        );

    \I__1474\ : InMux
    port map (
            O => \N__12022\,
            I => \N__12014\
        );

    \I__1473\ : InMux
    port map (
            O => \N__12021\,
            I => \N__12014\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__12014\,
            I => \N__12010\
        );

    \I__1471\ : InMux
    port map (
            O => \N__12013\,
            I => \N__12007\
        );

    \I__1470\ : Span4Mux_h
    port map (
            O => \N__12010\,
            I => \N__12004\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__12007\,
            I => \tok.uart.sentbits_1\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__12004\,
            I => \tok.uart.sentbits_1\
        );

    \I__1467\ : CEMux
    port map (
            O => \N__11999\,
            I => \N__11996\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__11996\,
            I => \N__11992\
        );

    \I__1465\ : CEMux
    port map (
            O => \N__11995\,
            I => \N__11989\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__11992\,
            I => \N__11984\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__11989\,
            I => \N__11984\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__11984\,
            I => \tok.uart.n1023\
        );

    \I__1461\ : SRMux
    port map (
            O => \N__11981\,
            I => \N__11977\
        );

    \I__1460\ : SRMux
    port map (
            O => \N__11980\,
            I => \N__11974\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__11977\,
            I => \N__11971\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__11974\,
            I => \N__11968\
        );

    \I__1457\ : Span4Mux_h
    port map (
            O => \N__11971\,
            I => \N__11965\
        );

    \I__1456\ : Span4Mux_h
    port map (
            O => \N__11968\,
            I => \N__11962\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__11965\,
            I => \tok.uart.n1093\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__11962\,
            I => \tok.uart.n1093\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__11957\,
            I => \N__11954\
        );

    \I__1452\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11951\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__11951\,
            I => \N__11948\
        );

    \I__1450\ : Span4Mux_v
    port map (
            O => \N__11948\,
            I => \N__11945\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__11945\,
            I => \tok.n4_adj_707\
        );

    \I__1448\ : InMux
    port map (
            O => \N__11942\,
            I => \N__11939\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__11939\,
            I => \N__11936\
        );

    \I__1446\ : Span4Mux_h
    port map (
            O => \N__11936\,
            I => \N__11933\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__11933\,
            I => \tok.n42\
        );

    \I__1444\ : InMux
    port map (
            O => \N__11930\,
            I => \N__11927\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__11927\,
            I => \tok.n5287\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__11924\,
            I => \tok.n5287_cascade_\
        );

    \I__1441\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11918\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__11918\,
            I => \N__11915\
        );

    \I__1439\ : Span4Mux_h
    port map (
            O => \N__11915\,
            I => \N__11912\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__11912\,
            I => \tok.n7\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__11909\,
            I => \tok.n5312_cascade_\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__11906\,
            I => \tok.n15_adj_817_cascade_\
        );

    \I__1435\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11900\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__11900\,
            I => \tok.n898\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__11897\,
            I => \tok.n898_cascade_\
        );

    \I__1432\ : InMux
    port map (
            O => \N__11894\,
            I => \N__11891\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__11891\,
            I => \tok.uart.n6\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__11888\,
            I => \N__11883\
        );

    \I__1429\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11876\
        );

    \I__1428\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11876\
        );

    \I__1427\ : InMux
    port map (
            O => \N__11883\,
            I => \N__11871\
        );

    \I__1426\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11871\
        );

    \I__1425\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11868\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__11876\,
            I => \tok.n59\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__11871\,
            I => \tok.n59\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__11868\,
            I => \tok.n59\
        );

    \I__1421\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11858\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__11858\,
            I => \tok.depth_3\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__11855\,
            I => \N__11850\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__11854\,
            I => \N__11847\
        );

    \I__1417\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11830\
        );

    \I__1416\ : InMux
    port map (
            O => \N__11850\,
            I => \N__11830\
        );

    \I__1415\ : InMux
    port map (
            O => \N__11847\,
            I => \N__11830\
        );

    \I__1414\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11830\
        );

    \I__1413\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11830\
        );

    \I__1412\ : InMux
    port map (
            O => \N__11844\,
            I => \N__11830\
        );

    \I__1411\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11827\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__11830\,
            I => \tok.n60\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__11827\,
            I => \tok.n60\
        );

    \I__1408\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11819\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__11819\,
            I => \tok.depth_2\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__11816\,
            I => \N__11813\
        );

    \I__1405\ : InMux
    port map (
            O => \N__11813\,
            I => \N__11810\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__11810\,
            I => \N__11807\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__11807\,
            I => \tok.n807\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__11804\,
            I => \n23_cascade_\
        );

    \I__1401\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11795\
        );

    \I__1400\ : InMux
    port map (
            O => \N__11800\,
            I => \N__11795\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__11795\,
            I => \N__11788\
        );

    \I__1398\ : SRMux
    port map (
            O => \N__11794\,
            I => \N__11785\
        );

    \I__1397\ : SRMux
    port map (
            O => \N__11793\,
            I => \N__11782\
        );

    \I__1396\ : InMux
    port map (
            O => \N__11792\,
            I => \N__11777\
        );

    \I__1395\ : InMux
    port map (
            O => \N__11791\,
            I => \N__11777\
        );

    \I__1394\ : Span4Mux_v
    port map (
            O => \N__11788\,
            I => \N__11774\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__11785\,
            I => txtick
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__11782\,
            I => txtick
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__11777\,
            I => txtick
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__11774\,
            I => txtick
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__11765\,
            I => \tok.A_stk_delta_1__N_4_cascade_\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__11762\,
            I => \tok.depth_1_cascade_\
        );

    \I__1387\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__1385\ : Span4Mux_h
    port map (
            O => \N__11753\,
            I => \N__11750\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__11750\,
            I => \tok.n37\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__11747\,
            I => \tok.n2585_cascade_\
        );

    \I__1382\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11738\
        );

    \I__1381\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11738\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__11738\,
            I => \tok.A_stk.tail_33\
        );

    \I__1379\ : InMux
    port map (
            O => \N__11735\,
            I => \N__11729\
        );

    \I__1378\ : InMux
    port map (
            O => \N__11734\,
            I => \N__11729\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__11729\,
            I => \tok.A_stk.tail_49\
        );

    \I__1376\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11720\
        );

    \I__1375\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11720\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__11720\,
            I => \tok.A_stk.tail_65\
        );

    \I__1373\ : InMux
    port map (
            O => \N__11717\,
            I => \N__11711\
        );

    \I__1372\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11711\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__11711\,
            I => \tok.A_stk.tail_81\
        );

    \I__1370\ : InMux
    port map (
            O => \N__11708\,
            I => \N__11702\
        );

    \I__1369\ : InMux
    port map (
            O => \N__11707\,
            I => \N__11702\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__11702\,
            I => \tok.A_stk.tail_1\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__11699\,
            I => \N__11696\
        );

    \I__1366\ : InMux
    port map (
            O => \N__11696\,
            I => \N__11693\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__11693\,
            I => \N__11689\
        );

    \I__1364\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11686\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__11689\,
            I => \tok.tail_62\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__11686\,
            I => \tok.tail_62\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__11681\,
            I => \N__11678\
        );

    \I__1360\ : InMux
    port map (
            O => \N__11678\,
            I => \N__11675\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__11675\,
            I => \tok.C_stk.n5444\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__11672\,
            I => \N__11669\
        );

    \I__1357\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11665\
        );

    \I__1356\ : InMux
    port map (
            O => \N__11668\,
            I => \N__11662\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__11665\,
            I => \tok.tail_54\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__11662\,
            I => \tok.tail_54\
        );

    \I__1353\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11651\
        );

    \I__1352\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11651\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__11651\,
            I => \tok.C_stk.tail_38\
        );

    \I__1350\ : InMux
    port map (
            O => \N__11648\,
            I => \N__11642\
        );

    \I__1349\ : InMux
    port map (
            O => \N__11647\,
            I => \N__11642\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__11642\,
            I => \tok.tail_46\
        );

    \I__1347\ : InMux
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__11636\,
            I => \N__11633\
        );

    \I__1345\ : Span12Mux_s6_v
    port map (
            O => \N__11633\,
            I => \N__11629\
        );

    \I__1344\ : InMux
    port map (
            O => \N__11632\,
            I => \N__11626\
        );

    \I__1343\ : Odrv12
    port map (
            O => \N__11629\,
            I => sender_1
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__11626\,
            I => sender_1
        );

    \I__1341\ : IoInMux
    port map (
            O => \N__11621\,
            I => \N__11618\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__11618\,
            I => \N__11615\
        );

    \I__1339\ : Span4Mux_s1_v
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__11612\,
            I => tx_c
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__1336\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11600\
        );

    \I__1335\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11600\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__11600\,
            I => \tok.A_stk.tail_17\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__11597\,
            I => \N__11594\
        );

    \I__1332\ : InMux
    port map (
            O => \N__11594\,
            I => \N__11591\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__11591\,
            I => \tok.tc_7\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__11588\,
            I => \tok.ram.n5600_cascade_\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__11585\,
            I => \N__11580\
        );

    \I__1328\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11576\
        );

    \I__1327\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11571\
        );

    \I__1326\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11571\
        );

    \I__1325\ : InMux
    port map (
            O => \N__11579\,
            I => \N__11568\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__11576\,
            I => \tok.c_stk_r_7\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__11571\,
            I => \tok.c_stk_r_7\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__11568\,
            I => \tok.c_stk_r_7\
        );

    \I__1321\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11558\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__11558\,
            I => \tok.n5511\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__11555\,
            I => \tok.n3_adj_719_cascade_\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__11552\,
            I => \tok.n5_adj_720_cascade_\
        );

    \I__1317\ : InMux
    port map (
            O => \N__11549\,
            I => \N__11546\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__11546\,
            I => n92_adj_869
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__11543\,
            I => \n92_adj_869_cascade_\
        );

    \I__1314\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11537\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__11537\,
            I => \N__11534\
        );

    \I__1312\ : Odrv4
    port map (
            O => \N__11534\,
            I => \tok.n5507\
        );

    \I__1311\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11527\
        );

    \I__1310\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11524\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__11527\,
            I => \tok.C_stk.tail_4\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__11524\,
            I => \tok.C_stk.tail_4\
        );

    \I__1307\ : InMux
    port map (
            O => \N__11519\,
            I => \N__11516\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__11516\,
            I => n10
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__11513\,
            I => \tok.n36_cascade_\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__11510\,
            I => \tok.n83_adj_842_cascade_\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__11507\,
            I => \tok.ram.n5597_cascade_\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__11504\,
            I => \N__11500\
        );

    \I__1301\ : InMux
    port map (
            O => \N__11503\,
            I => \N__11492\
        );

    \I__1300\ : InMux
    port map (
            O => \N__11500\,
            I => \N__11492\
        );

    \I__1299\ : InMux
    port map (
            O => \N__11499\,
            I => \N__11492\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__11492\,
            I => \N__11488\
        );

    \I__1297\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11485\
        );

    \I__1296\ : Span4Mux_h
    port map (
            O => \N__11488\,
            I => \N__11482\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__11485\,
            I => \tok.c_stk_r_0\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__11482\,
            I => \tok.c_stk_r_0\
        );

    \I__1293\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11474\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__11474\,
            I => \tok.n5583\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__11471\,
            I => \tok.n3_adj_863_cascade_\
        );

    \I__1290\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11465\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__11465\,
            I => \tok.n5_adj_864\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__11462\,
            I => \tok.n83_adj_714_cascade_\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__11459\,
            I => \N__11456\
        );

    \I__1286\ : InMux
    port map (
            O => \N__11456\,
            I => \N__11452\
        );

    \I__1285\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11449\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__11452\,
            I => \tok.tail_29\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__11449\,
            I => \tok.tail_29\
        );

    \I__1282\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11438\
        );

    \I__1281\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11438\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__11438\,
            I => \tok.C_stk.tail_37\
        );

    \I__1279\ : CascadeMux
    port map (
            O => \N__11435\,
            I => \N__11432\
        );

    \I__1278\ : InMux
    port map (
            O => \N__11432\,
            I => \N__11428\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__11431\,
            I => \N__11425\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__11428\,
            I => \N__11422\
        );

    \I__1275\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11419\
        );

    \I__1274\ : Span4Mux_v
    port map (
            O => \N__11422\,
            I => \N__11416\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11413\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__11416\,
            I => \tok.tail_53\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__11413\,
            I => \tok.tail_53\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__11408\,
            I => \N__11404\
        );

    \I__1269\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11401\
        );

    \I__1268\ : InMux
    port map (
            O => \N__11404\,
            I => \N__11398\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__11401\,
            I => \N__11395\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__11398\,
            I => \tok.tail_45\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__11395\,
            I => \tok.tail_45\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__11390\,
            I => \N__11387\
        );

    \I__1263\ : InMux
    port map (
            O => \N__11387\,
            I => \N__11384\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__11384\,
            I => \N__11381\
        );

    \I__1261\ : Span4Mux_v
    port map (
            O => \N__11381\,
            I => \N__11378\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__11378\,
            I => \tok.tc_0\
        );

    \I__1259\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11372\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__11372\,
            I => n92
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__11369\,
            I => \n92_cascade_\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__11366\,
            I => \N__11363\
        );

    \I__1255\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11360\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__11360\,
            I => \N__11357\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__11357\,
            I => \tok.tc_3\
        );

    \I__1252\ : InMux
    port map (
            O => \N__11354\,
            I => \N__11351\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__11351\,
            I => \N__11348\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__11348\,
            I => \tok.n13_adj_646\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__11345\,
            I => \n10_cascade_\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__1247\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__11336\,
            I => \N__11333\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__11333\,
            I => \tok.tc_2\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__11330\,
            I => \tok.n31_adj_795_cascade_\
        );

    \I__1243\ : InMux
    port map (
            O => \N__11327\,
            I => \N__11324\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__11324\,
            I => \tok.n5473\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__11321\,
            I => \tok.C_stk.n5441_cascade_\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__11318\,
            I => \N__11315\
        );

    \I__1239\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11309\
        );

    \I__1238\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11309\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__11309\,
            I => \tok.C_stk.tail_5\
        );

    \I__1236\ : InMux
    port map (
            O => \N__11306\,
            I => \N__11300\
        );

    \I__1235\ : InMux
    port map (
            O => \N__11305\,
            I => \N__11300\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__11300\,
            I => \tok.tail_13\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__11297\,
            I => \N__11293\
        );

    \I__1232\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11290\
        );

    \I__1231\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11287\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__11290\,
            I => \tok.C_stk.tail_21\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__11287\,
            I => \tok.C_stk.tail_21\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__11282\,
            I => \tok.uart.n2_cascade_\
        );

    \I__1227\ : SRMux
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__11276\,
            I => \N__11273\
        );

    \I__1225\ : Span4Mux_s2_h
    port map (
            O => \N__11273\,
            I => \N__11270\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__11270\,
            I => \tok.uart.rxclkcounter_6__N_477\
        );

    \I__1223\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11257\
        );

    \I__1222\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11257\
        );

    \I__1221\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11257\
        );

    \I__1220\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11254\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__11257\,
            I => \N__11251\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__11254\,
            I => \tok.uart.bytephase_2\
        );

    \I__1217\ : Odrv4
    port map (
            O => \N__11251\,
            I => \tok.uart.bytephase_2\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__11246\,
            I => \tok.uart.n13_cascade_\
        );

    \I__1215\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11233\
        );

    \I__1214\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11233\
        );

    \I__1213\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11233\
        );

    \I__1212\ : InMux
    port map (
            O => \N__11240\,
            I => \N__11230\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__11233\,
            I => \N__11227\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__11230\,
            I => \tok.uart.bytephase_4\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__11227\,
            I => \tok.uart.bytephase_4\
        );

    \I__1208\ : SRMux
    port map (
            O => \N__11222\,
            I => \N__11219\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__11219\,
            I => \N__11215\
        );

    \I__1206\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11212\
        );

    \I__1205\ : Span4Mux_s1_v
    port map (
            O => \N__11215\,
            I => \N__11207\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__11212\,
            I => \N__11207\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__11207\,
            I => \bytephase_5__N_510\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__11204\,
            I => \N__11198\
        );

    \I__1201\ : InMux
    port map (
            O => \N__11203\,
            I => \N__11195\
        );

    \I__1200\ : InMux
    port map (
            O => \N__11202\,
            I => \N__11188\
        );

    \I__1199\ : InMux
    port map (
            O => \N__11201\,
            I => \N__11188\
        );

    \I__1198\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11188\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__11195\,
            I => \N__11182\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__11188\,
            I => \N__11182\
        );

    \I__1195\ : InMux
    port map (
            O => \N__11187\,
            I => \N__11179\
        );

    \I__1194\ : Span4Mux_v
    port map (
            O => \N__11182\,
            I => \N__11176\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__11179\,
            I => \tok.uart.bytephase_0\
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__11176\,
            I => \tok.uart.bytephase_0\
        );

    \I__1191\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11165\
        );

    \I__1190\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11165\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__11165\,
            I => \N__11162\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__11162\,
            I => n813
        );

    \I__1187\ : InMux
    port map (
            O => \N__11159\,
            I => \N__11146\
        );

    \I__1186\ : InMux
    port map (
            O => \N__11158\,
            I => \N__11146\
        );

    \I__1185\ : InMux
    port map (
            O => \N__11157\,
            I => \N__11146\
        );

    \I__1184\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11146\
        );

    \I__1183\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11143\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__11146\,
            I => \N__11140\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__11143\,
            I => \tok.uart.bytephase_1\
        );

    \I__1180\ : Odrv12
    port map (
            O => \N__11140\,
            I => \tok.uart.bytephase_1\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__1178\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11127\
        );

    \I__1177\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11123\
        );

    \I__1176\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11120\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__11127\,
            I => \N__11117\
        );

    \I__1174\ : InMux
    port map (
            O => \N__11126\,
            I => \N__11114\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__11123\,
            I => \tok.c_stk_r_2\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__11120\,
            I => \tok.c_stk_r_2\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__11117\,
            I => \tok.c_stk_r_2\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__11114\,
            I => \tok.c_stk_r_2\
        );

    \I__1169\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11102\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__11102\,
            I => \tok.ram.n5585\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__11099\,
            I => \tok.n3_adj_645_cascade_\
        );

    \I__1166\ : InMux
    port map (
            O => \N__11096\,
            I => \N__11093\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__11093\,
            I => \tok.n83\
        );

    \I__1164\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__11087\,
            I => \tok.n5603\
        );

    \I__1162\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11080\
        );

    \I__1161\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11077\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__11080\,
            I => \N__11074\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__11077\,
            I => \tok.uart.txclkcounter_5\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__11074\,
            I => \tok.uart.txclkcounter_5\
        );

    \I__1157\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11065\
        );

    \I__1156\ : InMux
    port map (
            O => \N__11068\,
            I => \N__11062\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__11065\,
            I => \tok.uart.txclkcounter_2\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__11062\,
            I => \tok.uart.txclkcounter_2\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__11057\,
            I => \N__11053\
        );

    \I__1152\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11050\
        );

    \I__1151\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11047\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__11050\,
            I => \tok.uart.txclkcounter_8\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__11047\,
            I => \tok.uart.txclkcounter_8\
        );

    \I__1148\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11038\
        );

    \I__1147\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11035\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__11038\,
            I => \tok.uart.txclkcounter_3\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__11035\,
            I => \tok.uart.txclkcounter_3\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__11030\,
            I => \N__11025\
        );

    \I__1143\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11018\
        );

    \I__1142\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11018\
        );

    \I__1141\ : InMux
    port map (
            O => \N__11025\,
            I => \N__11018\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__11018\,
            I => \tok.uart.sentbits_2\
        );

    \I__1139\ : InMux
    port map (
            O => \N__11015\,
            I => \N__11011\
        );

    \I__1138\ : InMux
    port map (
            O => \N__11014\,
            I => \N__11008\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__11011\,
            I => \tok.uart.txclkcounter_4\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__11008\,
            I => \tok.uart.txclkcounter_4\
        );

    \I__1135\ : InMux
    port map (
            O => \N__11003\,
            I => \N__10999\
        );

    \I__1134\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10996\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__10999\,
            I => \tok.uart.txclkcounter_7\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__10996\,
            I => \tok.uart.txclkcounter_7\
        );

    \I__1131\ : InMux
    port map (
            O => \N__10991\,
            I => \N__10987\
        );

    \I__1130\ : InMux
    port map (
            O => \N__10990\,
            I => \N__10984\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__10987\,
            I => \tok.uart.txclkcounter_6\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__10984\,
            I => \tok.uart.txclkcounter_6\
        );

    \I__1127\ : InMux
    port map (
            O => \N__10979\,
            I => \N__10975\
        );

    \I__1126\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10972\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__10975\,
            I => \tok.uart.txclkcounter_0\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__10972\,
            I => \tok.uart.txclkcounter_0\
        );

    \I__1123\ : InMux
    port map (
            O => \N__10967\,
            I => \N__10963\
        );

    \I__1122\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10960\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__10963\,
            I => \tok.uart.txclkcounter_1\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__10960\,
            I => \tok.uart.txclkcounter_1\
        );

    \I__1119\ : CascadeMux
    port map (
            O => \N__10955\,
            I => \tok.uart.n5418_cascade_\
        );

    \I__1118\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10949\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__10949\,
            I => \tok.uart.n12\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__10946\,
            I => \txtick_cascade_\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__10943\,
            I => \N__10940\
        );

    \I__1114\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10937\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__10937\,
            I => \N__10934\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__10934\,
            I => \N__10930\
        );

    \I__1111\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10927\
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__10930\,
            I => \tok.tail_61\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__10927\,
            I => \tok.tail_61\
        );

    \I__1108\ : InMux
    port map (
            O => \N__10922\,
            I => \tok.uart.n4826\
        );

    \I__1107\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10915\
        );

    \I__1106\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10912\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__10915\,
            I => \tok.uart.rxclkcounter_5\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__10912\,
            I => \tok.uart.rxclkcounter_5\
        );

    \I__1103\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10903\
        );

    \I__1102\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10900\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__10903\,
            I => \tok.uart.rxclkcounter_3\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__10900\,
            I => \tok.uart.rxclkcounter_3\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__10895\,
            I => \N__10891\
        );

    \I__1098\ : InMux
    port map (
            O => \N__10894\,
            I => \N__10888\
        );

    \I__1097\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10885\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__10888\,
            I => \N__10880\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__10885\,
            I => \N__10880\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__10880\,
            I => \tok.uart.rxclkcounter_2\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__10877\,
            I => \n813_cascade_\
        );

    \I__1092\ : CEMux
    port map (
            O => \N__10874\,
            I => \N__10871\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__1090\ : Span4Mux_s2_v
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__10865\,
            I => n971
        );

    \I__1088\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10858\
        );

    \I__1087\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10855\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__10858\,
            I => \tok.uart.rxclkcounter_6\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__10855\,
            I => \tok.uart.rxclkcounter_6\
        );

    \I__1084\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10846\
        );

    \I__1083\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10843\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__10846\,
            I => \tok.uart.rxclkcounter_0\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__10843\,
            I => \tok.uart.rxclkcounter_0\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__10838\,
            I => \N__10834\
        );

    \I__1079\ : InMux
    port map (
            O => \N__10837\,
            I => \N__10831\
        );

    \I__1078\ : InMux
    port map (
            O => \N__10834\,
            I => \N__10828\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__10831\,
            I => \tok.uart.rxclkcounter_4\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__10828\,
            I => \tok.uart.rxclkcounter_4\
        );

    \I__1075\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10819\
        );

    \I__1074\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10816\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__10819\,
            I => \tok.uart.rxclkcounter_1\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__10816\,
            I => \tok.uart.rxclkcounter_1\
        );

    \I__1071\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10808\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__10808\,
            I => \tok.uart.n12_adj_640\
        );

    \I__1069\ : InMux
    port map (
            O => \N__10805\,
            I => \N__10799\
        );

    \I__1068\ : InMux
    port map (
            O => \N__10804\,
            I => \N__10799\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__10799\,
            I => \tok.uart.sentbits_3\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__10796\,
            I => \N__10793\
        );

    \I__1065\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10789\
        );

    \I__1064\ : InMux
    port map (
            O => \N__10792\,
            I => \N__10786\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__10789\,
            I => \N__10783\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__10786\,
            I => \tok.tail_12\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__10783\,
            I => \tok.tail_12\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__10778\,
            I => \N__10774\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__10777\,
            I => \N__10771\
        );

    \I__1058\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10766\
        );

    \I__1057\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10766\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__10766\,
            I => \tok.C_stk.tail_20\
        );

    \I__1055\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10757\
        );

    \I__1054\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10757\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__10757\,
            I => \tok.tail_28\
        );

    \I__1052\ : InMux
    port map (
            O => \N__10754\,
            I => \N__10748\
        );

    \I__1051\ : InMux
    port map (
            O => \N__10753\,
            I => \N__10748\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__10748\,
            I => \tok.C_stk.tail_36\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__10745\,
            I => \N__10741\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__10744\,
            I => \N__10738\
        );

    \I__1047\ : InMux
    port map (
            O => \N__10741\,
            I => \N__10735\
        );

    \I__1046\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10732\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__10735\,
            I => \N__10727\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__10732\,
            I => \N__10727\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__10727\,
            I => \tok.tail_52\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__10724\,
            I => \N__10720\
        );

    \I__1041\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10717\
        );

    \I__1040\ : InMux
    port map (
            O => \N__10720\,
            I => \N__10714\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__10717\,
            I => \N__10711\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__10714\,
            I => \tok.tail_44\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__10711\,
            I => \tok.tail_44\
        );

    \I__1036\ : InMux
    port map (
            O => \N__10706\,
            I => \bfn_2_2_0_\
        );

    \I__1035\ : InMux
    port map (
            O => \N__10703\,
            I => \tok.uart.n4822\
        );

    \I__1034\ : InMux
    port map (
            O => \N__10700\,
            I => \tok.uart.n4823\
        );

    \I__1033\ : InMux
    port map (
            O => \N__10697\,
            I => \tok.uart.n4824\
        );

    \I__1032\ : InMux
    port map (
            O => \N__10694\,
            I => \tok.uart.n4825\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__10691\,
            I => \tok.C_stk.n5435_cascade_\
        );

    \I__1030\ : InMux
    port map (
            O => \N__10688\,
            I => \N__10684\
        );

    \I__1029\ : InMux
    port map (
            O => \N__10687\,
            I => \N__10681\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__10684\,
            I => \tok.C_stk.tail_7\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__10681\,
            I => \tok.C_stk.tail_7\
        );

    \I__1026\ : InMux
    port map (
            O => \N__10676\,
            I => \N__10670\
        );

    \I__1025\ : InMux
    port map (
            O => \N__10675\,
            I => \N__10670\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__10670\,
            I => \tok.tail_15\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__10667\,
            I => \N__10663\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__10666\,
            I => \N__10660\
        );

    \I__1021\ : InMux
    port map (
            O => \N__10663\,
            I => \N__10655\
        );

    \I__1020\ : InMux
    port map (
            O => \N__10660\,
            I => \N__10655\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__10655\,
            I => \tok.C_stk.tail_23\
        );

    \I__1018\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10646\
        );

    \I__1017\ : InMux
    port map (
            O => \N__10651\,
            I => \N__10646\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__10646\,
            I => \tok.tail_31\
        );

    \I__1015\ : InMux
    port map (
            O => \N__10643\,
            I => \N__10637\
        );

    \I__1014\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10637\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__10637\,
            I => \tok.C_stk.tail_39\
        );

    \I__1012\ : CascadeMux
    port map (
            O => \N__10634\,
            I => \N__10630\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__10633\,
            I => \N__10627\
        );

    \I__1010\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10624\
        );

    \I__1009\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10621\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__10624\,
            I => \N__10618\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__10621\,
            I => \tok.tail_55\
        );

    \I__1006\ : Odrv4
    port map (
            O => \N__10618\,
            I => \tok.tail_55\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__10613\,
            I => \N__10610\
        );

    \I__1004\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10606\
        );

    \I__1003\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10603\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__10606\,
            I => \N__10600\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__10603\,
            I => \tok.tail_47\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__10600\,
            I => \tok.tail_47\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__998\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10588\
        );

    \I__997\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10585\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__10588\,
            I => \tok.tail_60\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__10585\,
            I => \tok.tail_60\
        );

    \I__994\ : CascadeMux
    port map (
            O => \N__10580\,
            I => \N__10576\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__10579\,
            I => \N__10573\
        );

    \I__992\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10570\
        );

    \I__991\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10567\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__10570\,
            I => \N__10564\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__10567\,
            I => \tok.tail_51\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__10564\,
            I => \tok.tail_51\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__10559\,
            I => \N__10556\
        );

    \I__986\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10552\
        );

    \I__985\ : InMux
    port map (
            O => \N__10555\,
            I => \N__10549\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__10552\,
            I => \tok.tail_59\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__10549\,
            I => \tok.tail_59\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__981\ : InMux
    port map (
            O => \N__10541\,
            I => \N__10537\
        );

    \I__980\ : InMux
    port map (
            O => \N__10540\,
            I => \N__10534\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__10537\,
            I => \N__10531\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__10534\,
            I => \tok.tail_50\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__10531\,
            I => \tok.tail_50\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__10526\,
            I => \N__10523\
        );

    \I__975\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10519\
        );

    \I__974\ : InMux
    port map (
            O => \N__10522\,
            I => \N__10516\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__10519\,
            I => \tok.tail_58\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__10516\,
            I => \tok.tail_58\
        );

    \I__971\ : InMux
    port map (
            O => \N__10511\,
            I => \N__10507\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__10510\,
            I => \N__10504\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__10507\,
            I => \N__10501\
        );

    \I__968\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10498\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__10501\,
            I => \tok.tail_49\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__10498\,
            I => \tok.tail_49\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__10493\,
            I => \N__10490\
        );

    \I__964\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10487\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__10487\,
            I => \N__10483\
        );

    \I__962\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10480\
        );

    \I__961\ : Odrv4
    port map (
            O => \N__10483\,
            I => \tok.tail_57\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__10480\,
            I => \tok.tail_57\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__10475\,
            I => \N__10471\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__10474\,
            I => \N__10468\
        );

    \I__957\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10465\
        );

    \I__956\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10462\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__10465\,
            I => \N__10459\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__10462\,
            I => \tok.tail_48\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__10459\,
            I => \tok.tail_48\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__951\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10447\
        );

    \I__950\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10444\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__10447\,
            I => \tok.tail_56\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__10444\,
            I => \tok.tail_56\
        );

    \I__947\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10435\
        );

    \I__946\ : InMux
    port map (
            O => \N__10438\,
            I => \N__10432\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__10435\,
            I => \tok.tail_63\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__10432\,
            I => \tok.tail_63\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__10427\,
            I => \N__10423\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__10426\,
            I => \N__10420\
        );

    \I__941\ : InMux
    port map (
            O => \N__10423\,
            I => \N__10415\
        );

    \I__940\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10415\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__10415\,
            I => \tok.C_stk.tail_18\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__10412\,
            I => \N__10408\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__10411\,
            I => \N__10405\
        );

    \I__936\ : InMux
    port map (
            O => \N__10408\,
            I => \N__10400\
        );

    \I__935\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10400\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__10400\,
            I => \tok.tail_26\
        );

    \I__933\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10391\
        );

    \I__932\ : InMux
    port map (
            O => \N__10396\,
            I => \N__10391\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__10391\,
            I => \tok.C_stk.tail_34\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__929\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10381\
        );

    \I__928\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10378\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__10381\,
            I => \tok.tail_43\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__10378\,
            I => \tok.tail_43\
        );

    \I__925\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10369\
        );

    \I__924\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10366\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__10369\,
            I => \tok.tail_42\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__10366\,
            I => \tok.tail_42\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__10361\,
            I => \N__10357\
        );

    \I__920\ : InMux
    port map (
            O => \N__10360\,
            I => \N__10354\
        );

    \I__919\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10351\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__10354\,
            I => \N__10348\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__10351\,
            I => \tok.tail_41\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__10348\,
            I => \tok.tail_41\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__10343\,
            I => \N__10339\
        );

    \I__914\ : InMux
    port map (
            O => \N__10342\,
            I => \N__10336\
        );

    \I__913\ : InMux
    port map (
            O => \N__10339\,
            I => \N__10333\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__10336\,
            I => \N__10330\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__10333\,
            I => \tok.tail_40\
        );

    \I__910\ : Odrv4
    port map (
            O => \N__10330\,
            I => \tok.tail_40\
        );

    \I__909\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10321\
        );

    \I__908\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10318\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__10321\,
            I => \tok.C_stk.tail_1\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__10318\,
            I => \tok.C_stk.tail_1\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__10313\,
            I => \N__10309\
        );

    \I__904\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10304\
        );

    \I__903\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10304\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__10304\,
            I => \tok.tail_9\
        );

    \I__901\ : InMux
    port map (
            O => \N__10301\,
            I => \N__10295\
        );

    \I__900\ : InMux
    port map (
            O => \N__10300\,
            I => \N__10295\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__10295\,
            I => \tok.C_stk.tail_17\
        );

    \I__898\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10286\
        );

    \I__897\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10286\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__10286\,
            I => \tok.tail_25\
        );

    \I__895\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10277\
        );

    \I__894\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10277\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__10277\,
            I => \tok.C_stk.tail_33\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__10274\,
            I => \tok.C_stk.n5450_cascade_\
        );

    \I__891\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10267\
        );

    \I__890\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10264\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__10267\,
            I => \tok.C_stk.tail_2\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__10264\,
            I => \tok.C_stk.tail_2\
        );

    \I__887\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10253\
        );

    \I__886\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10253\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__10253\,
            I => \tok.tail_10\
        );

    \I__884\ : InMux
    port map (
            O => \N__10250\,
            I => \tok.uart.n4816\
        );

    \I__883\ : InMux
    port map (
            O => \N__10247\,
            I => \tok.uart.n4817\
        );

    \I__882\ : InMux
    port map (
            O => \N__10244\,
            I => \tok.uart.n4818\
        );

    \I__881\ : InMux
    port map (
            O => \N__10241\,
            I => \tok.uart.n4819\
        );

    \I__880\ : InMux
    port map (
            O => \N__10238\,
            I => \tok.uart.n4820\
        );

    \I__879\ : InMux
    port map (
            O => \N__10235\,
            I => \bfn_1_5_0_\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__10232\,
            I => \tok.C_stk.n5453_cascade_\
        );

    \I__877\ : InMux
    port map (
            O => \N__10229\,
            I => \tok.uart.n4827\
        );

    \I__876\ : InMux
    port map (
            O => \N__10226\,
            I => \tok.uart.n4828\
        );

    \I__875\ : InMux
    port map (
            O => \N__10223\,
            I => \tok.uart.n4829\
        );

    \I__874\ : InMux
    port map (
            O => \N__10220\,
            I => \tok.uart.n4830\
        );

    \I__873\ : InMux
    port map (
            O => \N__10217\,
            I => \tok.uart.n4831\
        );

    \I__872\ : InMux
    port map (
            O => \N__10214\,
            I => \tok.uart.n4832\
        );

    \I__871\ : InMux
    port map (
            O => \N__10211\,
            I => \bfn_1_4_0_\
        );

    \I__870\ : InMux
    port map (
            O => \N__10208\,
            I => \tok.uart.n4814\
        );

    \I__869\ : InMux
    port map (
            O => \N__10205\,
            I => \tok.uart.n4815\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__10202\,
            I => \tok.C_stk.n5456_cascade_\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__10199\,
            I => \N__10196\
        );

    \I__866\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10190\
        );

    \I__865\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10190\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__10190\,
            I => \tok.C_stk.tail_0\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__10187\,
            I => \N__10183\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__10186\,
            I => \N__10180\
        );

    \I__861\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10175\
        );

    \I__860\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10175\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__10175\,
            I => \tok.tail_8\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__10172\,
            I => \N__10168\
        );

    \I__857\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10165\
        );

    \I__856\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10162\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10157\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__10162\,
            I => \N__10157\
        );

    \I__853\ : Odrv4
    port map (
            O => \N__10157\,
            I => \tok.C_stk.tail_16\
        );

    \I__852\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10148\
        );

    \I__851\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10148\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__10148\,
            I => \tok.tail_24\
        );

    \I__849\ : InMux
    port map (
            O => \N__10145\,
            I => \N__10139\
        );

    \I__848\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10139\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__10139\,
            I => \tok.C_stk.tail_32\
        );

    \I__846\ : InMux
    port map (
            O => \N__10136\,
            I => \bfn_1_3_0_\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__10133\,
            I => \tok.C_stk.n5447_cascade_\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__843\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10121\
        );

    \I__842\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10121\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__10121\,
            I => \tok.C_stk.tail_3\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__10118\,
            I => \N__10114\
        );

    \I__839\ : InMux
    port map (
            O => \N__10117\,
            I => \N__10111\
        );

    \I__838\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10108\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__10111\,
            I => \tok.tail_11\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__10108\,
            I => \tok.tail_11\
        );

    \I__835\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10097\
        );

    \I__834\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10097\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__10097\,
            I => \tok.C_stk.tail_19\
        );

    \I__832\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10088\
        );

    \I__831\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10088\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__10088\,
            I => \tok.tail_27\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__10085\,
            I => \N__10082\
        );

    \I__828\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10078\
        );

    \I__827\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10075\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__10078\,
            I => \tok.C_stk.tail_35\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__10075\,
            I => \tok.C_stk.tail_35\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_4_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.uart.n4821\,
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_2_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_2_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4776\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4783_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4768\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4806\,
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \tok.n4791\,
            carryinitout => \bfn_8_8_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \OSCInst0\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b01"
        )
    port map (
            CLKHFPU => \N__24259\,
            CLKHFEN => \N__24258\,
            CLKHF => clk
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i3_LC_0_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__13601\,
            in1 => \N__14010\,
            in2 => \N__15017\,
            in3 => \N__10117\,
            lcout => \tok.C_stk.tail_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28473\,
            ce => \N__13370\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i5274_3_lut_LC_0_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10126\,
            in1 => \N__14264\,
            in2 => \_gnd_net_\,
            in3 => \N__14981\,
            lcout => OPEN,
            ltout => \tok.C_stk.n5447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i3_LC_0_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__14188\,
            in1 => \N__15543\,
            in2 => \N__10133\,
            in3 => \N__13091\,
            lcout => \tok.c_stk_r_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28473\,
            ce => \N__13370\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i11_LC_0_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14007\,
            in1 => \N__10103\,
            in2 => \N__10130\,
            in3 => \N__13602\,
            lcout => \tok.tail_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28473\,
            ce => \N__13370\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i19_LC_0_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13599\,
            in1 => \N__10094\,
            in2 => \N__10118\,
            in3 => \N__14011\,
            lcout => \tok.C_stk.tail_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28473\,
            ce => \N__13370\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i27_LC_0_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14008\,
            in1 => \N__10102\,
            in2 => \N__10085\,
            in3 => \N__13603\,
            lcout => \tok.tail_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28473\,
            ce => \N__13370\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i35_LC_0_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13600\,
            in1 => \N__10093\,
            in2 => \N__10388\,
            in3 => \N__14012\,
            lcout => \tok.C_stk.tail_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28473\,
            ce => \N__13370\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i43_LC_0_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14009\,
            in1 => \N__10081\,
            in2 => \N__10579\,
            in3 => \N__13604\,
            lcout => \tok.tail_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28473\,
            ce => \N__13370\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i0_LC_0_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__13605\,
            in1 => \N__14020\,
            in2 => \N__10187\,
            in3 => \N__11491\,
            lcout => \tok.C_stk.tail_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28478\,
            ce => \N__13329\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i5283_3_lut_LC_0_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10195\,
            in1 => \N__14251\,
            in2 => \_gnd_net_\,
            in3 => \N__12758\,
            lcout => OPEN,
            ltout => \tok.C_stk.n5456_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i0_LC_0_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__14197\,
            in1 => \N__15544\,
            in2 => \N__10202\,
            in3 => \N__12785\,
            lcout => \tok.c_stk_r_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28478\,
            ce => \N__13329\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i8_LC_0_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14019\,
            in1 => \N__10171\,
            in2 => \N__10199\,
            in3 => \N__13610\,
            lcout => \tok.tail_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28478\,
            ce => \N__13329\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i16_LC_0_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13606\,
            in1 => \N__10154\,
            in2 => \N__10186\,
            in3 => \N__14021\,
            lcout => \tok.C_stk.tail_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28478\,
            ce => \N__13329\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i24_LC_0_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14017\,
            in1 => \N__10145\,
            in2 => \N__10172\,
            in3 => \N__13608\,
            lcout => \tok.tail_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28478\,
            ce => \N__13329\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i32_LC_0_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13607\,
            in1 => \N__10153\,
            in2 => \N__10343\,
            in3 => \N__14022\,
            lcout => \tok.C_stk.tail_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28478\,
            ce => \N__13329\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i40_LC_0_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14018\,
            in1 => \N__10144\,
            in2 => \N__10475\,
            in3 => \N__13609\,
            lcout => \tok.tail_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28478\,
            ce => \N__13329\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i52_LC_0_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14038\,
            in1 => \N__10723\,
            in2 => \N__10595\,
            in3 => \N__13694\,
            lcout => \tok.tail_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28483\,
            ce => \N__13371\,
            sr => \_gnd_net_\
        );

    \tok.uart.rxclkcounter_148__i0_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10850\,
            in2 => \_gnd_net_\,
            in3 => \N__10136\,
            lcout => \tok.uart.rxclkcounter_0\,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \tok.uart.n4827\,
            clk => \N__28466\,
            ce => 'H',
            sr => \N__11279\
        );

    \tok.uart.rxclkcounter_148__i1_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10823\,
            in2 => \_gnd_net_\,
            in3 => \N__10229\,
            lcout => \tok.uart.rxclkcounter_1\,
            ltout => OPEN,
            carryin => \tok.uart.n4827\,
            carryout => \tok.uart.n4828\,
            clk => \N__28466\,
            ce => 'H',
            sr => \N__11279\
        );

    \tok.uart.rxclkcounter_148__i2_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10894\,
            in2 => \_gnd_net_\,
            in3 => \N__10226\,
            lcout => \tok.uart.rxclkcounter_2\,
            ltout => OPEN,
            carryin => \tok.uart.n4828\,
            carryout => \tok.uart.n4829\,
            clk => \N__28466\,
            ce => 'H',
            sr => \N__11279\
        );

    \tok.uart.rxclkcounter_148__i3_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10907\,
            in2 => \_gnd_net_\,
            in3 => \N__10223\,
            lcout => \tok.uart.rxclkcounter_3\,
            ltout => OPEN,
            carryin => \tok.uart.n4829\,
            carryout => \tok.uart.n4830\,
            clk => \N__28466\,
            ce => 'H',
            sr => \N__11279\
        );

    \tok.uart.rxclkcounter_148__i4_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10837\,
            in2 => \_gnd_net_\,
            in3 => \N__10220\,
            lcout => \tok.uart.rxclkcounter_4\,
            ltout => OPEN,
            carryin => \tok.uart.n4830\,
            carryout => \tok.uart.n4831\,
            clk => \N__28466\,
            ce => 'H',
            sr => \N__11279\
        );

    \tok.uart.rxclkcounter_148__i5_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10919\,
            in2 => \_gnd_net_\,
            in3 => \N__10217\,
            lcout => \tok.uart.rxclkcounter_5\,
            ltout => OPEN,
            carryin => \tok.uart.n4831\,
            carryout => \tok.uart.n4832\,
            clk => \N__28466\,
            ce => 'H',
            sr => \N__11279\
        );

    \tok.uart.rxclkcounter_148__i6_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10862\,
            in2 => \_gnd_net_\,
            in3 => \N__10214\,
            lcout => \tok.uart.rxclkcounter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28466\,
            ce => 'H',
            sr => \N__11279\
        );

    \tok.uart.txclkcounter_145__i0_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10979\,
            in2 => \_gnd_net_\,
            in3 => \N__10211\,
            lcout => \tok.uart.txclkcounter_0\,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => \tok.uart.n4814\,
            clk => \N__28468\,
            ce => 'H',
            sr => \N__11793\
        );

    \tok.uart.txclkcounter_145__i1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10967\,
            in2 => \_gnd_net_\,
            in3 => \N__10208\,
            lcout => \tok.uart.txclkcounter_1\,
            ltout => OPEN,
            carryin => \tok.uart.n4814\,
            carryout => \tok.uart.n4815\,
            clk => \N__28468\,
            ce => 'H',
            sr => \N__11793\
        );

    \tok.uart.txclkcounter_145__i2_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11069\,
            in2 => \_gnd_net_\,
            in3 => \N__10205\,
            lcout => \tok.uart.txclkcounter_2\,
            ltout => OPEN,
            carryin => \tok.uart.n4815\,
            carryout => \tok.uart.n4816\,
            clk => \N__28468\,
            ce => 'H',
            sr => \N__11793\
        );

    \tok.uart.txclkcounter_145__i3_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11042\,
            in2 => \_gnd_net_\,
            in3 => \N__10250\,
            lcout => \tok.uart.txclkcounter_3\,
            ltout => OPEN,
            carryin => \tok.uart.n4816\,
            carryout => \tok.uart.n4817\,
            clk => \N__28468\,
            ce => 'H',
            sr => \N__11793\
        );

    \tok.uart.txclkcounter_145__i4_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11015\,
            in2 => \_gnd_net_\,
            in3 => \N__10247\,
            lcout => \tok.uart.txclkcounter_4\,
            ltout => OPEN,
            carryin => \tok.uart.n4817\,
            carryout => \tok.uart.n4818\,
            clk => \N__28468\,
            ce => 'H',
            sr => \N__11793\
        );

    \tok.uart.txclkcounter_145__i5_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11083\,
            in2 => \_gnd_net_\,
            in3 => \N__10244\,
            lcout => \tok.uart.txclkcounter_5\,
            ltout => OPEN,
            carryin => \tok.uart.n4818\,
            carryout => \tok.uart.n4819\,
            clk => \N__28468\,
            ce => 'H',
            sr => \N__11793\
        );

    \tok.uart.txclkcounter_145__i6_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10991\,
            in2 => \_gnd_net_\,
            in3 => \N__10241\,
            lcout => \tok.uart.txclkcounter_6\,
            ltout => OPEN,
            carryin => \tok.uart.n4819\,
            carryout => \tok.uart.n4820\,
            clk => \N__28468\,
            ce => 'H',
            sr => \N__11793\
        );

    \tok.uart.txclkcounter_145__i7_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11003\,
            in2 => \_gnd_net_\,
            in3 => \N__10238\,
            lcout => \tok.uart.txclkcounter_7\,
            ltout => OPEN,
            carryin => \tok.uart.n4820\,
            carryout => \tok.uart.n4821\,
            clk => \N__28468\,
            ce => 'H',
            sr => \N__11793\
        );

    \tok.uart.txclkcounter_145__i8_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11056\,
            in2 => \_gnd_net_\,
            in3 => \N__10235\,
            lcout => \tok.uart.txclkcounter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28470\,
            ce => 'H',
            sr => \N__11794\
        );

    \tok.C_stk.tail_i0_i1_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__10312\,
            in1 => \N__13899\,
            in2 => \N__13692\,
            in3 => \N__12611\,
            lcout => \tok.C_stk.tail_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28474\,
            ce => \N__13345\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i5280_3_lut_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10324\,
            in1 => \N__14269\,
            in2 => \_gnd_net_\,
            in3 => \N__12716\,
            lcout => OPEN,
            ltout => \tok.C_stk.n5453_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i1_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__14164\,
            in1 => \N__15545\,
            in2 => \N__10232\,
            in3 => \N__15731\,
            lcout => \tok.c_stk_r_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28474\,
            ce => \N__13345\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i9_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__13898\,
            in1 => \N__10301\,
            in2 => \N__13690\,
            in3 => \N__10325\,
            lcout => \tok.tail_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28474\,
            ce => \N__13345\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i17_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10292\,
            in1 => \N__13611\,
            in2 => \N__10313\,
            in3 => \N__13900\,
            lcout => \tok.C_stk.tail_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28474\,
            ce => \N__13345\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i25_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__13896\,
            in1 => \N__10300\,
            in2 => \N__13688\,
            in3 => \N__10283\,
            lcout => \tok.tail_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28474\,
            ce => \N__13345\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i33_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10291\,
            in1 => \N__13612\,
            in2 => \N__10361\,
            in3 => \N__13901\,
            lcout => \tok.C_stk.tail_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28474\,
            ce => \N__13345\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i41_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__13897\,
            in1 => \N__10511\,
            in2 => \N__13689\,
            in3 => \N__10282\,
            lcout => \tok.tail_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28474\,
            ce => \N__13345\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i2_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14001\,
            in1 => \N__11131\,
            in2 => \N__13691\,
            in3 => \N__10259\,
            lcout => \tok.C_stk.tail_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28479\,
            ce => \N__13361\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i5277_3_lut_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14260\,
            in1 => \N__10270\,
            in2 => \_gnd_net_\,
            in3 => \N__12659\,
            lcout => OPEN,
            ltout => \tok.C_stk.n5450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i2_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__14187\,
            in1 => \N__15542\,
            in2 => \N__10274\,
            in3 => \N__12682\,
            lcout => \tok.c_stk_r_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28479\,
            ce => \N__13361\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i10_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10271\,
            in1 => \N__13622\,
            in2 => \N__10427\,
            in3 => \N__14003\,
            lcout => \tok.tail_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28479\,
            ce => \N__13361\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i18_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14000\,
            in1 => \N__10258\,
            in2 => \N__10412\,
            in3 => \N__13631\,
            lcout => \tok.C_stk.tail_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28479\,
            ce => \N__13361\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i26_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10397\,
            in1 => \N__13623\,
            in2 => \N__10426\,
            in3 => \N__14004\,
            lcout => \tok.tail_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28479\,
            ce => \N__13361\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i34_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14002\,
            in1 => \N__10373\,
            in2 => \N__10411\,
            in3 => \N__13632\,
            lcout => \tok.C_stk.tail_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28479\,
            ce => \N__13361\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i42_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10396\,
            in1 => \N__13627\,
            in2 => \N__10544\,
            in3 => \N__14005\,
            lcout => \tok.tail_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28479\,
            ce => \N__13361\,
            sr => \_gnd_net_\
        );

    \tok.i2454_2_lut_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13549\,
            in2 => \_gnd_net_\,
            in3 => \N__13902\,
            lcout => \tok.C_stk_delta_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i51_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13904\,
            in1 => \N__10384\,
            in2 => \N__10559\,
            in3 => \N__13634\,
            lcout => \tok.tail_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28484\,
            ce => \N__13328\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i50_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10372\,
            in1 => \N__13551\,
            in2 => \N__10526\,
            in3 => \N__13907\,
            lcout => \tok.tail_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28484\,
            ce => \N__13328\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i49_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13903\,
            in1 => \N__10360\,
            in2 => \N__10493\,
            in3 => \N__13633\,
            lcout => \tok.tail_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28484\,
            ce => \N__13328\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i48_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10342\,
            in1 => \N__13550\,
            in2 => \N__10454\,
            in3 => \N__13906\,
            lcout => \tok.tail_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28484\,
            ce => \N__13328\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i55_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13905\,
            in1 => \N__10439\,
            in2 => \N__10613\,
            in3 => \N__13635\,
            lcout => \tok.tail_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28484\,
            ce => \N__13328\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i60_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__10591\,
            in1 => \N__13683\,
            in2 => \N__10744\,
            in3 => \N__14040\,
            lcout => \tok.tail_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i59_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__13977\,
            in1 => \N__10555\,
            in2 => \N__10580\,
            in3 => \N__13685\,
            lcout => \tok.tail_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i58_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__10522\,
            in1 => \N__13682\,
            in2 => \N__14045\,
            in3 => \N__10540\,
            lcout => \tok.tail_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i57_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__13976\,
            in1 => \N__10486\,
            in2 => \N__10510\,
            in3 => \N__13684\,
            lcout => \tok.tail_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i56_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__10450\,
            in1 => \N__13681\,
            in2 => \N__10474\,
            in3 => \N__14039\,
            lcout => \tok.tail_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i63_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__13979\,
            in1 => \N__10438\,
            in2 => \N__10633\,
            in3 => \N__13687\,
            lcout => \tok.tail_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.i547_4_lut_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__13244\,
            in1 => \N__17498\,
            in2 => \N__14195\,
            in3 => \N__13136\,
            lcout => \tok.C_stk.n602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i61_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__13978\,
            in1 => \N__10933\,
            in2 => \N__11435\,
            in3 => \N__13686\,
            lcout => \tok.tail_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i7_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14034\,
            in1 => \N__10676\,
            in2 => \N__13713\,
            in3 => \N__11584\,
            lcout => \tok.C_stk.tail_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28496\,
            ce => \N__13330\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i5262_3_lut_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14256\,
            in1 => \N__10687\,
            in2 => \_gnd_net_\,
            in3 => \N__12959\,
            lcout => OPEN,
            ltout => \tok.C_stk.n5435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i7_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14196\,
            in1 => \N__12983\,
            in2 => \N__10691\,
            in3 => \N__15527\,
            lcout => \tok.c_stk_r_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28496\,
            ce => \N__13330\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i15_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10688\,
            in1 => \N__13669\,
            in2 => \N__10667\,
            in3 => \N__14035\,
            lcout => \tok.tail_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28496\,
            ce => \N__13330\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i23_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14032\,
            in1 => \N__10652\,
            in2 => \N__13711\,
            in3 => \N__10675\,
            lcout => \tok.C_stk.tail_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28496\,
            ce => \N__13330\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i31_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__10643\,
            in1 => \N__13670\,
            in2 => \N__10666\,
            in3 => \N__14036\,
            lcout => \tok.tail_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28496\,
            ce => \N__13330\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i39_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14033\,
            in1 => \N__10609\,
            in2 => \N__13712\,
            in3 => \N__10651\,
            lcout => \tok.C_stk.tail_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28496\,
            ce => \N__13330\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i47_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10642\,
            in1 => \N__13671\,
            in2 => \N__10634\,
            in3 => \N__14037\,
            lcout => \tok.tail_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28496\,
            ce => \N__13330\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i4_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__13665\,
            in1 => \N__14029\,
            in2 => \N__16071\,
            in3 => \N__10792\,
            lcout => \tok.C_stk.tail_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28501\,
            ce => \N__13360\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i12_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14026\,
            in1 => \N__11531\,
            in2 => \N__10778\,
            in3 => \N__13666\,
            lcout => \tok.tail_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28501\,
            ce => \N__13360\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i20_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13663\,
            in1 => \N__10763\,
            in2 => \N__10796\,
            in3 => \N__14030\,
            lcout => \tok.C_stk.tail_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28501\,
            ce => \N__13360\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i28_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14027\,
            in1 => \N__10754\,
            in2 => \N__10777\,
            in3 => \N__13667\,
            lcout => \tok.tail_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28501\,
            ce => \N__13360\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i36_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13664\,
            in1 => \N__10762\,
            in2 => \N__10724\,
            in3 => \N__14031\,
            lcout => \tok.C_stk.tail_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28501\,
            ce => \N__13360\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i44_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14028\,
            in1 => \N__10753\,
            in2 => \N__10745\,
            in3 => \N__13668\,
            lcout => \tok.tail_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28501\,
            ce => \N__13360\,
            sr => \_gnd_net_\
        );

    \tok.uart.bytephase__i0_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11187\,
            in2 => \_gnd_net_\,
            in3 => \N__10706\,
            lcout => \tok.uart.bytephase_0\,
            ltout => OPEN,
            carryin => \bfn_2_2_0_\,
            carryout => \tok.uart.n4822\,
            clk => \N__28467\,
            ce => \N__10874\,
            sr => \N__11222\
        );

    \tok.uart.bytephase__i1_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11155\,
            in2 => \_gnd_net_\,
            in3 => \N__10703\,
            lcout => \tok.uart.bytephase_1\,
            ltout => OPEN,
            carryin => \tok.uart.n4822\,
            carryout => \tok.uart.n4823\,
            clk => \N__28467\,
            ce => \N__10874\,
            sr => \N__11222\
        );

    \tok.uart.bytephase__i2_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11264\,
            in2 => \_gnd_net_\,
            in3 => \N__10700\,
            lcout => \tok.uart.bytephase_2\,
            ltout => OPEN,
            carryin => \tok.uart.n4823\,
            carryout => \tok.uart.n4824\,
            clk => \N__28467\,
            ce => \N__10874\,
            sr => \N__11222\
        );

    \tok.uart.bytephase__i3_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17067\,
            in2 => \_gnd_net_\,
            in3 => \N__10697\,
            lcout => \tok.uart.bytephase_3\,
            ltout => OPEN,
            carryin => \tok.uart.n4824\,
            carryout => \tok.uart.n4825\,
            clk => \N__28467\,
            ce => \N__10874\,
            sr => \N__11222\
        );

    \tok.uart.bytephase__i4_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11240\,
            in2 => \_gnd_net_\,
            in3 => \N__10694\,
            lcout => \tok.uart.bytephase_4\,
            ltout => OPEN,
            carryin => \tok.uart.n4825\,
            carryout => \tok.uart.n4826\,
            clk => \N__28467\,
            ce => \N__10874\,
            sr => \N__11222\
        );

    \tok.uart.bytephase__i5_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17097\,
            in2 => \_gnd_net_\,
            in3 => \N__10922\,
            lcout => \tok.uart.bytephase_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28467\,
            ce => \N__10874\,
            sr => \N__11222\
        );

    \tok.uart.i6_4_lut_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__10918\,
            in1 => \N__10906\,
            in2 => \N__10895\,
            in3 => \N__10811\,
            lcout => n813,
            ltout => \n813_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10877\,
            in3 => \N__11218\,
            lcout => n971,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i10_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001010100"
        )
    port map (
            in0 => \N__14374\,
            in1 => \N__11791\,
            in2 => \N__14401\,
            in3 => \N__22326\,
            lcout => sender_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i2_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__11792\,
            in1 => \N__11632\,
            in2 => \N__13226\,
            in3 => \N__14373\,
            lcout => sender_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i127_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__16516\,
            in1 => \N__26057\,
            in2 => \N__17186\,
            in3 => \N__26581\,
            lcout => tail_127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i5_4_lut_adj_27_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__10861\,
            in1 => \N__10849\,
            in2 => \N__10838\,
            in3 => \N__10822\,
            lcout => \tok.uart.n12_adj_640\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i2_4_lut_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__10804\,
            in1 => \N__12048\,
            in2 => \N__11030\,
            in3 => \N__12021\,
            lcout => \tok.uart_tx_busy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sentbits_147__i3_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12023\,
            in1 => \N__11029\,
            in2 => \N__12056\,
            in3 => \N__10805\,
            lcout => \tok.uart.sentbits_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28471\,
            ce => \N__11999\,
            sr => \N__11981\
        );

    \tok.uart.i5_4_lut_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__11084\,
            in1 => \N__11068\,
            in2 => \N__11057\,
            in3 => \N__11041\,
            lcout => \tok.uart.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sentbits_147__i2_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__12022\,
            in1 => \_gnd_net_\,
            in2 => \N__12055\,
            in3 => \N__11028\,
            lcout => \tok.uart.sentbits_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28471\,
            ce => \N__11999\,
            sr => \N__11981\
        );

    \tok.uart.i5246_3_lut_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11014\,
            in1 => \N__11002\,
            in2 => \_gnd_net_\,
            in3 => \N__10990\,
            lcout => OPEN,
            ltout => \tok.uart.n5418_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i5618_4_lut_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10978\,
            in1 => \N__10966\,
            in2 => \N__10955\,
            in3 => \N__10952\,
            lcout => txtick,
            ltout => \txtick_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i5612_2_lut_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10946\,
            in3 => \N__14365\,
            lcout => \tok.uart.n1017\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i53_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__11407\,
            in1 => \N__13648\,
            in2 => \N__10943\,
            in3 => \N__14006\,
            lcout => \tok.tail_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28475\,
            ce => \N__13363\,
            sr => \_gnd_net_\
        );

    \tok.ram.i5523_4_lut_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__15963\,
            in1 => \N__12658\,
            in2 => \N__11135\,
            in3 => \N__19903\,
            lcout => \tok.ram.n5585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_4_lut_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__11156\,
            in1 => \N__11265\,
            in2 => \N__11204\,
            in3 => \N__11241\,
            lcout => \tok.uart.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i2_2_lut_3_lut_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__11266\,
            in1 => \N__11159\,
            in2 => \_gnd_net_\,
            in3 => \N__11202\,
            lcout => OPEN,
            ltout => \tok.uart.n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rxrst_I_0_4_lut_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011101"
        )
    port map (
            in0 => \N__11171\,
            in1 => \N__17123\,
            in2 => \N__11282\,
            in3 => \N__11243\,
            lcout => \tok.uart.rxclkcounter_6__N_477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i24_3_lut_4_lut_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010100000"
        )
    port map (
            in0 => \N__17101\,
            in1 => \N__17159\,
            in2 => \N__17078\,
            in3 => \N__11157\,
            lcout => OPEN,
            ltout => \tok.uart.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_3_lut_4_lut_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11201\,
            in1 => \N__11267\,
            in2 => \N__11246\,
            in3 => \N__11242\,
            lcout => \bytephase_5__N_510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i2_3_lut_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__11203\,
            in1 => \N__11170\,
            in2 => \_gnd_net_\,
            in3 => \N__11158\,
            lcout => n4858,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__11126\,
            in1 => \N__18340\,
            in2 => \N__17719\,
            in3 => \N__20292\,
            lcout => \tok.n83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6_4_lut_adj_20_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__11130\,
            in1 => \N__11105\,
            in2 => \N__15889\,
            in3 => \N__29997\,
            lcout => OPEN,
            ltout => \tok.n3_adj_645_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_29_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__19236\,
            in1 => \N__11090\,
            in2 => \N__11099\,
            in3 => \N__20295\,
            lcout => \tok.n13_adj_646\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5540_2_lut_3_lut_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11096\,
            in1 => \N__19056\,
            in2 => \_gnd_net_\,
            in3 => \N__29996\,
            lcout => \tok.n5603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111101111111"
        )
    port map (
            in0 => \N__29995\,
            in1 => \N__18341\,
            in2 => \N__19255\,
            in3 => \N__20294\,
            lcout => \tok.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i59_3_lut_adj_127_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__18339\,
            in1 => \N__19055\,
            in2 => \_gnd_net_\,
            in3 => \N__29994\,
            lcout => OPEN,
            ltout => \tok.n31_adj_795_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i58_4_lut_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__19232\,
            in1 => \N__11327\,
            in2 => \N__11330\,
            in3 => \N__20293\,
            lcout => \tok.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5450_4_lut_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010000000"
        )
    port map (
            in0 => \N__20291\,
            in1 => \N__19054\,
            in2 => \N__18359\,
            in3 => \N__29993\,
            lcout => \tok.n5473\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i5_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__13644\,
            in1 => \N__13997\,
            in2 => \N__12128\,
            in3 => \N__11306\,
            lcout => \tok.C_stk.tail_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28485\,
            ce => \N__13372\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i5268_3_lut_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11314\,
            in1 => \N__14265\,
            in2 => \_gnd_net_\,
            in3 => \N__13022\,
            lcout => OPEN,
            ltout => \tok.C_stk.n5441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i5_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__14186\,
            in1 => \N__15528\,
            in2 => \N__11321\,
            in3 => \N__13049\,
            lcout => \tok.c_stk_r_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28485\,
            ce => \N__13372\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i13_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13994\,
            in1 => \N__11296\,
            in2 => \N__11318\,
            in3 => \N__13645\,
            lcout => \tok.tail_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28485\,
            ce => \N__13372\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i21_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13642\,
            in1 => \N__11305\,
            in2 => \N__11459\,
            in3 => \N__13998\,
            lcout => \tok.C_stk.tail_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28485\,
            ce => \N__13372\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i29_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__13995\,
            in1 => \N__11444\,
            in2 => \N__11297\,
            in3 => \N__13646\,
            lcout => \tok.tail_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28485\,
            ce => \N__13372\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i37_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13643\,
            in1 => \N__11455\,
            in2 => \N__11408\,
            in3 => \N__13999\,
            lcout => \tok.C_stk.tail_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28485\,
            ce => \N__13372\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i45_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__13996\,
            in1 => \N__11443\,
            in2 => \N__11431\,
            in3 => \N__13647\,
            lcout => \tok.tail_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28485\,
            ce => \N__13372\,
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_89_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11375\,
            in1 => \N__16196\,
            in2 => \_gnd_net_\,
            in3 => \N__12779\,
            lcout => \tok.tc_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_197_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__16310\,
            in1 => \N__12752\,
            in2 => \N__16382\,
            in3 => \N__11468\,
            lcout => n92,
            ltout => \n92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i0_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16197\,
            in2 => \N__11369\,
            in3 => \N__12780\,
            lcout => tc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28489\,
            ce => 'H',
            sr => \N__28238\
        );

    \tok.tc_i3_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__16201\,
            in1 => \N__14945\,
            in2 => \N__13086\,
            in3 => \_gnd_net_\,
            lcout => tc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28489\,
            ce => 'H',
            sr => \N__28238\
        );

    \tok.i26_3_lut_adj_86_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14944\,
            in1 => \N__13076\,
            in2 => \_gnd_net_\,
            in3 => \N__16194\,
            lcout => \tok.tc_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_32_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__16311\,
            in1 => \N__12654\,
            in2 => \N__16383\,
            in3 => \N__11354\,
            lcout => n10,
            ltout => \n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_87_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16195\,
            in2 => \N__11345\,
            in3 => \N__12680\,
            lcout => \tok.tc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i2_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__12681\,
            in1 => \_gnd_net_\,
            in2 => \N__16205\,
            in3 => \N__11519\,
            lcout => tc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28489\,
            ce => 'H',
            sr => \N__28238\
        );

    \tok.i57_3_lut_3_lut_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__19017\,
            in1 => \N__18293\,
            in2 => \_gnd_net_\,
            in3 => \N__29942\,
            lcout => OPEN,
            ltout => \tok.n36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i59_4_lut_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__20265\,
            in1 => \N__11540\,
            in2 => \N__11513\,
            in3 => \N__19198\,
            lcout => \tok.n42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_194_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__11499\,
            in1 => \N__18294\,
            in2 => \N__17560\,
            in3 => \N__20266\,
            lcout => OPEN,
            ltout => \tok.n83_adj_842_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5522_2_lut_3_lut_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__29943\,
            in1 => \_gnd_net_\,
            in2 => \N__11510\,
            in3 => \N__19018\,
            lcout => \tok.n5583\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5531_4_lut_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__15961\,
            in1 => \N__12757\,
            in2 => \N__11504\,
            in3 => \N__19896\,
            lcout => OPEN,
            ltout => \tok.ram.n5597_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6_4_lut_adj_26_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__29944\,
            in1 => \N__15875\,
            in2 => \N__11507\,
            in3 => \N__11503\,
            lcout => OPEN,
            ltout => \tok.n3_adj_863_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i18_4_lut_adj_196_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__19199\,
            in1 => \N__11477\,
            in2 => \N__11471\,
            in3 => \N__20267\,
            lcout => \tok.n5_adj_864\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_68_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__11579\,
            in1 => \N__18295\,
            in2 => \N__19300\,
            in3 => \N__20268\,
            lcout => OPEN,
            ltout => \tok.n83_adj_714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5495_2_lut_3_lut_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18924\,
            in2 => \N__11462\,
            in3 => \N__29945\,
            lcout => \tok.n5511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12987\,
            in1 => \N__16202\,
            in2 => \_gnd_net_\,
            in3 => \N__11549\,
            lcout => \tok.tc_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5535_4_lut_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__15962\,
            in1 => \N__19902\,
            in2 => \N__11585\,
            in3 => \N__12957\,
            lcout => OPEN,
            ltout => \tok.ram.n5600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6_4_lut_adj_25_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__29946\,
            in1 => \N__15890\,
            in2 => \N__11588\,
            in3 => \N__11583\,
            lcout => OPEN,
            ltout => \tok.n3_adj_719_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i18_4_lut_adj_70_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__20269\,
            in1 => \N__11561\,
            in2 => \N__11555\,
            in3 => \N__19166\,
            lcout => OPEN,
            ltout => \tok.n5_adj_720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_77_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__12958\,
            in1 => \N__16390\,
            in2 => \N__11552\,
            in3 => \N__16312\,
            lcout => n92_adj_869,
            ltout => \n92_adj_869_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i7_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__16203\,
            in1 => \_gnd_net_\,
            in2 => \N__11543\,
            in3 => \N__12988\,
            lcout => tc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28502\,
            ce => 'H',
            sr => \N__28226\
        );

    \tok.i5492_3_lut_4_lut_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__18214\,
            in1 => \N__20145\,
            in2 => \N__18963\,
            in3 => \N__29878\,
            lcout => \tok.n5507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i62_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__11692\,
            in1 => \N__13693\,
            in2 => \N__11672\,
            in3 => \N__14044\,
            lcout => \tok.tail_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.i5271_3_lut_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11530\,
            in1 => \N__14255\,
            in2 => \_gnd_net_\,
            in3 => \N__16253\,
            lcout => \tok.C_stk.n5444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i30_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11657\,
            in1 => \N__13695\,
            in2 => \N__13397\,
            in3 => \N__14015\,
            lcout => \tok.tail_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28514\,
            ce => \N__13376\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i38_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14013\,
            in1 => \N__11648\,
            in2 => \N__13714\,
            in3 => \N__13732\,
            lcout => \tok.C_stk.tail_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28514\,
            ce => \N__13376\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i54_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__11647\,
            in1 => \N__13696\,
            in2 => \N__11699\,
            in3 => \N__14016\,
            lcout => \tok.tail_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28514\,
            ce => \N__13376\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i4_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__14204\,
            in1 => \N__15535\,
            in2 => \N__11681\,
            in3 => \N__16105\,
            lcout => \tok.c_stk_r_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28514\,
            ce => \N__13376\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i46_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14014\,
            in1 => \N__11668\,
            in2 => \N__13715\,
            in3 => \N__11656\,
            lcout => \tok.tail_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28514\,
            ce => \N__13376\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i1_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11639\,
            lcout => tx_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28522\,
            ce => \N__14293\,
            sr => \N__14381\
        );

    \tok.A_stk.tail_i0_i17_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11744\,
            in1 => \N__11708\,
            in2 => \_gnd_net_\,
            in3 => \N__26553\,
            lcout => \tok.A_stk.tail_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28472\,
            ce => \N__26072\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i1_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26554\,
            in1 => \_gnd_net_\,
            in2 => \N__11609\,
            in3 => \N__23980\,
            lcout => \tok.A_stk.tail_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28472\,
            ce => \N__26072\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i33_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11735\,
            in1 => \N__11605\,
            in2 => \_gnd_net_\,
            in3 => \N__26555\,
            lcout => \tok.A_stk.tail_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28472\,
            ce => \N__26072\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i49_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26556\,
            in1 => \N__11743\,
            in2 => \_gnd_net_\,
            in3 => \N__11726\,
            lcout => \tok.A_stk.tail_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28472\,
            ce => \N__26072\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i65_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11734\,
            in1 => \N__11717\,
            in2 => \_gnd_net_\,
            in3 => \N__26557\,
            lcout => \tok.A_stk.tail_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28472\,
            ce => \N__26072\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i81_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26558\,
            in1 => \N__12313\,
            in2 => \_gnd_net_\,
            in3 => \N__11725\,
            lcout => \tok.A_stk.tail_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28472\,
            ce => \N__26072\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i97_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12302\,
            in1 => \N__11716\,
            in2 => \_gnd_net_\,
            in3 => \N__26559\,
            lcout => tail_97,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28472\,
            ce => \N__26072\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i1_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11707\,
            in1 => \N__25467\,
            in2 => \_gnd_net_\,
            in3 => \N__21142\,
            lcout => \tok.S_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28472\,
            ce => \N__26072\,
            sr => \_gnd_net_\
        );

    \tok.depth_i1_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001011010101010"
        )
    port map (
            in0 => \N__12359\,
            in1 => \N__12379\,
            in2 => \N__16497\,
            in3 => \N__16435\,
            lcout => \tok.n61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28476\,
            ce => 'H',
            sr => \N__28235\
        );

    \tok.i1_2_lut_3_lut_adj_156_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__12355\,
            in1 => \_gnd_net_\,
            in2 => \N__16493\,
            in3 => \N__18833\,
            lcout => \tok.n4_adj_707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_4_lut_adj_167_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__12358\,
            in1 => \N__22150\,
            in2 => \N__18058\,
            in3 => \N__16480\,
            lcout => \tok.n807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_i0_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16488\,
            lcout => \tok.n62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28476\,
            ce => 'H',
            sr => \N__28235\
        );

    \tok.i1_2_lut_adj_147_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16476\,
            in2 => \_gnd_net_\,
            in3 => \N__12354\,
            lcout => \tok.n890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_4_lut_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12353\,
            in1 => \N__11881\,
            in2 => \N__16492\,
            in3 => \N__11843\,
            lcout => \tok.A_stk_delta_1__N_4\,
            ltout => \tok.A_stk_delta_1__N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_4_lut_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011011001100"
        )
    port map (
            in0 => \N__16484\,
            in1 => \N__12356\,
            in2 => \N__11765\,
            in3 => \N__16433\,
            lcout => OPEN,
            ltout => \tok.depth_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5236_3_lut_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11861\,
            in2 => \N__11762\,
            in3 => \N__11822\,
            lcout => \tok.n5408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_4_lut_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__12419\,
            in1 => \N__12451\,
            in2 => \N__19334\,
            in3 => \N__18053\,
            lcout => \tok.n820\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5173_2_lut_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11882\,
            in2 => \_gnd_net_\,
            in3 => \N__11844\,
            lcout => \tok.n5338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2525_2_lut_3_lut_4_lut_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__11845\,
            in1 => \N__12450\,
            in2 => \N__11888\,
            in3 => \N__16944\,
            lcout => \tok.n2585\,
            ltout => \tok.n2585_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_4_lut_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__18054\,
            in1 => \N__11759\,
            in2 => \N__11747\,
            in3 => \N__19333\,
            lcout => \tok.n29_adj_787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.depth_i3_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101101100100100"
        )
    port map (
            in0 => \N__12329\,
            in1 => \N__12467\,
            in2 => \N__11855\,
            in3 => \N__11887\,
            lcout => \tok.n59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28480\,
            ce => 'H',
            sr => \N__28236\
        );

    \tok.depth_i2_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12466\,
            in1 => \N__11853\,
            in2 => \_gnd_net_\,
            in3 => \N__12328\,
            lcout => \tok.n60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28480\,
            ce => 'H',
            sr => \N__28236\
        );

    \tok.i2_4_lut_adj_139_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101100100100"
        )
    port map (
            in0 => \N__12327\,
            in1 => \N__12465\,
            in2 => \N__11854\,
            in3 => \N__11886\,
            lcout => \tok.depth_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_134_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12464\,
            in1 => \N__11846\,
            in2 => \_gnd_net_\,
            in3 => \N__12326\,
            lcout => \tok.depth_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_48_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12420\,
            in1 => \N__11903\,
            in2 => \N__11816\,
            in3 => \N__18306\,
            lcout => \tok.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_220_i9_2_lut_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__18305\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20228\,
            lcout => \tok.n9_adj_766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i5605_4_lut_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11894\,
            in1 => \N__18051\,
            in2 => \N__17812\,
            in3 => \N__18307\,
            lcout => n23,
            ltout => \n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i5610_2_lut_3_lut_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__11800\,
            in1 => \_gnd_net_\,
            in2 => \N__11804\,
            in3 => \N__17807\,
            lcout => \tok.uart.n1093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_119_i9_2_lut_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__20227\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18304\,
            lcout => \tok.n9_adj_798\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_3_lut_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__11801\,
            in1 => \N__17808\,
            in2 => \_gnd_net_\,
            in3 => \N__14332\,
            lcout => \tok.uart.n1023\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sentbits_147__i0_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12039\,
            lcout => \tok.uart.sentbits_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28486\,
            ce => \N__11995\,
            sr => \N__11980\
        );

    \tok.uart.sentbits_147__i1_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12040\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12013\,
            lcout => \tok.uart.sentbits_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28486\,
            ce => \N__11995\,
            sr => \N__11980\
        );

    \tok.i2_4_lut_adj_64_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__11930\,
            in1 => \N__12422\,
            in2 => \N__11957\,
            in3 => \N__11942\,
            lcout => \tok.n5298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_119_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22134\,
            in2 => \_gnd_net_\,
            in3 => \N__18026\,
            lcout => \tok.n5287\,
            ltout => \tok.n5287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_122_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__12233\,
            in1 => \N__12278\,
            in2 => \N__11924\,
            in3 => \N__16584\,
            lcout => \tok.n241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5149_2_lut_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18835\,
            in2 => \_gnd_net_\,
            in3 => \N__18027\,
            lcout => OPEN,
            ltout => \tok.n5312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_124_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__19060\,
            in1 => \N__11921\,
            in2 => \N__11909\,
            in3 => \N__14930\,
            lcout => \tok.n2515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_143_i15_2_lut_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19059\,
            in2 => \_gnd_net_\,
            in3 => \N__18834\,
            lcout => OPEN,
            ltout => \tok.n15_adj_817_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i3_4_lut_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19239\,
            in1 => \N__20232\,
            in2 => \N__11906\,
            in3 => \N__29984\,
            lcout => \tok.n898\,
            ltout => \tok.n898_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11897\,
            in3 => \N__22135\,
            lcout => \tok.uart.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5546_4_lut_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__15953\,
            in1 => \N__19895\,
            in2 => \N__12134\,
            in3 => \N__13013\,
            lcout => OPEN,
            ltout => \tok.ram.n5608_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6_4_lut_adj_23_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__15861\,
            in1 => \N__12132\,
            in2 => \N__12137\,
            in3 => \N__29985\,
            lcout => \tok.n3_adj_683\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_45_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__12133\,
            in1 => \N__18313\,
            in2 => \N__27106\,
            in3 => \N__20238\,
            lcout => OPEN,
            ltout => \tok.n83_adj_678_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5458_2_lut_3_lut_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19038\,
            in2 => \N__12104\,
            in3 => \N__29986\,
            lcout => OPEN,
            ltout => \tok.n5483_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i18_4_lut_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__12101\,
            in1 => \N__19240\,
            in2 => \N__12095\,
            in3 => \N__20239\,
            lcout => OPEN,
            ltout => \tok.n5_adj_684_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_49_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__13014\,
            in1 => \N__16293\,
            in2 => \N__12092\,
            in3 => \N__16369\,
            lcout => n92_adj_868,
            ltout => \n92_adj_868_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_83_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16171\,
            in2 => \N__12089\,
            in3 => \N__13041\,
            lcout => \tok.tc_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i5_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16172\,
            in1 => \_gnd_net_\,
            in2 => \N__13048\,
            in3 => \N__12071\,
            lcout => tc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28497\,
            ce => 'H',
            sr => \N__28212\
        );

    \tok.i1546_3_lut_4_lut_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__23793\,
            in1 => \N__16242\,
            in2 => \N__22541\,
            in3 => \N__15619\,
            lcout => \tok.table_wr_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2569_2_lut_3_lut_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__15625\,
            in1 => \_gnd_net_\,
            in2 => \N__24782\,
            in3 => \N__22502\,
            lcout => \tok.table_wr_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2570_2_lut_3_lut_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__22501\,
            in1 => \N__28867\,
            in2 => \_gnd_net_\,
            in3 => \N__15626\,
            lcout => \tok.table_wr_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1584_3_lut_4_lut_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__15620\,
            in1 => \N__22492\,
            in2 => \N__25375\,
            in3 => \N__14967\,
            lcout => \tok.table_wr_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1622_3_lut_4_lut_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__23932\,
            in1 => \N__12650\,
            in2 => \N__22540\,
            in3 => \N__15621\,
            lcout => \tok.table_wr_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1660_3_lut_4_lut_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__15622\,
            in1 => \N__22496\,
            in2 => \N__24028\,
            in3 => \N__12710\,
            lcout => \tok.table_wr_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1812_3_lut_4_lut_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__27213\,
            in1 => \N__13018\,
            in2 => \N__22542\,
            in3 => \N__15624\,
            lcout => \tok.table_wr_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1736_3_lut_4_lut_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__15623\,
            in1 => \N__22497\,
            in2 => \N__23553\,
            in3 => \N__12948\,
            lcout => \tok.table_wr_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2445_2_lut_3_lut_4_lut_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__22504\,
            in1 => \N__24351\,
            in2 => \N__15672\,
            in3 => \N__12923\,
            lcout => \tok.table_wr_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2446_2_lut_3_lut_4_lut_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__12925\,
            in1 => \N__15663\,
            in2 => \N__24488\,
            in3 => \N__22507\,
            lcout => \tok.table_wr_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2453_2_lut_3_lut_4_lut_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__22505\,
            in1 => \N__25060\,
            in2 => \N__15673\,
            in3 => \N__12924\,
            lcout => \tok.table_wr_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2462_2_lut_3_lut_4_lut_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__12926\,
            in1 => \N__15667\,
            in2 => \N__27464\,
            in3 => \N__22508\,
            lcout => \tok.table_wr_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2469_2_lut_3_lut_4_lut_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__22506\,
            in1 => \N__27538\,
            in2 => \N__15674\,
            in3 => \N__12928\,
            lcout => \tok.table_wr_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2470_2_lut_3_lut_4_lut_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__12927\,
            in1 => \N__15671\,
            in2 => \N__28073\,
            in3 => \N__22509\,
            lcout => \tok.table_wr_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1698_3_lut_4_lut_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__22503\,
            in1 => \N__22853\,
            in2 => \N__12756\,
            in3 => \N__15594\,
            lcout => \tok.table_wr_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_121_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18262\,
            in1 => \N__20231\,
            in2 => \_gnd_net_\,
            in3 => \N__29947\,
            lcout => \tok.n8_adj_790\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_219_i11_2_lut_4_lut_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__20166\,
            in1 => \N__17974\,
            in2 => \N__18315\,
            in3 => \N__29911\,
            lcout => \tok.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_118_i10_2_lut_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__29913\,
            in1 => \_gnd_net_\,
            in2 => \N__18023\,
            in3 => \_gnd_net_\,
            lcout => \tok.n10_adj_803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_2_lut_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__20162\,
            in1 => \_gnd_net_\,
            in2 => \N__18314\,
            in3 => \_gnd_net_\,
            lcout => \tok.n5318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_4_lut_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111101"
        )
    port map (
            in0 => \N__29914\,
            in1 => \N__18258\,
            in2 => \N__18024\,
            in3 => \N__20167\,
            lcout => \tok.n5293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_135_i11_2_lut_4_lut_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__20164\,
            in1 => \N__17975\,
            in2 => \N__18316\,
            in3 => \N__29912\,
            lcout => \tok.n11_adj_694\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_128_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111110111"
        )
    port map (
            in0 => \N__29910\,
            in1 => \N__18250\,
            in2 => \N__18022\,
            in3 => \N__20165\,
            lcout => \tok.n10_adj_796\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_233_i11_2_lut_4_lut_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__20168\,
            in1 => \N__17982\,
            in2 => \N__18317\,
            in3 => \N__29915\,
            lcout => \tok.n11_adj_681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_116_i9_2_lut_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18251\,
            in2 => \_gnd_net_\,
            in3 => \N__20163\,
            lcout => \tok.n9_adj_802\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_213_i11_2_lut_4_lut_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__20122\,
            in1 => \N__17934\,
            in2 => \N__18280\,
            in3 => \N__29853\,
            lcout => \tok.n11_adj_788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_111_i11_2_lut_4_lut_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29850\,
            in1 => \N__18194\,
            in2 => \N__17997\,
            in3 => \N__20120\,
            lcout => \tok.n11_adj_680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_122_i11_2_lut_4_lut_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__20121\,
            in1 => \N__17933\,
            in2 => \N__18279\,
            in3 => \N__29852\,
            lcout => \tok.n11_adj_706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_237_i11_2_lut_4_lut_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20119\,
            in1 => \N__17926\,
            in2 => \N__29927\,
            in3 => \N__18193\,
            lcout => \tok.n11_adj_793\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_214_i14_2_lut_3_lut_4_lut_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__18761\,
            in1 => \N__22063\,
            in2 => \N__18962\,
            in3 => \N__19153\,
            lcout => \tok.n14_adj_644\,
            ltout => \tok.n14_adj_644_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_154_i16_2_lut_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12269\,
            in3 => \N__13129\,
            lcout => \tok.n399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_4_lut_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100100110000"
        )
    port map (
            in0 => \N__18192\,
            in1 => \N__20118\,
            in2 => \N__17996\,
            in3 => \N__29851\,
            lcout => \tok.n8_adj_805\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_4_lut_adj_142_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__29854\,
            in1 => \N__18201\,
            in2 => \N__17998\,
            in3 => \N__20123\,
            lcout => \tok.n26_adj_750\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5256_4_lut_4_lut_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111000111"
        )
    port map (
            in0 => \N__17962\,
            in1 => \N__20124\,
            in2 => \N__18281\,
            in3 => \N__29855\,
            lcout => \tok.n5429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_67_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18908\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18213\,
            lcout => \tok.n4_adj_712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19154\,
            in1 => \N__18765\,
            in2 => \_gnd_net_\,
            in3 => \N__18909\,
            lcout => \tok.n7_adj_785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_adj_153_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000001"
        )
    port map (
            in0 => \N__29858\,
            in1 => \N__18208\,
            in2 => \N__20194\,
            in3 => \N__17965\,
            lcout => \tok.n4848\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i12_1_lut_2_lut_4_lut_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17966\,
            in1 => \N__20132\,
            in2 => \N__18283\,
            in3 => \N__29860\,
            lcout => \tok.n20_adj_663\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i20_1_lut_2_lut_4_lut_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__29859\,
            in1 => \N__18209\,
            in2 => \N__20195\,
            in3 => \N__17967\,
            lcout => \tok.n8_adj_792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5220_2_lut_4_lut_4_lut_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101111111111"
        )
    port map (
            in0 => \N__17963\,
            in1 => \N__20125\,
            in2 => \N__18282\,
            in3 => \N__29856\,
            lcout => \tok.n5391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2547_2_lut_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17964\,
            lcout => \tok.n2607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i113_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__26502\,
            in1 => \N__12298\,
            in2 => \N__26056\,
            in3 => \N__12314\,
            lcout => tail_113,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i112_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__14431\,
            in1 => \N__26012\,
            in2 => \N__14459\,
            in3 => \N__26501\,
            lcout => tail_112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_151_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__16940\,
            in1 => \N__29607\,
            in2 => \N__16859\,
            in3 => \N__14735\,
            lcout => \tok.n27_adj_825\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_154_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__14657\,
            in1 => \N__16941\,
            in2 => \N__27353\,
            in3 => \N__16853\,
            lcout => OPEN,
            ltout => \tok.n27_adj_828_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i5_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__16700\,
            in1 => \N__14697\,
            in2 => \N__12287\,
            in3 => \N__16734\,
            lcout => \tok.idx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28481\,
            ce => 'H',
            sr => \N__28234\
        );

    \tok.i50_4_lut_adj_157_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__16942\,
            in1 => \N__16854\,
            in2 => \N__21894\,
            in3 => \N__14582\,
            lcout => OPEN,
            ltout => \tok.n27_adj_831_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i6_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__16701\,
            in1 => \N__14622\,
            in2 => \N__12284\,
            in3 => \N__16735\,
            lcout => \tok.idx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28481\,
            ce => 'H',
            sr => \N__28234\
        );

    \tok.i50_4_lut_adj_160_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__16943\,
            in1 => \N__16855\,
            in2 => \N__22321\,
            in3 => \N__14513\,
            lcout => OPEN,
            ltout => \tok.n27_adj_833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i7_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__16702\,
            in1 => \N__14545\,
            in2 => \N__12281\,
            in3 => \N__16736\,
            lcout => \tok.idx_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28481\,
            ce => 'H',
            sr => \N__28234\
        );

    \tok.idx_i4_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__16733\,
            in1 => \N__16699\,
            in2 => \N__14778\,
            in3 => \N__12479\,
            lcout => \tok.idx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28481\,
            ce => 'H',
            sr => \N__28234\
        );

    \tok.i1_2_lut_3_lut_4_lut_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16923\,
            in1 => \N__12446\,
            in2 => \N__12421\,
            in3 => \N__22140\,
            lcout => \tok.n17_adj_777\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_136_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000100"
        )
    port map (
            in0 => \N__18351\,
            in1 => \N__18052\,
            in2 => \N__12380\,
            in3 => \N__20297\,
            lcout => OPEN,
            ltout => \tok.n5285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_137_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17416\,
            in1 => \N__12388\,
            in2 => \N__12473\,
            in3 => \N__30025\,
            lcout => \tok.n1_adj_715\,
            ltout => \tok.n1_adj_715_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2571_2_lut_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__12378\,
            in1 => \_gnd_net_\,
            in2 => \N__12470\,
            in3 => \_gnd_net_\,
            lcout => \tok.n190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_108_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__20298\,
            in1 => \N__18352\,
            in2 => \N__17420\,
            in3 => \N__18059\,
            lcout => OPEN,
            ltout => \tok.n10_adj_763_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_4_lut_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12389\,
            in1 => \N__12452\,
            in2 => \N__12425\,
            in3 => \N__12415\,
            lcout => \tok.n238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5175_2_lut_3_lut_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__16922\,
            in1 => \N__22139\,
            in2 => \_gnd_net_\,
            in3 => \N__19246\,
            lcout => \tok.n5340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_162_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__12377\,
            in1 => \N__12357\,
            in2 => \N__16499\,
            in3 => \N__16432\,
            lcout => \tok.n4_adj_813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_54_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__20278\,
            in1 => \N__12503\,
            in2 => \N__12494\,
            in3 => \N__19256\,
            lcout => OPEN,
            ltout => \tok.n13_adj_691_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_55_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__16353\,
            in1 => \N__16294\,
            in2 => \N__12530\,
            in3 => \N__15313\,
            lcout => n10_adj_871,
            ltout => \n10_adj_871_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_82_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16134\,
            in2 => \N__12527\,
            in3 => \N__14105\,
            lcout => \tok.tc_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5541_4_lut_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__15964\,
            in1 => \N__19897\,
            in2 => \N__14084\,
            in3 => \N__15312\,
            lcout => OPEN,
            ltout => \tok.ram.n5605_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6_4_lut_adj_24_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__14083\,
            in1 => \N__15874\,
            in2 => \N__12506\,
            in3 => \N__30031\,
            lcout => \tok.n3_adj_690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_51_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__14079\,
            in1 => \N__18350\,
            in2 => \N__17279\,
            in3 => \N__20277\,
            lcout => OPEN,
            ltout => \tok.n83_adj_687_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5480_2_lut_3_lut_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19070\,
            in2 => \N__12497\,
            in3 => \N__30030\,
            lcout => \tok.n5505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i6_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16135\,
            in1 => \_gnd_net_\,
            in2 => \N__14113\,
            in3 => \N__12485\,
            lcout => tc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28492\,
            ce => 'H',
            sr => \N__28213\
        );

    \tok.i125_4_lut_adj_198_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__18361\,
            in1 => \N__12612\,
            in2 => \N__17459\,
            in3 => \N__20311\,
            lcout => OPEN,
            ltout => \tok.n83_adj_848_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5545_2_lut_3_lut_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19058\,
            in2 => \N__12620\,
            in3 => \N__30026\,
            lcout => \tok.n5610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5527_4_lut_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__15960\,
            in1 => \N__12711\,
            in2 => \N__12617\,
            in3 => \N__19901\,
            lcout => OPEN,
            ltout => \tok.ram.n5594_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6_4_lut_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__15860\,
            in1 => \N__12616\,
            in2 => \N__12590\,
            in3 => \N__30027\,
            lcout => OPEN,
            ltout => \tok.n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__12587\,
            in1 => \N__19245\,
            in2 => \N__12581\,
            in3 => \N__20312\,
            lcout => OPEN,
            ltout => \tok.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__12712\,
            in1 => \N__16281\,
            in2 => \N__12578\,
            in3 => \N__16357\,
            lcout => n10_adj_866,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i1_4_lut_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__15995\,
            in1 => \N__17048\,
            in2 => \N__17330\,
            in3 => \N__12575\,
            lcout => \rx_data_7__N_511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_65_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19057\,
            in2 => \_gnd_net_\,
            in3 => \N__18360\,
            lcout => \tok.n101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i11_4_lut_adj_103_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12872\,
            in1 => \N__12560\,
            in2 => \N__12548\,
            in3 => \N__12887\,
            lcout => \tok.n27_adj_757\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_adj_81_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__12559\,
            in1 => \N__12544\,
            in2 => \N__21631\,
            in3 => \N__29266\,
            lcout => OPEN,
            ltout => \tok.n21_adj_733_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i14_4_lut_adj_107_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12845\,
            in1 => \N__12857\,
            in2 => \N__12533\,
            in3 => \N__12851\,
            lcout => \tok.n30_adj_761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_71_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__12886\,
            in1 => \N__12871\,
            in2 => \N__22320\,
            in3 => \N__22757\,
            lcout => \tok.n22_adj_721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_79_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__12838\,
            in1 => \N__12796\,
            in2 => \N__25765\,
            in3 => \N__25158\,
            lcout => \tok.n23_adj_731\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_4_lut_adj_33_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__12826\,
            in1 => \N__12808\,
            in2 => \N__24862\,
            in3 => \N__29070\,
            lcout => \tok.n24_adj_651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i12_4_lut_adj_101_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12839\,
            in1 => \N__12827\,
            in2 => \N__12812\,
            in3 => \N__12797\,
            lcout => \tok.n28_adj_755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__21619\,
            in1 => \N__24481\,
            in2 => \N__27460\,
            in3 => \N__29267\,
            lcout => \tok.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_2_lut_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12784\,
            in2 => \_gnd_net_\,
            in3 => \N__12719\,
            lcout => \tok.tc_plus_1_0\,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \tok.n4754\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_3_lut_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15726\,
            in2 => \_gnd_net_\,
            in3 => \N__12686\,
            lcout => \tok.tc_plus_1_1\,
            ltout => OPEN,
            carryin => \tok.n4754\,
            carryout => \tok.n4755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_4_lut_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12683\,
            in2 => \_gnd_net_\,
            in3 => \N__12623\,
            lcout => \tok.tc_plus_1_2\,
            ltout => OPEN,
            carryin => \tok.n4755\,
            carryout => \tok.n4756\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_5_lut_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13090\,
            in3 => \N__13055\,
            lcout => \tok.tc_plus_1_3\,
            ltout => OPEN,
            carryin => \tok.n4756\,
            carryout => \tok.n4757\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_6_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16106\,
            in2 => \_gnd_net_\,
            in3 => \N__13052\,
            lcout => \tok.tc_plus_1_4\,
            ltout => OPEN,
            carryin => \tok.n4757\,
            carryout => \tok.n4758\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_7_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13040\,
            in2 => \_gnd_net_\,
            in3 => \N__12995\,
            lcout => \tok.tc_plus_1_5\,
            ltout => OPEN,
            carryin => \tok.n4758\,
            carryout => \tok.n4759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_8_lut_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14112\,
            in2 => \_gnd_net_\,
            in3 => \N__12992\,
            lcout => \tok.tc_plus_1_6\,
            ltout => OPEN,
            carryin => \tok.n4759\,
            carryout => \tok.n4760\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_7__I_0_9_lut_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12989\,
            in2 => \_gnd_net_\,
            in3 => \N__12962\,
            lcout => \tok.tc_plus_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5608_2_lut_3_lut_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000100"
        )
    port map (
            in0 => \N__17611\,
            in1 => \N__18386\,
            in2 => \N__22510\,
            in3 => \_gnd_net_\,
            lcout => \tok.write_flag\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5234_4_lut_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__18385\,
            in1 => \N__17610\,
            in2 => \N__12932\,
            in3 => \N__15589\,
            lcout => \tok.n5406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_157_i15_2_lut_3_lut_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__17528\,
            in1 => \N__15815\,
            in2 => \_gnd_net_\,
            in3 => \N__15423\,
            lcout => \tok.n15_adj_671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__12893\,
            in1 => \_gnd_net_\,
            in2 => \N__23278\,
            in3 => \N__15590\,
            lcout => OPEN,
            ltout => \tok.n14_adj_688_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2652_4_lut_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__13178\,
            in1 => \N__15814\,
            in2 => \N__13166\,
            in3 => \N__13097\,
            lcout => \tok.n2735\,
            ltout => \tok.n2735_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_4_i1_3_lut_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27756\,
            in2 => \N__13163\,
            in3 => \N__19042\,
            lcout => OPEN,
            ltout => \tok.n1_adj_850_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_186_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__23212\,
            in1 => \N__13253\,
            in2 => \N__13160\,
            in3 => \N__21632\,
            lcout => \tok.n17_adj_853\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_155_i16_2_lut_3_lut_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__15424\,
            in1 => \N__22450\,
            in2 => \_gnd_net_\,
            in3 => \N__17529\,
            lcout => \tok.n400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_98_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__13157\,
            in1 => \N__13151\,
            in2 => \N__16004\,
            in3 => \N__19681\,
            lcout => \tok.n5254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5210_4_lut_4_lut_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__15419\,
            in1 => \N__23258\,
            in2 => \N__17531\,
            in3 => \N__15451\,
            lcout => \tok.n5380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_129_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111111"
        )
    port map (
            in0 => \N__17598\,
            in1 => \N__15417\,
            in2 => \N__13145\,
            in3 => \N__13128\,
            lcout => OPEN,
            ltout => \tok.n5271_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_130_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111111"
        )
    port map (
            in0 => \N__15418\,
            in1 => \N__15450\,
            in2 => \N__13112\,
            in3 => \N__23377\,
            lcout => \tok.n5272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_56_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__13109\,
            in1 => \N__13103\,
            in2 => \N__17612\,
            in3 => \N__19680\,
            lcout => \tok.n15_adj_695\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i4_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13262\,
            in1 => \N__23039\,
            in2 => \_gnd_net_\,
            in3 => \N__25679\,
            lcout => uart_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_4_i12_2_lut_3_lut_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__23259\,
            in1 => \N__13261\,
            in2 => \_gnd_net_\,
            in3 => \N__22411\,
            lcout => \tok.n12_adj_826\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_213_i15_2_lut_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__13237\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17487\,
            lcout => \tok.n15_adj_789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i3_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13208\,
            in1 => \N__14366\,
            in2 => \_gnd_net_\,
            in3 => \N__27755\,
            lcout => sender_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28527\,
            ce => \N__14300\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i4_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14367\,
            in1 => \N__13202\,
            in2 => \_gnd_net_\,
            in3 => \N__21131\,
            lcout => \tok.uart.sender_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28527\,
            ce => \N__14300\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i5_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13196\,
            in1 => \N__14368\,
            in2 => \_gnd_net_\,
            in3 => \N__22758\,
            lcout => \tok.uart.sender_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28527\,
            ce => \N__14300\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i6_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14369\,
            in1 => \N__13190\,
            in2 => \_gnd_net_\,
            in3 => \N__29731\,
            lcout => \tok.uart.sender_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28527\,
            ce => \N__14300\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i7_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13184\,
            in1 => \N__14370\,
            in2 => \_gnd_net_\,
            in3 => \N__29596\,
            lcout => \tok.uart.sender_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28527\,
            ce => \N__14300\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i8_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14371\,
            in1 => \N__14306\,
            in2 => \_gnd_net_\,
            in3 => \N__27347\,
            lcout => \tok.uart.sender_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28527\,
            ce => \N__14300\,
            sr => \_gnd_net_\
        );

    \tok.uart.sender_i9_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14408\,
            in1 => \N__14372\,
            in2 => \_gnd_net_\,
            in3 => \N__21893\,
            lcout => \tok.uart.sender_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28527\,
            ce => \N__14300\,
            sr => \_gnd_net_\
        );

    \tok.equal_114_i10_2_lut_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18002\,
            in2 => \_gnd_net_\,
            in3 => \N__29958\,
            lcout => \tok.n10_adj_643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i6_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14024\,
            in1 => \N__14070\,
            in2 => \N__13721\,
            in3 => \N__13748\,
            lcout => \tok.C_stk.tail_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28530\,
            ce => \N__13362\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.i5265_3_lut_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14053\,
            in1 => \N__14270\,
            in2 => \_gnd_net_\,
            in3 => \N__15314\,
            lcout => OPEN,
            ltout => \tok.C_stk.n5438_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.C_stk.head_i0_i6_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__14185\,
            in1 => \N__15517\,
            in2 => \N__14117\,
            in3 => \N__14114\,
            lcout => \tok.c_stk_r_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28530\,
            ce => \N__13362\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i14_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__14054\,
            in1 => \N__13716\,
            in2 => \N__13396\,
            in3 => \N__14025\,
            lcout => \tok.tail_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28530\,
            ce => \N__13362\,
            sr => \_gnd_net_\
        );

    \tok.C_stk.tail_i0_i22_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14023\,
            in1 => \N__13747\,
            in2 => \N__13739\,
            in3 => \N__13720\,
            lcout => \tok.C_stk.tail_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28530\,
            ce => \N__13362\,
            sr => \_gnd_net_\
        );

    \tok.tc_i1_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15752\,
            in1 => \N__16204\,
            in2 => \_gnd_net_\,
            in3 => \N__15722\,
            lcout => tc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28535\,
            ce => 'H',
            sr => \N__28128\
        );

    \tok.inv_106_i14_1_lut_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23154\,
            lcout => \tok.n289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.reset_I_0_1_lut_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14507\,
            lcout => \tok.reset_N_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i16_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14486\,
            in1 => \N__14417\,
            in2 => \_gnd_net_\,
            in3 => \N__26402\,
            lcout => \tok.A_stk.tail_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28482\,
            ce => \N__26019\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i0_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26401\,
            in1 => \_gnd_net_\,
            in2 => \N__14498\,
            in3 => \N__22840\,
            lcout => \tok.A_stk.tail_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28482\,
            ce => \N__26019\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i32_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14477\,
            in1 => \N__14494\,
            in2 => \_gnd_net_\,
            in3 => \N__26403\,
            lcout => \tok.A_stk.tail_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28482\,
            ce => \N__26019\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i48_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26404\,
            in1 => \N__14485\,
            in2 => \_gnd_net_\,
            in3 => \N__14468\,
            lcout => \tok.A_stk.tail_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28482\,
            ce => \N__26019\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i64_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14476\,
            in1 => \N__14441\,
            in2 => \_gnd_net_\,
            in3 => \N__26405\,
            lcout => \tok.A_stk.tail_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28482\,
            ce => \N__26019\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i80_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26406\,
            in1 => \_gnd_net_\,
            in2 => \N__14432\,
            in3 => \N__14467\,
            lcout => \tok.A_stk.tail_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28482\,
            ce => \N__26019\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i96_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14458\,
            in1 => \N__14440\,
            in2 => \_gnd_net_\,
            in3 => \N__26407\,
            lcout => tail_96,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28482\,
            ce => \N__26019\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i0_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14416\,
            in1 => \N__25466\,
            in2 => \_gnd_net_\,
            in3 => \N__27783\,
            lcout => \tok.S_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28482\,
            ce => \N__26019\,
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_2_lut_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__14849\,
            in1 => \N__14848\,
            in2 => \N__15229\,
            in3 => \N__14813\,
            lcout => \tok.n33\,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \tok.n4747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_3_lut_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__16631\,
            in1 => \N__16630\,
            in2 => \N__15233\,
            in3 => \N__14810\,
            lcout => \tok.n33_adj_814\,
            ltout => OPEN,
            carryin => \tok.n4747\,
            carryout => \tok.n4748\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_4_lut_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__16974\,
            in1 => \N__16973\,
            in2 => \N__15230\,
            in3 => \N__14807\,
            lcout => \tok.n33_adj_816\,
            ltout => OPEN,
            carryin => \tok.n4748\,
            carryout => \tok.n4749\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_5_lut_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__16769\,
            in1 => \N__16768\,
            in2 => \N__15234\,
            in3 => \N__14804\,
            lcout => \tok.n33_adj_821\,
            ltout => OPEN,
            carryin => \tok.n4749\,
            carryout => \tok.n4750\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_6_lut_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__14768\,
            in1 => \N__14767\,
            in2 => \N__15231\,
            in3 => \N__14729\,
            lcout => \tok.n33_adj_819\,
            ltout => OPEN,
            carryin => \tok.n4750\,
            carryout => \tok.n4751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_7_lut_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__14696\,
            in1 => \N__14695\,
            in2 => \N__15235\,
            in3 => \N__14651\,
            lcout => \tok.n33_adj_811\,
            ltout => OPEN,
            carryin => \tok.n4751\,
            carryout => \tok.n4752\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_8_lut_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__14615\,
            in1 => \N__14614\,
            in2 => \N__15232\,
            in3 => \N__14576\,
            lcout => \tok.n33_adj_804\,
            ltout => OPEN,
            carryin => \tok.n4752\,
            carryout => \tok.n4753\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_7__I_0_9_lut_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__14552\,
            in1 => \N__14553\,
            in2 => \N__15236\,
            in3 => \N__14516\,
            lcout => \tok.n33_adj_801\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16837\,
            in2 => \_gnd_net_\,
            in3 => \N__15186\,
            lcout => \tok.n5\,
            ltout => \tok.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_72_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010111011"
        )
    port map (
            in0 => \N__17768\,
            in1 => \N__15560\,
            in2 => \N__14897\,
            in3 => \N__16930\,
            lcout => \stall_\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.stall_200_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111111001101"
        )
    port map (
            in0 => \N__16933\,
            in1 => \N__17771\,
            in2 => \N__15566\,
            in3 => \N__14894\,
            lcout => \tok.stall\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28493\,
            ce => 'H',
            sr => \N__28237\
        );

    \tok.i1_4_lut_adj_132_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__17770\,
            in1 => \N__15562\,
            in2 => \N__16857\,
            in3 => \N__16931\,
            lcout => \tok.n5282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.search_clk_198_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16844\,
            lcout => \tok.search_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28493\,
            ce => 'H',
            sr => \N__28237\
        );

    \tok.i50_4_lut_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__27770\,
            in1 => \N__14888\,
            in2 => \N__16856\,
            in3 => \N__16932\,
            lcout => OPEN,
            ltout => \tok.n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i0_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__14850\,
            in1 => \N__16693\,
            in2 => \N__14882\,
            in3 => \N__16729\,
            lcout => \tok.idx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28493\,
            ce => 'H',
            sr => \N__28237\
        );

    \tok.i2622_2_lut_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__17769\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15561\,
            lcout => \tok.n2699\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_34_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__18367\,
            in1 => \N__15018\,
            in2 => \N__15395\,
            in3 => \N__20313\,
            lcout => OPEN,
            ltout => \tok.n83_adj_652_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5442_2_lut_3_lut_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19071\,
            in2 => \N__14816\,
            in3 => \N__30028\,
            lcout => \tok.n5460\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5518_4_lut_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__15965\,
            in1 => \N__14976\,
            in2 => \N__19904\,
            in3 => \N__15019\,
            lcout => OPEN,
            ltout => \tok.ram.n5580_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6_4_lut_adj_21_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__15020\,
            in1 => \N__15873\,
            in2 => \N__14993\,
            in3 => \N__30029\,
            lcout => OPEN,
            ltout => \tok.n3_adj_659_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_37_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__14990\,
            in1 => \N__19258\,
            in2 => \N__14984\,
            in3 => \N__20315\,
            lcout => OPEN,
            ltout => \tok.n13_adj_660_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_39_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__14977\,
            in1 => \N__16370\,
            in2 => \N__14948\,
            in3 => \N__16309\,
            lcout => n92_adj_867,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_4_lut_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__18368\,
            in1 => \N__19257\,
            in2 => \N__18836\,
            in3 => \N__20314\,
            lcout => OPEN,
            ltout => \tok.n4_adj_778_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_115_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18046\,
            in1 => \N__14923\,
            in2 => \N__14912\,
            in3 => \N__19072\,
            lcout => \tok.n797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_106_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111110"
        )
    port map (
            in0 => \N__29468\,
            in1 => \N__17018\,
            in2 => \N__15113\,
            in3 => \N__15274\,
            lcout => OPEN,
            ltout => \tok.n26_adj_760_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5526_4_lut_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15026\,
            in1 => \N__15104\,
            in2 => \N__14909\,
            in3 => \N__14906\,
            lcout => OPEN,
            ltout => \tok.n5587_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_138_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001000100"
        )
    port map (
            in0 => \N__15640\,
            in1 => \N__16949\,
            in2 => \N__14900\,
            in3 => \N__15242\,
            lcout => \tok.found_slot\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_102_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15128\,
            in1 => \N__17036\,
            in2 => \N__15275\,
            in3 => \N__15143\,
            lcout => OPEN,
            ltout => \tok.n26_adj_756_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i15_4_lut_adj_126_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15257\,
            in1 => \N__15062\,
            in2 => \N__15251\,
            in3 => \N__15248\,
            lcout => \tok.found_slot_N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_adj_145_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15641\,
            in2 => \_gnd_net_\,
            in3 => \N__15185\,
            lcout => \tok.write_slot\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__15142\,
            in1 => \N__15127\,
            in2 => \N__27351\,
            in3 => \N__29724\,
            lcout => \tok.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_105_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__21109\,
            in1 => \N__15076\,
            in2 => \N__15098\,
            in3 => \N__29597\,
            lcout => \tok.n18_adj_759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_104_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15040\,
            in1 => \N__15094\,
            in2 => \N__15080\,
            in3 => \N__15055\,
            lcout => \tok.n25_adj_758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5505_4_lut_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__15056\,
            in1 => \N__21886\,
            in2 => \N__27782\,
            in3 => \N__15041\,
            lcout => \tok.n5590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_175_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__25159\,
            in1 => \N__20657\,
            in2 => \_gnd_net_\,
            in3 => \N__23402\,
            lcout => \tok.n6_adj_843\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i6_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22916\,
            in1 => \N__25660\,
            in2 => \_gnd_net_\,
            in3 => \N__15356\,
            lcout => uart_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_6_i12_2_lut_3_lut_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__15355\,
            in1 => \N__22511\,
            in2 => \_gnd_net_\,
            in3 => \N__23314\,
            lcout => \tok.n12_adj_824\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_176_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101110"
        )
    port map (
            in0 => \N__15347\,
            in1 => \N__23813\,
            in2 => \N__23335\,
            in3 => \N__15337\,
            lcout => OPEN,
            ltout => \tok.n31_adj_844_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_177_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__22539\,
            in1 => \N__18047\,
            in2 => \N__15341\,
            in3 => \N__19511\,
            lcout => \tok.n10_adj_845\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i3_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__15338\,
            in1 => \_gnd_net_\,
            in2 => \N__15329\,
            in3 => \N__25680\,
            lcout => uart_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_4_lut_adj_188_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__28730\,
            in1 => \N__23665\,
            in2 => \N__18509\,
            in3 => \N__29167\,
            lcout => \tok.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i2_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21183\,
            in1 => \N__17344\,
            in2 => \_gnd_net_\,
            in3 => \N__22975\,
            lcout => capture_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i4_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22977\,
            in1 => \N__23035\,
            in2 => \_gnd_net_\,
            in3 => \N__15324\,
            lcout => capture_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i3_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15325\,
            in1 => \N__17343\,
            in2 => \_gnd_net_\,
            in3 => \N__22976\,
            lcout => capture_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1774_3_lut_4_lut_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__23667\,
            in1 => \N__15311\,
            in2 => \N__22547\,
            in3 => \N__15629\,
            lcout => \tok.table_wr_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_219_i10_2_lut_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18034\,
            in2 => \_gnd_net_\,
            in3 => \N__30013\,
            lcout => \tok.n10_adj_747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2573_3_lut_4_lut_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__15432\,
            in1 => \N__15627\,
            in2 => \N__22545\,
            in3 => \N__17613\,
            lcout => \tok.n2635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2620_3_lut_4_lut_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__15628\,
            in1 => \N__15464\,
            in2 => \N__26979\,
            in3 => \N__22523\,
            lcout => \tok.n2697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2460_3_lut_4_lut_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__15433\,
            in1 => \N__15508\,
            in2 => \N__22546\,
            in3 => \N__17614\,
            lcout => \tok.n2520\,
            ltout => \tok.n2520_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2587_4_lut_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__22527\,
            in1 => \N__15458\,
            in2 => \N__15437\,
            in3 => \N__15434\,
            lcout => \tok.n2661\,
            ltout => \tok.n2661_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_179_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__15391\,
            in1 => \N__25369\,
            in2 => \N__15368\,
            in3 => \N__26958\,
            lcout => OPEN,
            ltout => \tok.n9_adj_847_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5562_4_lut_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__15365\,
            in1 => \N__18398\,
            in2 => \N__15359\,
            in3 => \N__19754\,
            lcout => \tok.n5566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__15971\,
            in1 => \N__18420\,
            in2 => \_gnd_net_\,
            in3 => \N__18983\,
            lcout => \tok.n880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_116_i14_2_lut_3_lut_4_lut_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__22109\,
            in1 => \N__18791\,
            in2 => \N__19043\,
            in3 => \N__19217\,
            lcout => \tok.n14_adj_701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__19216\,
            in1 => \N__18979\,
            in2 => \N__18815\,
            in3 => \N__22108\,
            lcout => \tok.n14_adj_807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5260_4_lut_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__15806\,
            in1 => \N__17483\,
            in2 => \N__16013\,
            in3 => \N__15794\,
            lcout => OPEN,
            ltout => \tok.n5433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_133_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__15767\,
            in1 => \N__15758\,
            in2 => \N__15788\,
            in3 => \N__15785\,
            lcout => \tok.n2743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_131_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100000"
        )
    port map (
            in0 => \N__15680\,
            in1 => \N__17482\,
            in2 => \N__15779\,
            in3 => \N__15766\,
            lcout => \tok.n5175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_88_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15748\,
            in1 => \N__16162\,
            in2 => \_gnd_net_\,
            in3 => \N__15727\,
            lcout => \tok.tc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i8_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22993\,
            in1 => \N__15991\,
            in2 => \_gnd_net_\,
            in3 => \N__22978\,
            lcout => capture_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28528\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_213_i14_2_lut_3_lut_4_lut_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__18777\,
            in1 => \N__19167\,
            in2 => \N__22107\,
            in3 => \N__19044\,
            lcout => \tok.n14_adj_765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_174_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101011"
        )
    port map (
            in0 => \N__18016\,
            in1 => \N__20240\,
            in2 => \N__30014\,
            in3 => \N__18354\,
            lcout => \tok.n2_adj_808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5250_3_lut_4_lut_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29962\,
            in2 => \N__20279\,
            in3 => \N__18017\,
            lcout => \tok.n5423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_4_lut_adj_143_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__18019\,
            in1 => \N__20245\,
            in2 => \N__30016\,
            in3 => \N__18356\,
            lcout => \tok.n42_adj_751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i9_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17151\,
            in1 => \N__15990\,
            in2 => \_gnd_net_\,
            in3 => \N__22982\,
            lcout => capture_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_3_lut_adj_173_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__19168\,
            in1 => \N__22077\,
            in2 => \_gnd_net_\,
            in3 => \N__18778\,
            lcout => \tok.n878\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5588_4_lut_4_lut_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000101110101"
        )
    port map (
            in0 => \N__18357\,
            in1 => \N__29969\,
            in2 => \N__20280\,
            in3 => \N__18020\,
            lcout => \tok.n5470\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2549_2_lut_4_lut_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18018\,
            in1 => \N__20244\,
            in2 => \N__30015\,
            in3 => \N__18355\,
            lcout => \tok.n2609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i5514_4_lut_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__15946\,
            in1 => \N__16251\,
            in2 => \N__16072\,
            in3 => \N__19888\,
            lcout => OPEN,
            ltout => \tok.ram.n5577_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.ram.i6_4_lut_adj_22_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__30020\,
            in1 => \N__16067\,
            in2 => \N__15893\,
            in3 => \N__15882\,
            lcout => \tok.n3_adj_672\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i27_4_lut_adj_42_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__15821\,
            in1 => \N__19215\,
            in2 => \N__16034\,
            in3 => \N__20276\,
            lcout => OPEN,
            ltout => \tok.n13_adj_673_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_44_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__16394\,
            in1 => \N__16316\,
            in2 => \N__16256\,
            in3 => \N__16252\,
            lcout => n10_adj_870,
            ltout => \n10_adj_870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i26_3_lut_adj_85_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16094\,
            in2 => \N__16223\,
            in3 => \N__16163\,
            lcout => \tok.tc_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.tc_i4_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16164\,
            in1 => \_gnd_net_\,
            in2 => \N__16104\,
            in3 => \N__16112\,
            lcout => tc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28536\,
            ce => 'H',
            sr => \N__28174\
        );

    \tok.i5568_3_lut_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__28751\,
            in1 => \N__18083\,
            in2 => \_gnd_net_\,
            in3 => \N__23931\,
            lcout => \tok.n5571\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i125_4_lut_adj_40_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__16073\,
            in1 => \N__18334\,
            in2 => \N__17402\,
            in3 => \N__20230\,
            lcout => OPEN,
            ltout => \tok.n83_adj_665_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5463_2_lut_3_lut_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19053\,
            in2 => \N__16037\,
            in3 => \N__30021\,
            lcout => \tok.n5487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i110_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17201\,
            in1 => \N__16024\,
            in2 => \_gnd_net_\,
            in3 => \N__26393\,
            lcout => tail_110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28487\,
            ce => \N__26047\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i94_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26400\,
            in1 => \N__17215\,
            in2 => \_gnd_net_\,
            in3 => \N__16561\,
            lcout => \tok.A_stk.tail_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28487\,
            ce => \N__26047\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i78_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16025\,
            in1 => \N__16552\,
            in2 => \_gnd_net_\,
            in3 => \N__26399\,
            lcout => \tok.A_stk.tail_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28487\,
            ce => \N__26047\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i62_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26398\,
            in1 => \N__16543\,
            in2 => \_gnd_net_\,
            in3 => \N__16562\,
            lcout => \tok.A_stk.tail_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28487\,
            ce => \N__26047\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i46_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16534\,
            in1 => \N__16553\,
            in2 => \_gnd_net_\,
            in3 => \N__26397\,
            lcout => \tok.A_stk.tail_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28487\,
            ce => \N__26047\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i30_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26396\,
            in1 => \N__25072\,
            in2 => \_gnd_net_\,
            in3 => \N__16544\,
            lcout => \tok.A_stk.tail_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28487\,
            ce => \N__26047\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i14_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16535\,
            in1 => \N__26395\,
            in2 => \_gnd_net_\,
            in3 => \N__28868\,
            lcout => \tok.A_stk.tail_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28487\,
            ce => \N__26047\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i111_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26394\,
            in1 => \N__16526\,
            in2 => \_gnd_net_\,
            in3 => \N__24667\,
            lcout => tail_111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28487\,
            ce => \N__26047\,
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_140_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__16939\,
            in1 => \N__16505\,
            in2 => \N__16858\,
            in3 => \N__21143\,
            lcout => \tok.n27_adj_815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_69_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16498\,
            in2 => \_gnd_net_\,
            in3 => \N__16442\,
            lcout => OPEN,
            ltout => \tok.depth_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_96_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__28582\,
            in1 => \N__16934\,
            in2 => \N__16412\,
            in3 => \N__16409\,
            lcout => \tok.n995\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i50_4_lut_adj_144_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__22761\,
            in1 => \N__16848\,
            in2 => \N__16948\,
            in3 => \N__16400\,
            lcout => OPEN,
            ltout => \tok.n27_adj_818_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i2_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__16975\,
            in1 => \N__16697\,
            in2 => \N__17009\,
            in3 => \N__16731\,
            lcout => \tok.idx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28494\,
            ce => 'H',
            sr => \N__28232\
        );

    \tok.i50_4_lut_adj_148_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__16935\,
            in1 => \N__16865\,
            in2 => \N__29738\,
            in3 => \N__16849\,
            lcout => OPEN,
            ltout => \tok.n27_adj_822_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.idx_i3_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__16770\,
            in1 => \N__16698\,
            in2 => \N__16805\,
            in3 => \N__16732\,
            lcout => \tok.idx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28494\,
            ce => 'H',
            sr => \N__28232\
        );

    \tok.idx_i1_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110100001100"
        )
    port map (
            in0 => \N__16730\,
            in1 => \N__16632\,
            in2 => \N__16703\,
            in3 => \N__16667\,
            lcout => \tok.idx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28494\,
            ce => 'H',
            sr => \N__28232\
        );

    \tok.i567_2_lut_4_lut_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001111"
        )
    port map (
            in0 => \N__16586\,
            in1 => \N__17677\,
            in2 => \N__16598\,
            in3 => \N__19324\,
            lcout => \rd_15__N_301\,
            ltout => \rd_15__N_301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i120_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__26194\,
            in1 => \N__18616\,
            in2 => \N__16601\,
            in3 => \N__18596\,
            lcout => tail_120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i119_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__18653\,
            in1 => \N__25870\,
            in2 => \N__18682\,
            in3 => \N__26193\,
            lcout => tail_119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2563_2_lut_4_lut_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19323\,
            in1 => \N__16594\,
            in2 => \N__17678\,
            in3 => \N__16585\,
            lcout => \A_stk_delta_1\,
            ltout => \A_stk_delta_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i117_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__24914\,
            in1 => \N__24925\,
            in2 => \N__16565\,
            in3 => \N__25869\,
            lcout => tail_117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i121_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__26195\,
            in1 => \N__18481\,
            in2 => \N__25926\,
            in3 => \N__18470\,
            lcout => tail_121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i115_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__18536\,
            in1 => \N__25868\,
            in2 => \N__18551\,
            in3 => \N__26192\,
            lcout => tail_115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i126_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__26196\,
            in1 => \N__17219\,
            in2 => \N__25927\,
            in3 => \N__17197\,
            lcout => tail_126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i95_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17176\,
            in1 => \N__24641\,
            in2 => \_gnd_net_\,
            in3 => \N__26246\,
            lcout => \tok.A_stk.tail_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28505\,
            ce => \N__26020\,
            sr => \_gnd_net_\
        );

    \tok.or_99_i9_2_lut_3_lut_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__22170\,
            in1 => \N__29586\,
            in2 => \_gnd_net_\,
            in3 => \N__22144\,
            lcout => \tok.n181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i2_3_lut_adj_28_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__17077\,
            in1 => \_gnd_net_\,
            in2 => \N__17111\,
            in3 => \N__17158\,
            lcout => \tok.uart.n5235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.i5204_2_lut_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17107\,
            in2 => \_gnd_net_\,
            in3 => \N__17076\,
            lcout => \tok.uart.n5374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.key_rd_15__I_0_241_i14_2_lut_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17035\,
            in2 => \_gnd_net_\,
            in3 => \N__23157\,
            lcout => \tok.n14_adj_647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25661\,
            in1 => \N__17306\,
            in2 => \_gnd_net_\,
            in3 => \N__17293\,
            lcout => uart_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i0_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17305\,
            in1 => \N__17320\,
            in2 => \_gnd_net_\,
            in3 => \N__22973\,
            lcout => capture_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i1_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22974\,
            in1 => \N__17304\,
            in2 => \_gnd_net_\,
            in3 => \N__21184\,
            lcout => capture_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_125_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__23410\,
            in1 => \N__29469\,
            in2 => \N__17294\,
            in3 => \N__23334\,
            lcout => OPEN,
            ltout => \tok.n6_adj_794_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_159_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__22781\,
            in1 => \N__20477\,
            in2 => \N__17282\,
            in3 => \N__22550\,
            lcout => \tok.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_5_i3_3_lut_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28949\,
            in1 => \N__27754\,
            in2 => \_gnd_net_\,
            in3 => \N__18818\,
            lcout => \tok.n3_adj_859\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5577_4_lut_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110110"
        )
    port map (
            in0 => \N__21111\,
            in1 => \N__19259\,
            in2 => \N__19430\,
            in3 => \N__28950\,
            lcout => OPEN,
            ltout => \tok.n5553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5576_4_lut_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__17275\,
            in1 => \N__23573\,
            in2 => \N__17249\,
            in3 => \N__26973\,
            lcout => \tok.n5552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_adj_111_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__26974\,
            in1 => \N__17246\,
            in2 => \_gnd_net_\,
            in3 => \N__19613\,
            lcout => \tok.n15_adj_770\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_adj_84_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__17234\,
            in1 => \N__26972\,
            in2 => \_gnd_net_\,
            in3 => \N__19625\,
            lcout => OPEN,
            ltout => \tok.n14_adj_735_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_adj_91_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__27940\,
            in1 => \N__20798\,
            in2 => \N__17423\,
            in3 => \N__29598\,
            lcout => \tok.n18_adj_739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_99_i6_3_lut_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__19049\,
            in1 => \N__18817\,
            in2 => \_gnd_net_\,
            in3 => \N__21110\,
            lcout => \tok.n184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_100_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__18816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19048\,
            lcout => \tok.n6_adj_754\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_185_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__27850\,
            in1 => \N__20642\,
            in2 => \N__29608\,
            in3 => \N__27633\,
            lcout => \tok.n13_adj_852\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_adj_184_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__17401\,
            in1 => \N__23696\,
            in2 => \_gnd_net_\,
            in3 => \N__26954\,
            lcout => OPEN,
            ltout => \tok.n16_adj_851_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5507_4_lut_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__19037\,
            in1 => \N__19442\,
            in2 => \N__17375\,
            in3 => \N__28971\,
            lcout => OPEN,
            ltout => \tok.n5562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5569_4_lut_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17372\,
            in1 => \N__17351\,
            in2 => \N__17360\,
            in3 => \N__17357\,
            lcout => \tok.n5561\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_4_lut_adj_187_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__23776\,
            in1 => \N__17825\,
            in2 => \N__28762\,
            in3 => \N__29149\,
            lcout => \tok.n14_adj_854\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i2_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17345\,
            in1 => \N__23365\,
            in2 => \_gnd_net_\,
            in3 => \N__25681\,
            lcout => uart_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5570_4_lut_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__19349\,
            in1 => \N__26960\,
            in2 => \N__17570\,
            in3 => \N__20012\,
            lcout => OPEN,
            ltout => \tok.n5463_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5555_4_lut_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__19913\,
            in1 => \N__17543\,
            in2 => \N__17534\,
            in3 => \N__27563\,
            lcout => \tok.n5462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_109_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011101"
        )
    port map (
            in0 => \N__29148\,
            in1 => \N__17530\,
            in2 => \N__17638\,
            in3 => \N__17491\,
            lcout => \tok.n8_adj_767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_215_i15_2_lut_3_lut_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__18421\,
            in1 => \N__19693\,
            in2 => \_gnd_net_\,
            in3 => \N__19050\,
            lcout => \tok.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5170_2_lut_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26710\,
            in2 => \_gnd_net_\,
            in3 => \N__28904\,
            lcout => \tok.n5334\,
            ltout => \tok.n5334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_166_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__26959\,
            in1 => \N__17458\,
            in2 => \N__17426\,
            in3 => \N__18335\,
            lcout => \tok.n8_adj_837\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_181_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__19051\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18422\,
            lcout => \tok.n14_adj_679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i2_1_lut_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21103\,
            lcout => \tok.n301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i11_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__27452\,
            in1 => \N__26858\,
            in2 => \N__28636\,
            in3 => \N__19919\,
            lcout => \tok.A_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28532\,
            ce => \N__28285\,
            sr => \N__28192\
        );

    \tok.A_i12_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011111000100"
        )
    port map (
            in0 => \N__26859\,
            in1 => \N__28618\,
            in2 => \N__20942\,
            in3 => \N__25061\,
            lcout => \tok.A_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28532\,
            ce => \N__28285\,
            sr => \N__28192\
        );

    \tok.A_i1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__28619\,
            in1 => \N__26860\,
            in2 => \N__17663\,
            in3 => \N__22886\,
            lcout => \tok.A_low_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28532\,
            ce => \N__28285\,
            sr => \N__28192\
        );

    \tok.A_i2_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111110101010"
        )
    port map (
            in0 => \N__24031\,
            in1 => \N__19517\,
            in2 => \N__26869\,
            in3 => \N__28620\,
            lcout => \tok.A_low_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28532\,
            ce => \N__28285\,
            sr => \N__28192\
        );

    \tok.A_i3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__23924\,
            in1 => \N__26864\,
            in2 => \N__28637\,
            in3 => \N__19760\,
            lcout => \tok.A_low_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28532\,
            ce => \N__28285\,
            sr => \N__28192\
        );

    \tok.A_i4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000101110"
        )
    port map (
            in0 => \N__25374\,
            in1 => \N__28624\,
            in2 => \N__26870\,
            in3 => \N__17654\,
            lcout => \tok.A_low_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28532\,
            ce => \N__28285\,
            sr => \N__28192\
        );

    \tok.A_i5_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__28625\,
            in1 => \N__26868\,
            in2 => \N__23794\,
            in3 => \N__17648\,
            lcout => \tok.A_low_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28532\,
            ce => \N__28285\,
            sr => \N__28192\
        );

    \tok.i2_4_lut_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24030\,
            in1 => \N__29545\,
            in2 => \N__23792\,
            in3 => \N__21084\,
            lcout => \tok.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i7_1_lut_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21867\,
            lcout => \tok.n296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_110_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__21868\,
            in1 => \N__20783\,
            in2 => \_gnd_net_\,
            in3 => \N__27914\,
            lcout => \tok.n14_adj_769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_220_i15_2_lut_3_lut_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__17639\,
            in1 => \N__22480\,
            in2 => \_gnd_net_\,
            in3 => \N__17615\,
            lcout => \tok.n15_adj_655\,
            ltout => \tok.n15_adj_655_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_135_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001011101"
        )
    port map (
            in0 => \N__17745\,
            in1 => \N__17813\,
            in2 => \N__17774\,
            in3 => \N__27913\,
            lcout => \tok.uart_stall\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.valid_54_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__17749\,
            in1 => \N__22481\,
            in2 => \_gnd_net_\,
            in3 => \N__23308\,
            lcout => \tok.uart_rx_valid\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28537\,
            ce => \N__17732\,
            sr => \_gnd_net_\
        );

    \tok.uart.i1_2_lut_3_lut_4_lut_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__23307\,
            in1 => \N__25688\,
            in2 => \N__17750\,
            in3 => \N__22485\,
            lcout => \tok.uart.n953\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.T_7__I_0_233_i15_2_lut_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22479\,
            in2 => \_gnd_net_\,
            in3 => \N__23306\,
            lcout => \tok.n15_adj_667\,
            ltout => \tok.n15_adj_667_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_117_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__22303\,
            in1 => \N__24861\,
            in2 => \N__17723\,
            in3 => \N__27649\,
            lcout => \tok.n13_adj_780\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_171_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__30019\,
            in1 => \N__26975\,
            in2 => \N__17720\,
            in3 => \N__26762\,
            lcout => \tok.n11_adj_840\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_2_lut_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18358\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30018\,
            lcout => OPEN,
            ltout => \tok.n28_adj_771_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5446_4_lut_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__20270\,
            in1 => \N__19046\,
            in2 => \N__17690\,
            in3 => \N__18021\,
            lcout => OPEN,
            ltout => \tok.n5467_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i49_4_lut_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__19047\,
            in1 => \N__17687\,
            in2 => \N__17681\,
            in3 => \N__19244\,
            lcout => \tok.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2626_1_lut_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29119\,
            lcout => \tok.n82\,
            ltout => \tok.n82_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_2_lut_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24190\,
            in2 => \N__18425\,
            in3 => \N__20271\,
            lcout => \tok.n14_adj_764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2625_2_lut_3_lut_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__19738\,
            in1 => \N__18414\,
            in2 => \_gnd_net_\,
            in3 => \N__19045\,
            lcout => \tok.n2703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_178_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__19457\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17837\,
            lcout => \tok.n8_adj_846\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_80_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20229\,
            in2 => \_gnd_net_\,
            in3 => \N__18318\,
            lcout => \tok.n41\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \tok.n4761\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_3_lut_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18072\,
            in1 => \_gnd_net_\,
            in2 => \N__18353\,
            in3 => \N__18086\,
            lcout => \tok.n23_adj_718\,
            ltout => OPEN,
            carryin => \tok.n4761\,
            carryout => \tok.n4762\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_4_lut_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18074\,
            in1 => \N__30017\,
            in2 => \_gnd_net_\,
            in3 => \N__18077\,
            lcout => \tok.n15_adj_664\,
            ltout => OPEN,
            carryin => \tok.n4762\,
            carryout => \tok.n4763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_5_lut_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18073\,
            in1 => \N__18025\,
            in2 => \N__24219\,
            in3 => \N__17828\,
            lcout => \tok.n11_adj_830\,
            ltout => OPEN,
            carryin => \tok.n4763\,
            carryout => \tok.n4764\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_6_lut_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__27725\,
            in1 => \N__19052\,
            in2 => \_gnd_net_\,
            in3 => \N__17816\,
            lcout => \tok.n212\,
            ltout => OPEN,
            carryin => \tok.n4764\,
            carryout => \tok.n4765\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_7_lut_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21115\,
            in1 => \N__18804\,
            in2 => \_gnd_net_\,
            in3 => \N__18512\,
            lcout => \tok.n211\,
            ltout => OPEN,
            carryin => \tok.n4765\,
            carryout => \tok.n4766\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_8_lut_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__22750\,
            in1 => \N__19214\,
            in2 => \N__24209\,
            in3 => \N__18494\,
            lcout => \tok.n210\,
            ltout => OPEN,
            carryin => \tok.n4766\,
            carryout => \tok.n4767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_9_lut_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__29702\,
            in1 => \N__22110\,
            in2 => \N__24220\,
            in3 => \N__18491\,
            lcout => \tok.n209\,
            ltout => OPEN,
            carryin => \tok.n4767\,
            carryout => \tok.n4768\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_100_add_2_10_lut_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24189\,
            in2 => \_gnd_net_\,
            in3 => \N__18488\,
            lcout => \tok.n191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i105_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26408\,
            in1 => \N__18485\,
            in2 => \_gnd_net_\,
            in3 => \N__18451\,
            lcout => tail_105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28495\,
            ce => \N__26048\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i89_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18463\,
            in1 => \N__18442\,
            in2 => \_gnd_net_\,
            in3 => \N__26413\,
            lcout => \tok.A_stk.tail_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28495\,
            ce => \N__26048\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i73_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26412\,
            in1 => \N__18452\,
            in2 => \_gnd_net_\,
            in3 => \N__18433\,
            lcout => \tok.A_stk.tail_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28495\,
            ce => \N__26048\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i57_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18580\,
            in1 => \N__18443\,
            in2 => \_gnd_net_\,
            in3 => \N__26411\,
            lcout => \tok.A_stk.tail_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28495\,
            ce => \N__26048\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i41_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26410\,
            in1 => \N__18571\,
            in2 => \_gnd_net_\,
            in3 => \N__18434\,
            lcout => \tok.A_stk.tail_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28495\,
            ce => \N__26048\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i25_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__18581\,
            in1 => \_gnd_net_\,
            in2 => \N__18563\,
            in3 => \N__26409\,
            lcout => \tok.A_stk.tail_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28495\,
            ce => \N__26048\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i9_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26414\,
            in1 => \N__18572\,
            in2 => \_gnd_net_\,
            in3 => \N__27513\,
            lcout => \tok.A_stk.tail_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28495\,
            ce => \N__26048\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i9_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18559\,
            in1 => \N__25473\,
            in2 => \_gnd_net_\,
            in3 => \N__29081\,
            lcout => \tok.S_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28495\,
            ce => \N__26048\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i99_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26286\,
            in1 => \N__18550\,
            in2 => \_gnd_net_\,
            in3 => \N__20560\,
            lcout => tail_99,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28499\,
            ce => \N__26061\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i83_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26623\,
            in1 => \N__18535\,
            in2 => \_gnd_net_\,
            in3 => \N__26284\,
            lcout => \tok.A_stk.tail_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28499\,
            ce => \N__26061\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i20_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26280\,
            in1 => \N__18692\,
            in2 => \_gnd_net_\,
            in3 => \N__20548\,
            lcout => \tok.A_stk.tail_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28499\,
            ce => \N__26061\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i100_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20453\,
            in1 => \N__18523\,
            in2 => \_gnd_net_\,
            in3 => \N__26279\,
            lcout => tail_100,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28499\,
            ce => \N__26061\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i84_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26285\,
            in1 => \N__20464\,
            in2 => \_gnd_net_\,
            in3 => \N__18709\,
            lcout => \tok.A_stk.tail_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28499\,
            ce => \N__26061\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i68_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18524\,
            in1 => \N__18700\,
            in2 => \_gnd_net_\,
            in3 => \N__26283\,
            lcout => \tok.A_stk.tail_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28499\,
            ce => \N__26061\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i52_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26282\,
            in1 => \N__18691\,
            in2 => \_gnd_net_\,
            in3 => \N__18710\,
            lcout => \tok.A_stk.tail_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28499\,
            ce => \N__26061\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i36_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18664\,
            in1 => \N__18701\,
            in2 => \_gnd_net_\,
            in3 => \N__26281\,
            lcout => \tok.A_stk.tail_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28499\,
            ce => \N__26061\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i103_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18683\,
            in1 => \N__18628\,
            in2 => \_gnd_net_\,
            in3 => \N__26238\,
            lcout => tail_103,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28506\,
            ce => \N__25968\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i55_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26241\,
            in1 => \_gnd_net_\,
            in2 => \N__18641\,
            in3 => \N__20575\,
            lcout => \tok.A_stk.tail_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28506\,
            ce => \N__25968\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i71_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18629\,
            in1 => \N__20587\,
            in2 => \_gnd_net_\,
            in3 => \N__26242\,
            lcout => \tok.A_stk.tail_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28506\,
            ce => \N__25968\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i88_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26245\,
            in1 => \N__18592\,
            in2 => \_gnd_net_\,
            in3 => \N__20392\,
            lcout => \tok.A_stk.tail_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28506\,
            ce => \N__25968\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i4_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18665\,
            in1 => \N__26240\,
            in2 => \_gnd_net_\,
            in3 => \N__23742\,
            lcout => \tok.A_stk.tail_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28506\,
            ce => \N__25968\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i72_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26243\,
            in1 => \N__18605\,
            in2 => \_gnd_net_\,
            in3 => \N__21988\,
            lcout => \tok.A_stk.tail_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28506\,
            ce => \N__25968\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i87_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18652\,
            in1 => \N__18637\,
            in2 => \_gnd_net_\,
            in3 => \N__26244\,
            lcout => \tok.A_stk.tail_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28506\,
            ce => \N__25968\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i104_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26239\,
            in1 => \N__18617\,
            in2 => \_gnd_net_\,
            in3 => \N__18604\,
            lcout => tail_104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28506\,
            ce => \N__25968\,
            sr => \_gnd_net_\
        );

    \tok.i1_2_lut_adj_123_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18830\,
            in2 => \_gnd_net_\,
            in3 => \N__22141\,
            lcout => \tok.n9_adj_786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5447_4_lut_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110110"
        )
    port map (
            in0 => \N__22143\,
            in1 => \N__22760\,
            in2 => \N__19418\,
            in3 => \N__28978\,
            lcout => OPEN,
            ltout => \tok.n5548_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5445_4_lut_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__19307\,
            in1 => \N__23432\,
            in2 => \N__19283\,
            in3 => \N__26994\,
            lcout => \tok.n5547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i227_2_lut_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__18832\,
            in1 => \_gnd_net_\,
            in2 => \N__19073\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \tok.n285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_6_i1_4_lut_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101101"
        )
    port map (
            in0 => \N__19238\,
            in1 => \N__22759\,
            in2 => \N__19280\,
            in3 => \N__26763\,
            lcout => OPEN,
            ltout => \tok.n1_adj_862_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_199_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__19277\,
            in1 => \N__23213\,
            in2 => \N__19262\,
            in3 => \N__25771\,
            lcout => \tok.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i237_2_lut_3_lut_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__19237\,
            in1 => \N__19066\,
            in2 => \_gnd_net_\,
            in3 => \N__18831\,
            lcout => \tok.n6_adj_650\,
            ltout => \tok.n6_adj_650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i245_2_lut_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__22142\,
            in1 => \_gnd_net_\,
            in2 => \N__18713\,
            in3 => \_gnd_net_\,
            lcout => \tok.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_35_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__27652\,
            in1 => \N__20615\,
            in2 => \N__22313\,
            in3 => \N__27882\,
            lcout => OPEN,
            ltout => \tok.n13_adj_654_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5578_4_lut_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20351\,
            in1 => \N__20927\,
            in2 => \N__19391\,
            in3 => \N__19388\,
            lcout => OPEN,
            ltout => \tok.n5546_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i8_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011111000100"
        )
    port map (
            in0 => \N__26828\,
            in1 => \N__28589\,
            in2 => \N__19382\,
            in3 => \N__23543\,
            lcout => \A_low_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28518\,
            ce => \N__28300\,
            sr => \N__28205\
        );

    \tok.i2_4_lut_adj_195_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__21834\,
            in1 => \N__20624\,
            in2 => \N__27887\,
            in3 => \N__27651\,
            lcout => OPEN,
            ltout => \tok.n13_adj_641_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5582_4_lut_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19379\,
            in1 => \N__19367\,
            in2 => \N__19361\,
            in3 => \N__19358\,
            lcout => OPEN,
            ltout => \tok.n5551_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i7_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__28588\,
            in1 => \N__26827\,
            in2 => \N__19352\,
            in3 => \N__23633\,
            lcout => \tok.A_low_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28518\,
            ce => \N__28300\,
            sr => \N__28205\
        );

    \tok.add_104_2_lut_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27738\,
            in2 => \N__22880\,
            in3 => \N__19598\,
            lcout => \tok.n5465\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \tok.n4784\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_3_lut_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19595\,
            in1 => \N__21107\,
            in2 => \N__24035\,
            in3 => \N__19340\,
            lcout => \tok.n17_adj_812\,
            ltout => OPEN,
            carryin => \tok.n4784\,
            carryout => \tok.n4785\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_4_lut_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19591\,
            in1 => \N__22732\,
            in2 => \N__23920\,
            in3 => \N__19337\,
            lcout => \tok.n16_adj_810\,
            ltout => OPEN,
            carryin => \tok.n4785\,
            carryout => \tok.n4786\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_5_lut_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19594\,
            in1 => \N__29700\,
            in2 => \N__25373\,
            in3 => \N__19445\,
            lcout => \tok.n4_adj_806\,
            ltout => OPEN,
            carryin => \tok.n4786\,
            carryout => \tok.n4787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_6_lut_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19593\,
            in1 => \N__29585\,
            in2 => \N__23762\,
            in3 => \N__19436\,
            lcout => \tok.n5564\,
            ltout => OPEN,
            carryin => \tok.n4787\,
            carryout => \tok.n4788\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_7_lut_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19597\,
            in1 => \N__27303\,
            in2 => \N__27209\,
            in3 => \N__19433\,
            lcout => \tok.n5_adj_800\,
            ltout => OPEN,
            carryin => \tok.n4788\,
            carryout => \tok.n4789\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_8_lut_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19592\,
            in1 => \N__21830\,
            in2 => \N__23666\,
            in3 => \N__19421\,
            lcout => \tok.n5554\,
            ltout => OPEN,
            carryin => \tok.n4789\,
            carryout => \tok.n4790\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_9_lut_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19596\,
            in1 => \N__22258\,
            in2 => \N__23533\,
            in3 => \N__19406\,
            lcout => \tok.n5549\,
            ltout => OPEN,
            carryin => \tok.n4790\,
            carryout => \tok.n4791\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_10_lut_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19590\,
            in1 => \N__29447\,
            in2 => \N__28066\,
            in3 => \N__19403\,
            lcout => \tok.n5_adj_669\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \tok.n4792\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_11_lut_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19601\,
            in1 => \N__29061\,
            in2 => \N__27531\,
            in3 => \N__19400\,
            lcout => \tok.n25\,
            ltout => OPEN,
            carryin => \tok.n4792\,
            carryout => \tok.n4793\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_12_lut_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19587\,
            in1 => \N__29249\,
            in2 => \N__27459\,
            in3 => \N__19397\,
            lcout => \tok.n24_adj_703\,
            ltout => OPEN,
            carryin => \tok.n4793\,
            carryout => \tok.n4794\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_13_lut_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19599\,
            in1 => \N__25146\,
            in2 => \N__25059\,
            in3 => \N__19394\,
            lcout => \tok.n5_adj_726\,
            ltout => OPEN,
            carryin => \tok.n4794\,
            carryout => \tok.n4795\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_14_lut_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19586\,
            in1 => \N__21611\,
            in2 => \N__24477\,
            in3 => \N__19619\,
            lcout => \tok.n5_adj_734\,
            ltout => OPEN,
            carryin => \tok.n4795\,
            carryout => \tok.n4796\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_15_lut_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19600\,
            in1 => \N__23150\,
            in2 => \N__24369\,
            in3 => \N__19616\,
            lcout => \tok.n5_adj_732\,
            ltout => OPEN,
            carryin => \tok.n4796\,
            carryout => \tok.n4797\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_16_lut_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19589\,
            in1 => \N__28859\,
            in2 => \N__25772\,
            in3 => \N__19604\,
            lcout => \tok.n5_adj_716\,
            ltout => OPEN,
            carryin => \tok.n4797\,
            carryout => \tok.n4798\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_104_17_lut_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__24860\,
            in1 => \N__19588\,
            in2 => \N__24778\,
            in3 => \N__19526\,
            lcout => \tok.n5_adj_713\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5561_4_lut_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__22340\,
            in1 => \N__19523\,
            in2 => \N__20882\,
            in3 => \N__21011\,
            lcout => \tok.n5574\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5242_4_lut_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26940\,
            in1 => \N__21910\,
            in2 => \N__27878\,
            in3 => \N__19510\,
            lcout => OPEN,
            ltout => \tok.n5414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_149_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001111"
        )
    port map (
            in0 => \N__22528\,
            in1 => \N__19499\,
            in2 => \N__19487\,
            in3 => \N__19484\,
            lcout => \tok.n904\,
            ltout => \tok.n904_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i47_3_lut_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27855\,
            in1 => \_gnd_net_\,
            in2 => \N__19478\,
            in3 => \N__22710\,
            lcout => OPEN,
            ltout => \tok.n5346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_172_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001111"
        )
    port map (
            in0 => \N__22529\,
            in1 => \N__19475\,
            in2 => \N__19460\,
            in3 => \N__23225\,
            lcout => OPEN,
            ltout => \tok.n14_adj_841_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5557_4_lut_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__19790\,
            in1 => \N__29750\,
            in2 => \N__19775\,
            in3 => \N__19772\,
            lcout => \tok.n5569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i49_3_lut_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29687\,
            in1 => \N__27854\,
            in2 => \_gnd_net_\,
            in3 => \N__27629\,
            lcout => \tok.n45_adj_849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i3_1_lut_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22709\,
            lcout => \tok.n300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_57_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__29345\,
            in1 => \N__21875\,
            in2 => \_gnd_net_\,
            in3 => \N__19745\,
            lcout => \tok.n45_adj_696\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_50_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101111"
        )
    port map (
            in0 => \N__27325\,
            in1 => \N__19706\,
            in2 => \N__21314\,
            in3 => \N__26751\,
            lcout => \tok.n10_adj_686\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__29344\,
            in1 => \N__27324\,
            in2 => \_gnd_net_\,
            in3 => \N__19744\,
            lcout => OPEN,
            ltout => \tok.n45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_46_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110010"
        )
    port map (
            in0 => \N__19724\,
            in1 => \N__19642\,
            in2 => \N__19709\,
            in3 => \N__19699\,
            lcout => \tok.n39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_58_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000100"
        )
    port map (
            in0 => \N__19700\,
            in1 => \N__19667\,
            in2 => \N__19646\,
            in3 => \N__19634\,
            lcout => OPEN,
            ltout => \tok.n39_adj_697_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_60_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__21876\,
            in1 => \N__21311\,
            in2 => \N__19628\,
            in3 => \N__26752\,
            lcout => OPEN,
            ltout => \tok.n10_adj_700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5441_4_lut_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__27371\,
            in1 => \N__22616\,
            in2 => \N__19922\,
            in3 => \N__20852\,
            lcout => \tok.n5536\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_180_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000111011"
        )
    port map (
            in0 => \N__22882\,
            in1 => \N__20296\,
            in2 => \N__28789\,
            in3 => \N__28939\,
            lcout => \tok.n11_adj_730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_66_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27327\,
            in1 => \N__23111\,
            in2 => \N__29470\,
            in3 => \N__29701\,
            lcout => OPEN,
            ltout => \tok.n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i15_4_lut_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19805\,
            in1 => \N__19796\,
            in2 => \N__19907\,
            in3 => \N__19811\,
            lcout => \tok.tc__7__N_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27690\,
            in1 => \N__29552\,
            in2 => \N__21108\,
            in3 => \N__21865\,
            lcout => \tok.n25_adj_710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i12_4_lut_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29038\,
            in1 => \N__25767\,
            in2 => \N__24844\,
            in3 => \N__25116\,
            lcout => \tok.n28_adj_708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i11_4_lut_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22268\,
            in1 => \N__29215\,
            in2 => \N__22731\,
            in3 => \N__21595\,
            lcout => \tok.n27_adj_709\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_94_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001011101"
        )
    port map (
            in0 => \N__23112\,
            in1 => \N__29464\,
            in2 => \N__28979\,
            in3 => \N__27876\,
            lcout => \tok.n12_adj_745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_74_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__27874\,
            in1 => \N__28972\,
            in2 => \N__25145\,
            in3 => \N__21866\,
            lcout => \tok.n12_adj_723\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_116_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001111"
        )
    port map (
            in0 => \N__28973\,
            in1 => \N__29240\,
            in2 => \N__24845\,
            in3 => \N__27875\,
            lcout => \tok.n12_adj_779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_191_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__26747\,
            in1 => \N__20321\,
            in2 => \_gnd_net_\,
            in3 => \N__20272\,
            lcout => \tok.n10_adj_858\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_adj_97_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__26984\,
            in1 => \N__20003\,
            in2 => \_gnd_net_\,
            in3 => \N__19988\,
            lcout => \tok.n16_adj_749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_114_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001101"
        )
    port map (
            in0 => \N__26748\,
            in1 => \N__20342\,
            in2 => \N__21313\,
            in3 => \N__25167\,
            lcout => OPEN,
            ltout => \tok.n14_adj_776_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_120_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24071\,
            in1 => \N__19979\,
            in2 => \N__19973\,
            in3 => \N__19970\,
            lcout => OPEN,
            ltout => \tok.n20_adj_784_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5572_4_lut_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20699\,
            in1 => \N__19928\,
            in2 => \N__19964\,
            in3 => \N__19961\,
            lcout => \tok.n5513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_15_i9_2_lut_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24767\,
            in2 => \_gnd_net_\,
            in3 => \N__28777\,
            lcout => \tok.n9_adj_781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_adj_118_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__19955\,
            in1 => \N__19946\,
            in2 => \_gnd_net_\,
            in3 => \N__26983\,
            lcout => \tok.n16_adj_782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_4_lut_adj_182_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__28781\,
            in1 => \N__20357\,
            in2 => \N__23554\,
            in3 => \N__29139\,
            lcout => \tok.n14_adj_658\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_11_i2_3_lut_3_lut_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__29310\,
            in1 => \N__29138\,
            in2 => \_gnd_net_\,
            in3 => \N__22269\,
            lcout => \tok.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_15_i2_3_lut_3_lut_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__29319\,
            in1 => \N__29160\,
            in2 => \_gnd_net_\,
            in3 => \N__25166\,
            lcout => \tok.n2_adj_775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i102_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20333\,
            in1 => \N__20603\,
            in2 => \_gnd_net_\,
            in3 => \N__26526\,
            lcout => tail_102,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28500\,
            ce => \N__26049\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i125_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__21443\,
            in1 => \N__26011\,
            in2 => \N__21460\,
            in3 => \N__26455\,
            lcout => tail_125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i123_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__26453\,
            in1 => \N__21557\,
            in2 => \N__26055\,
            in3 => \N__21361\,
            lcout => tail_123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i124_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__21509\,
            in1 => \N__26010\,
            in2 => \N__21530\,
            in3 => \N__26454\,
            lcout => tail_124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i118_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__26451\,
            in1 => \N__20332\,
            in2 => \N__26054\,
            in3 => \N__20380\,
            lcout => tail_118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i122_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__25211\,
            in1 => \N__26006\,
            in2 => \N__25228\,
            in3 => \N__26452\,
            lcout => tail_122,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i116_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__26450\,
            in1 => \N__20468\,
            in2 => \N__26053\,
            in3 => \N__20449\,
            lcout => tail_116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i114_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__20419\,
            in1 => \N__25999\,
            in2 => \N__20437\,
            in3 => \N__26449\,
            lcout => tail_114,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i23_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20576\,
            in1 => \N__21745\,
            in2 => \_gnd_net_\,
            in3 => \N__26343\,
            lcout => \tok.A_stk.tail_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28512\,
            ce => \N__26031\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i70_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26347\,
            in1 => \N__20602\,
            in2 => \_gnd_net_\,
            in3 => \N__20524\,
            lcout => \tok.A_stk.tail_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28512\,
            ce => \N__26031\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i98_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20438\,
            in1 => \N__20401\,
            in2 => \_gnd_net_\,
            in3 => \N__26350\,
            lcout => tail_98,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28512\,
            ce => \N__26031\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i66_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26346\,
            in1 => \_gnd_net_\,
            in2 => \N__20405\,
            in3 => \N__21692\,
            lcout => \tok.A_stk.tail_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28512\,
            ce => \N__26031\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i82_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20420\,
            in1 => \N__21703\,
            in2 => \_gnd_net_\,
            in3 => \N__26348\,
            lcout => \tok.A_stk.tail_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28512\,
            ce => \N__26031\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i56_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26345\,
            in1 => \N__21977\,
            in2 => \_gnd_net_\,
            in3 => \N__20393\,
            lcout => \tok.A_stk.tail_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28512\,
            ce => \N__26031\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i54_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20366\,
            in1 => \N__20500\,
            in2 => \_gnd_net_\,
            in3 => \N__26344\,
            lcout => \tok.A_stk.tail_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28512\,
            ce => \N__26031\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i86_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26349\,
            in1 => \N__20381\,
            in2 => \_gnd_net_\,
            in3 => \N__20365\,
            lcout => \tok.A_stk.tail_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28512\,
            ce => \N__26031\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i39_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26508\,
            in1 => \N__20488\,
            in2 => \_gnd_net_\,
            in3 => \N__20588\,
            lcout => \tok.A_stk.tail_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28519\,
            ce => \N__26021\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i67_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26096\,
            in1 => \N__20564\,
            in2 => \_gnd_net_\,
            in3 => \N__26509\,
            lcout => \tok.A_stk.tail_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28519\,
            ce => \N__26021\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i4_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20549\,
            in1 => \N__25498\,
            in2 => \_gnd_net_\,
            in3 => \N__29599\,
            lcout => \tok.S_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28519\,
            ce => \N__26021\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i6_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25499\,
            in1 => \N__20536\,
            in2 => \_gnd_net_\,
            in3 => \N__21835\,
            lcout => \tok.S_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28519\,
            ce => \N__26021\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i6_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26510\,
            in1 => \N__20513\,
            in2 => \_gnd_net_\,
            in3 => \N__23648\,
            lcout => \tok.A_stk.tail_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28519\,
            ce => \N__26021\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i22_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20504\,
            in1 => \N__20537\,
            in2 => \_gnd_net_\,
            in3 => \N__26506\,
            lcout => \tok.A_stk.tail_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28519\,
            ce => \N__26021\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i38_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26507\,
            in1 => \_gnd_net_\,
            in2 => \N__20528\,
            in3 => \N__20512\,
            lcout => \tok.A_stk.tail_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28519\,
            ce => \N__26021\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23523\,
            in1 => \N__20489\,
            in2 => \_gnd_net_\,
            in3 => \N__26511\,
            lcout => \tok.A_stk.tail_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28519\,
            ce => \N__26021\,
            sr => \_gnd_net_\
        );

    \tok.add_109_2_lut_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20843\,
            in1 => \N__22881\,
            in2 => \_gnd_net_\,
            in3 => \N__20666\,
            lcout => \tok.n3_adj_692\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \tok.n4799\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_3_lut_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20839\,
            in1 => \N__24029\,
            in2 => \_gnd_net_\,
            in3 => \N__20663\,
            lcout => \tok.n14_adj_662\,
            ltout => OPEN,
            carryin => \tok.n4799\,
            carryout => \tok.n4800\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_4_lut_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20842\,
            in1 => \N__23913\,
            in2 => \_gnd_net_\,
            in3 => \N__20660\,
            lcout => \tok.n12_adj_832\,
            ltout => OPEN,
            carryin => \tok.n4800\,
            carryout => \tok.n4801\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_5_lut_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20838\,
            in1 => \N__25335\,
            in2 => \_gnd_net_\,
            in3 => \N__20645\,
            lcout => \tok.n22_adj_829\,
            ltout => OPEN,
            carryin => \tok.n4801\,
            carryout => \tok.n4802\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_6_lut_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20765\,
            in1 => \N__23732\,
            in2 => \_gnd_net_\,
            in3 => \N__20630\,
            lcout => \tok.n10_adj_827\,
            ltout => OPEN,
            carryin => \tok.n4802\,
            carryout => \tok.n4803\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_7_lut_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20767\,
            in1 => \N__27188\,
            in2 => \_gnd_net_\,
            in3 => \N__20627\,
            lcout => \tok.n10_adj_823\,
            ltout => OPEN,
            carryin => \tok.n4803\,
            carryout => \tok.n4804\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_8_lut_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20766\,
            in1 => \N__23629\,
            in2 => \_gnd_net_\,
            in3 => \N__20618\,
            lcout => \tok.n10_adj_820\,
            ltout => OPEN,
            carryin => \tok.n4804\,
            carryout => \tok.n4805\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_9_lut_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20768\,
            in1 => \N__23519\,
            in2 => \_gnd_net_\,
            in3 => \N__20609\,
            lcout => \tok.n10_adj_653\,
            ltout => OPEN,
            carryin => \tok.n4805\,
            carryout => \tok.n4806\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_10_lut_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20750\,
            in1 => \N__28057\,
            in2 => \_gnd_net_\,
            in3 => \N__20606\,
            lcout => \tok.n10_adj_666\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \tok.n4807\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_11_lut_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20841\,
            in1 => \N__27539\,
            in2 => \_gnd_net_\,
            in3 => \N__20846\,
            lcout => \tok.n23_adj_682\,
            ltout => OPEN,
            carryin => \tok.n4807\,
            carryout => \tok.n4808\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_12_lut_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20840\,
            in1 => \N__27441\,
            in2 => \_gnd_net_\,
            in3 => \N__20804\,
            lcout => \tok.n22_adj_698\,
            ltout => OPEN,
            carryin => \tok.n4808\,
            carryout => \tok.n4809\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_13_lut_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20762\,
            in1 => \N__25054\,
            in2 => \_gnd_net_\,
            in3 => \N__20801\,
            lcout => \tok.n5534\,
            ltout => OPEN,
            carryin => \tok.n4809\,
            carryout => \tok.n4810\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_14_lut_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20748\,
            in1 => \N__24464\,
            in2 => \_gnd_net_\,
            in3 => \N__20789\,
            lcout => \tok.n10_adj_738\,
            ltout => OPEN,
            carryin => \tok.n4810\,
            carryout => \tok.n4811\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_15_lut_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20763\,
            in1 => \N__24365\,
            in2 => \_gnd_net_\,
            in3 => \N__20786\,
            lcout => \tok.n5525\,
            ltout => OPEN,
            carryin => \tok.n4811\,
            carryout => \tok.n4812\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_16_lut_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20749\,
            in1 => \N__28866\,
            in2 => \_gnd_net_\,
            in3 => \N__20771\,
            lcout => \tok.n10_adj_768\,
            ltout => OPEN,
            carryin => \tok.n4812\,
            carryout => \tok.n4813\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.add_109_17_lut_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__24777\,
            in1 => \N__20751\,
            in2 => \_gnd_net_\,
            in3 => \N__20702\,
            lcout => \tok.n5516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_90_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__21612\,
            in1 => \N__26760\,
            in2 => \N__20900\,
            in3 => \N__27624\,
            lcout => OPEN,
            ltout => \tok.n12_adj_737_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_92_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__20684\,
            in1 => \N__22322\,
            in2 => \N__20669\,
            in3 => \N__28970\,
            lcout => \tok.n20_adj_740\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_7_i1_4_lut_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001000101"
        )
    port map (
            in0 => \N__26761\,
            in1 => \N__29728\,
            in2 => \N__22187\,
            in3 => \N__22146\,
            lcout => OPEN,
            ltout => \tok.n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_36_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__23208\,
            in1 => \N__20915\,
            in2 => \N__20930\,
            in3 => \N__24843\,
            lcout => \tok.n17_adj_656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_7_i12_2_lut_3_lut_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__20908\,
            in1 => \N__22548\,
            in2 => \_gnd_net_\,
            in3 => \N__23332\,
            lcout => \tok.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i7_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23008\,
            in1 => \N__25692\,
            in2 => \_gnd_net_\,
            in3 => \N__20909\,
            lcout => uart_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_99_i13_2_lut_3_lut_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__22182\,
            in1 => \N__29448\,
            in2 => \_gnd_net_\,
            in3 => \N__22145\,
            lcout => \tok.n177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_168_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__20891\,
            in1 => \N__28758\,
            in2 => \_gnd_net_\,
            in3 => \N__24039\,
            lcout => \tok.n9_adj_838\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_47_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__20873\,
            in1 => \N__21135\,
            in2 => \_gnd_net_\,
            in3 => \N__23336\,
            lcout => OPEN,
            ltout => \tok.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_53_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111110"
        )
    port map (
            in0 => \N__20861\,
            in1 => \N__24608\,
            in2 => \N__20855\,
            in3 => \N__22549\,
            lcout => \tok.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i59_3_lut_adj_63_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29270\,
            in1 => \N__27857\,
            in2 => \_gnd_net_\,
            in3 => \N__27631\,
            lcout => \tok.n5350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i1_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21188\,
            in1 => \N__25694\,
            in2 => \_gnd_net_\,
            in3 => \N__22600\,
            lcout => uart_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i59_3_lut_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29079\,
            in1 => \N__27858\,
            in2 => \_gnd_net_\,
            in3 => \N__27632\,
            lcout => OPEN,
            ltout => \tok.n5342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5560_4_lut_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__27476\,
            in1 => \N__21158\,
            in2 => \N__21152\,
            in3 => \N__21149\,
            lcout => \tok.n5539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i44_3_lut_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21136\,
            in1 => \N__27856\,
            in2 => \_gnd_net_\,
            in3 => \N__27630\,
            lcout => \tok.n5336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_11_i9_2_lut_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28782\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25055\,
            lcout => \tok.n9_adj_725\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_3_lut_adj_76_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__21005\,
            in1 => \N__20987\,
            in2 => \_gnd_net_\,
            in3 => \N__26993\,
            lcout => \tok.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_75_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__25157\,
            in1 => \N__29704\,
            in2 => \N__27953\,
            in3 => \N__27625\,
            lcout => OPEN,
            ltout => \tok.n13_adj_724_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_78_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24509\,
            in1 => \N__21230\,
            in2 => \N__20975\,
            in3 => \N__20972\,
            lcout => OPEN,
            ltout => \tok.n20_adj_729_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5567_4_lut_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20966\,
            in1 => \N__20957\,
            in2 => \N__20951\,
            in3 => \N__20948\,
            lcout => \tok.n5531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_73_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101111"
        )
    port map (
            in0 => \N__21239\,
            in1 => \N__22299\,
            in2 => \N__21312\,
            in3 => \N__26749\,
            lcout => \tok.n14_adj_722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i11_1_lut_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29253\,
            lcout => \tok.n292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i12_1_lut_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25156\,
            lcout => \tok.n291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5583_4_lut_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__24404\,
            in1 => \N__21248\,
            in2 => \N__21197\,
            in3 => \N__21224\,
            lcout => OPEN,
            ltout => \tok.n5527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i13_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011101110"
        )
    port map (
            in0 => \N__28652\,
            in1 => \N__24480\,
            in2 => \N__21215\,
            in3 => \N__26855\,
            lcout => \tok.A_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28542\,
            ce => \N__28296\,
            sr => \N__28230\
        );

    \tok.A_i14_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__26856\,
            in1 => \N__28653\,
            in2 => \N__24374\,
            in3 => \N__21320\,
            lcout => \tok.A_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28542\,
            ce => \N__28296\,
            sr => \N__28230\
        );

    \tok.A_i16_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__24746\,
            in1 => \N__26857\,
            in2 => \N__28658\,
            in3 => \N__21212\,
            lcout => \tok.A_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28542\,
            ce => \N__28296\,
            sr => \N__28230\
        );

    \tok.A_i10_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__27550\,
            in1 => \N__26854\,
            in2 => \N__28657\,
            in3 => \N__21206\,
            lcout => \tok.A_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28542\,
            ce => \N__28296\,
            sr => \N__28230\
        );

    \tok.i5181_2_lut_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27877\,
            in2 => \_gnd_net_\,
            in3 => \N__21599\,
            lcout => \tok.n5348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_4_lut_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__27549\,
            in1 => \N__24825\,
            in2 => \N__24760\,
            in3 => \N__29039\,
            lcout => \tok.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_95_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__27343\,
            in1 => \N__23116\,
            in2 => \N__27959\,
            in3 => \N__27650\,
            lcout => OPEN,
            ltout => \tok.n13_adj_746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i9_4_lut_adj_99_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24278\,
            in1 => \N__21269\,
            in2 => \N__21350\,
            in3 => \N__21347\,
            lcout => OPEN,
            ltout => \tok.n20_adj_753_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5581_4_lut_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21341\,
            in1 => \N__21329\,
            in2 => \N__21323\,
            in3 => \N__21263\,
            lcout => \tok.n5522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_93_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111011"
        )
    port map (
            in0 => \N__21257\,
            in1 => \N__21304\,
            in2 => \N__29065\,
            in3 => \N__26750\,
            lcout => \tok.n14_adj_744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_13_i9_2_lut_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24370\,
            in2 => \_gnd_net_\,
            in3 => \N__28783\,
            lcout => \tok.n9_adj_748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.select_73_Select_13_i2_3_lut_3_lut_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__29343\,
            in1 => \N__29153\,
            in2 => \_gnd_net_\,
            in3 => \N__29040\,
            lcout => \tok.n2_adj_743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_101_i13_2_lut_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29349\,
            in2 => \_gnd_net_\,
            in3 => \N__29460\,
            lcout => OPEN,
            ltout => \tok.n204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5_4_lut_4_lut_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__29171\,
            in1 => \N__24479\,
            in2 => \N__21251\,
            in3 => \N__28790\,
            lcout => \tok.n16_adj_741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i109_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21467\,
            in1 => \N__21424\,
            in2 => \_gnd_net_\,
            in3 => \N__26574\,
            lcout => tail_109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28508\,
            ce => \N__26073\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i93_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26580\,
            in1 => \N__21436\,
            in2 => \_gnd_net_\,
            in3 => \N__21412\,
            lcout => \tok.A_stk.tail_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28508\,
            ce => \N__26073\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i77_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21425\,
            in1 => \N__21403\,
            in2 => \_gnd_net_\,
            in3 => \N__26579\,
            lcout => \tok.A_stk.tail_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28508\,
            ce => \N__26073\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i61_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26578\,
            in1 => \N__21394\,
            in2 => \_gnd_net_\,
            in3 => \N__21413\,
            lcout => \tok.A_stk.tail_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28508\,
            ce => \N__26073\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i45_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21385\,
            in1 => \N__21404\,
            in2 => \_gnd_net_\,
            in3 => \N__26577\,
            lcout => \tok.A_stk.tail_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28508\,
            ce => \N__26073\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i29_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__26576\,
            in1 => \_gnd_net_\,
            in2 => \N__21377\,
            in3 => \N__21395\,
            lcout => \tok.A_stk.tail_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28508\,
            ce => \N__26073\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i13_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21386\,
            in1 => \N__26575\,
            in2 => \_gnd_net_\,
            in3 => \N__24319\,
            lcout => \tok.A_stk.tail_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28508\,
            ce => \N__26073\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i13_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21373\,
            in1 => \N__25512\,
            in2 => \_gnd_net_\,
            in3 => \N__23162\,
            lcout => \tok.S_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28508\,
            ce => \N__26073\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i107_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21365\,
            in1 => \N__21541\,
            in2 => \_gnd_net_\,
            in3 => \N__26560\,
            lcout => tail_107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28513\,
            ce => \N__26058\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i91_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26566\,
            in1 => \N__21553\,
            in2 => \_gnd_net_\,
            in3 => \N__25564\,
            lcout => \tok.A_stk.tail_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28513\,
            ce => \N__26058\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i75_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21542\,
            in1 => \N__25553\,
            in2 => \_gnd_net_\,
            in3 => \N__26564\,
            lcout => \tok.A_stk.tail_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28513\,
            ce => \N__26058\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i108_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26561\,
            in1 => \N__21529\,
            in2 => \_gnd_net_\,
            in3 => \N__21493\,
            lcout => tail_108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28513\,
            ce => \N__26058\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i92_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21505\,
            in1 => \N__21484\,
            in2 => \_gnd_net_\,
            in3 => \N__26567\,
            lcout => \tok.A_stk.tail_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28513\,
            ce => \N__26058\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i76_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26565\,
            in1 => \N__21494\,
            in2 => \_gnd_net_\,
            in3 => \N__21475\,
            lcout => \tok.A_stk.tail_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28513\,
            ce => \N__26058\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i60_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21673\,
            in1 => \N__21485\,
            in2 => \_gnd_net_\,
            in3 => \N__26563\,
            lcout => \tok.A_stk.tail_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28513\,
            ce => \N__26058\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i44_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26562\,
            in1 => \N__21662\,
            in2 => \_gnd_net_\,
            in3 => \N__21476\,
            lcout => \tok.A_stk.tail_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28513\,
            ce => \N__26058\,
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23880\,
            in1 => \N__22311\,
            in2 => \N__23507\,
            in3 => \N__22762\,
            lcout => \tok.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i2_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21733\,
            in1 => \N__25450\,
            in2 => \_gnd_net_\,
            in3 => \N__22763\,
            lcout => \tok.S_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28520\,
            ce => \N__26035\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i7_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22312\,
            in1 => \N__21752\,
            in2 => \_gnd_net_\,
            in3 => \N__25451\,
            lcout => \tok.S_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28520\,
            ce => \N__26035\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i2_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23881\,
            in1 => \_gnd_net_\,
            in2 => \N__26582\,
            in3 => \N__21725\,
            lcout => \tok.A_stk.tail_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28520\,
            ce => \N__26035\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i18_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21716\,
            in1 => \N__21734\,
            in2 => \_gnd_net_\,
            in3 => \N__26512\,
            lcout => \tok.A_stk.tail_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28520\,
            ce => \N__26035\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i34_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26516\,
            in1 => \N__21724\,
            in2 => \_gnd_net_\,
            in3 => \N__21691\,
            lcout => \tok.A_stk.tail_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28520\,
            ce => \N__26035\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i50_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21715\,
            in1 => \N__21707\,
            in2 => \_gnd_net_\,
            in3 => \N__26517\,
            lcout => \tok.A_stk.tail_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28520\,
            ce => \N__26035\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i12_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21661\,
            in1 => \N__26527\,
            in2 => \_gnd_net_\,
            in3 => \N__24457\,
            lcout => \tok.A_stk.tail_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28525\,
            ce => \N__26059\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i28_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__26529\,
            in1 => \_gnd_net_\,
            in2 => \N__21647\,
            in3 => \N__21677\,
            lcout => \tok.A_stk.tail_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28525\,
            ce => \N__26059\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i12_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21635\,
            in1 => \N__21643\,
            in2 => \_gnd_net_\,
            in3 => \N__25500\,
            lcout => \tok.S_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28525\,
            ce => \N__26059\,
            sr => \_gnd_net_\
        );

    \tok.inv_106_i13_1_lut_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21634\,
            lcout => \tok.n290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i8_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29452\,
            in1 => \N__22018\,
            in2 => \_gnd_net_\,
            in3 => \N__25501\,
            lcout => \tok.S_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28525\,
            ce => \N__26059\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i8_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26531\,
            in1 => \_gnd_net_\,
            in2 => \N__22010\,
            in3 => \N__28035\,
            lcout => \tok.A_stk.tail_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28525\,
            ce => \N__26059\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i24_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21973\,
            in1 => \N__22019\,
            in2 => \_gnd_net_\,
            in3 => \N__26528\,
            lcout => \tok.A_stk.tail_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28525\,
            ce => \N__26059\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i40_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__26530\,
            in1 => \_gnd_net_\,
            in2 => \N__22009\,
            in3 => \N__21995\,
            lcout => \tok.A_stk.tail_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28525\,
            ce => \N__26059\,
            sr => \_gnd_net_\
        );

    \tok.i14_4_lut_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21959\,
            in1 => \N__25190\,
            in2 => \N__21950\,
            in3 => \N__21932\,
            lcout => OPEN,
            ltout => \tok.n30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5151_3_lut_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21758\,
            in2 => \N__21917\,
            in3 => \N__21914\,
            lcout => \tok.n4908\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__28028\,
            in1 => \N__29459\,
            in2 => \N__24341\,
            in3 => \N__23158\,
            lcout => \tok.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_38_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__22872\,
            in1 => \N__21864\,
            in2 => \N__23677\,
            in3 => \N__27774\,
            lcout => OPEN,
            ltout => \tok.n17_adj_661_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i13_4_lut_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25535\,
            in1 => \N__21782\,
            in2 => \N__21767\,
            in3 => \N__21764\,
            lcout => \tok.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_163_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__23951\,
            in1 => \N__29075\,
            in2 => \_gnd_net_\,
            in3 => \N__23406\,
            lcout => \tok.n6_adj_834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_59_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__22764\,
            in1 => \N__22646\,
            in2 => \_gnd_net_\,
            in3 => \N__23331\,
            lcout => OPEN,
            ltout => \tok.n4_adj_699_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_4_lut_adj_62_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111110"
        )
    port map (
            in0 => \N__24536\,
            in1 => \N__22634\,
            in2 => \N__22619\,
            in3 => \N__22544\,
            lcout => \tok.n9_adj_705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_3_lut_adj_164_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__22604\,
            in1 => \N__22586\,
            in2 => \_gnd_net_\,
            in3 => \N__23330\,
            lcout => OPEN,
            ltout => \tok.n5_adj_835_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_165_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111110"
        )
    port map (
            in0 => \N__22574\,
            in1 => \N__22568\,
            in2 => \N__22553\,
            in3 => \N__22543\,
            lcout => \tok.n10_adj_836\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i8_1_lut_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22310\,
            lcout => \tok.n295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i10_1_lut_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29074\,
            lcout => \tok.n293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_99_i15_2_lut_3_lut_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__29269\,
            in1 => \N__22186\,
            in2 => \_gnd_net_\,
            in3 => \N__22151\,
            lcout => \tok.n175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_inv_0_i1_1_lut_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27766\,
            lcout => \tok.n17_adj_711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_169_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__23825\,
            in1 => \N__29271\,
            in2 => \_gnd_net_\,
            in3 => \N__23411\,
            lcout => OPEN,
            ltout => \tok.n6_adj_839_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_4_lut_adj_170_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__23366\,
            in1 => \N__23351\,
            in2 => \N__23339\,
            in3 => \N__23333\,
            lcout => \tok.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5550_2_lut_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__23204\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23155\,
            lcout => \tok.n5559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_4_lut_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__23069\,
            in1 => \N__29178\,
            in2 => \N__23054\,
            in3 => \N__26765\,
            lcout => \tok.n16_adj_855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i6_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22906\,
            in1 => \_gnd_net_\,
            in2 => \N__25615\,
            in3 => \N__22971\,
            lcout => capture_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i5_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22970\,
            in1 => \N__23023\,
            in2 => \_gnd_net_\,
            in3 => \N__25611\,
            lcout => capture_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.capture_i0_i7_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22905\,
            in1 => \N__23012\,
            in2 => \_gnd_net_\,
            in3 => \N__22972\,
            lcout => capture_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_2_lut_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24592\,
            in1 => \N__22892\,
            in2 => \N__22871\,
            in3 => \N__22769\,
            lcout => \tok.n11_adj_809\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \tok.n4769\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_3_lut_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24588\,
            in1 => \N__24059\,
            in2 => \N__24043\,
            in3 => \N__23942\,
            lcout => \tok.n20_adj_799\,
            ltout => OPEN,
            carryin => \tok.n4769\,
            carryout => \tok.n4770\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_4_lut_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24591\,
            in1 => \N__23906\,
            in2 => \N__23840\,
            in3 => \N__23816\,
            lcout => \tok.n22_adj_797\,
            ltout => OPEN,
            carryin => \tok.n4770\,
            carryout => \tok.n4771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_5_lut_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24589\,
            in1 => \N__25339\,
            in2 => \N__25529\,
            in3 => \N__23798\,
            lcout => \tok.n10_adj_791\,
            ltout => OPEN,
            carryin => \tok.n4771\,
            carryout => \tok.n4772\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_6_lut_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24141\,
            in1 => \N__23775\,
            in2 => \N__27362\,
            in3 => \N__23684\,
            lcout => \tok.n6_adj_762\,
            ltout => OPEN,
            carryin => \tok.n4772\,
            carryout => \tok.n4773\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_7_lut_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24135\,
            in1 => \N__27227\,
            in2 => \N__27214\,
            in3 => \N__23681\,
            lcout => \tok.n6_adj_717\,
            ltout => OPEN,
            carryin => \tok.n4773\,
            carryout => \tok.n4774\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_8_lut_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24142\,
            in1 => \N__23664\,
            in2 => \N__23588\,
            in3 => \N__23561\,
            lcout => \tok.n6\,
            ltout => OPEN,
            carryin => \tok.n4774\,
            carryout => \tok.n4775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_9_lut_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24134\,
            in1 => \N__23506\,
            in2 => \N__23444\,
            in3 => \N__23417\,
            lcout => \tok.n6_adj_657\,
            ltout => OPEN,
            carryin => \tok.n4775\,
            carryout => \tok.n4776\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_10_lut_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24139\,
            in1 => \N__29360\,
            in2 => \N__28067\,
            in3 => \N__23414\,
            lcout => \tok.n5544\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \tok.n4777\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_11_lut_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24590\,
            in1 => \N__27545\,
            in2 => \N__24620\,
            in3 => \N__24596\,
            lcout => \tok.n28\,
            ltout => OPEN,
            carryin => \tok.n4777\,
            carryout => \tok.n4778\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_12_lut_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24593\,
            in1 => \N__27440\,
            in2 => \N__24548\,
            in3 => \N__24527\,
            lcout => \tok.n27_adj_704\,
            ltout => OPEN,
            carryin => \tok.n4778\,
            carryout => \tok.n4779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_13_lut_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24136\,
            in1 => \N__25041\,
            in2 => \N__24524\,
            in3 => \N__24500\,
            lcout => \tok.n6_adj_728\,
            ltout => OPEN,
            carryin => \tok.n4779\,
            carryout => \tok.n4780\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_14_lut_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24140\,
            in1 => \N__24497\,
            in2 => \N__24478\,
            in3 => \N__24392\,
            lcout => \tok.n6_adj_742\,
            ltout => OPEN,
            carryin => \tok.n4780\,
            carryout => \tok.n4781\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_15_lut_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24137\,
            in1 => \N__24389\,
            in2 => \N__24364\,
            in3 => \N__24266\,
            lcout => \tok.n6_adj_752\,
            ltout => OPEN,
            carryin => \tok.n4781\,
            carryout => \tok.n4782\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_16_lut_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__24138\,
            in1 => \N__28857\,
            in2 => \N__25184\,
            in3 => \N__24263\,
            lcout => \tok.n5520\,
            ltout => OPEN,
            carryin => \tok.n4782\,
            carryout => \tok.n4783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_16_THRU_CRY_0_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24226\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \tok.n4783\,
            carryout => \tok.n4783_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.sub_105_add_2_17_lut_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__24758\,
            in1 => \N__24143\,
            in2 => \N__24872\,
            in3 => \N__24074\,
            lcout => \tok.n6_adj_783\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i16_1_lut_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24846\,
            lcout => \tok.n287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i15_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24847\,
            in1 => \N__24703\,
            in2 => \_gnd_net_\,
            in3 => \N__25514\,
            lcout => \tok.S_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28544\,
            ce => \N__26078\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i15_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24695\,
            in1 => \N__26602\,
            in2 => \_gnd_net_\,
            in3 => \N__24759\,
            lcout => \tok.A_stk.tail_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28544\,
            ce => \N__26078\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i31_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26603\,
            in1 => \N__24704\,
            in2 => \_gnd_net_\,
            in3 => \N__24686\,
            lcout => \tok.A_stk.tail_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28544\,
            ce => \N__26078\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i47_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24694\,
            in1 => \N__26604\,
            in2 => \_gnd_net_\,
            in3 => \N__24650\,
            lcout => \tok.A_stk.tail_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28544\,
            ce => \N__26078\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i63_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26605\,
            in1 => \N__24685\,
            in2 => \_gnd_net_\,
            in3 => \N__24634\,
            lcout => \tok.A_stk.tail_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28544\,
            ce => \N__26078\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i79_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24677\,
            in1 => \N__26606\,
            in2 => \_gnd_net_\,
            in3 => \N__24649\,
            lcout => \tok.A_stk.tail_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28544\,
            ce => \N__26078\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i90_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25207\,
            in1 => \N__24982\,
            in2 => \_gnd_net_\,
            in3 => \N__26573\,
            lcout => \tok.A_stk.tail_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28521\,
            ce => \N__26071\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i42_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26570\,
            in1 => \_gnd_net_\,
            in2 => \N__24974\,
            in3 => \N__24952\,
            lcout => \tok.A_stk.tail_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28521\,
            ce => \N__26071\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i74_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25247\,
            in1 => \N__24970\,
            in2 => \_gnd_net_\,
            in3 => \N__26572\,
            lcout => \tok.A_stk.tail_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28521\,
            ce => \N__26071\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i58_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26571\,
            in1 => \_gnd_net_\,
            in2 => \N__24986\,
            in3 => \N__24961\,
            lcout => \tok.A_stk.tail_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28521\,
            ce => \N__26071\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i26_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__26569\,
            in1 => \_gnd_net_\,
            in2 => \N__24944\,
            in3 => \N__24962\,
            lcout => \tok.A_stk.tail_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28521\,
            ce => \N__26071\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i10_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24953\,
            in1 => \N__26568\,
            in2 => \_gnd_net_\,
            in3 => \N__27414\,
            lcout => \tok.A_stk.tail_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28521\,
            ce => \N__26071\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i10_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24940\,
            in1 => \N__25511\,
            in2 => \_gnd_net_\,
            in3 => \N__29282\,
            lcout => \tok.S_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28521\,
            ce => \N__26071\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i101_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24932\,
            in1 => \N__24892\,
            in2 => \_gnd_net_\,
            in3 => \N__26518\,
            lcout => tail_101,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28526\,
            ce => \N__25986\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i85_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26525\,
            in1 => \N__24904\,
            in2 => \_gnd_net_\,
            in3 => \N__24880\,
            lcout => \tok.A_stk.tail_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28526\,
            ce => \N__25986\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i69_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24893\,
            in1 => \N__25273\,
            in2 => \_gnd_net_\,
            in3 => \N__26524\,
            lcout => \tok.A_stk.tail_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28526\,
            ce => \N__25986\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i53_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26522\,
            in1 => \N__25264\,
            in2 => \_gnd_net_\,
            in3 => \N__24881\,
            lcout => \tok.A_stk.tail_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28526\,
            ce => \N__25986\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i37_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25255\,
            in1 => \N__25274\,
            in2 => \_gnd_net_\,
            in3 => \N__26521\,
            lcout => \tok.A_stk.tail_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28526\,
            ce => \N__25986\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i21_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26520\,
            in1 => \N__25265\,
            in2 => \_gnd_net_\,
            in3 => \N__25390\,
            lcout => \tok.A_stk.tail_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28526\,
            ce => \N__25986\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i5_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25256\,
            in1 => \N__26523\,
            in2 => \_gnd_net_\,
            in3 => \N__27187\,
            lcout => \tok.A_stk.tail_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28526\,
            ce => \N__25986\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i106_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26519\,
            in1 => \N__25246\,
            in2 => \_gnd_net_\,
            in3 => \N__25235\,
            lcout => tail_106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28526\,
            ce => \N__25986\,
            sr => \_gnd_net_\
        );

    \tok.i7_4_lut_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__25762\,
            in1 => \N__25009\,
            in2 => \N__28837\,
            in3 => \N__25168\,
            lcout => \tok.n23_adj_642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i15_1_lut_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25761\,
            lcout => \tok.n288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i11_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25594\,
            in1 => \N__25502\,
            in2 => \_gnd_net_\,
            in3 => \N__25169\,
            lcout => \tok.S_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28529\,
            ce => \N__26060\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i14_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25503\,
            in1 => \N__25082\,
            in2 => \_gnd_net_\,
            in3 => \N__25763\,
            lcout => \tok.S_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28529\,
            ce => \N__26060\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i11_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25586\,
            in1 => \N__26583\,
            in2 => \_gnd_net_\,
            in3 => \N__25010\,
            lcout => \tok.A_stk.tail_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28529\,
            ce => \N__26060\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i27_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26584\,
            in1 => \N__25595\,
            in2 => \_gnd_net_\,
            in3 => \N__25577\,
            lcout => \tok.A_stk.tail_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28529\,
            ce => \N__26060\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i43_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25585\,
            in1 => \N__25549\,
            in2 => \_gnd_net_\,
            in3 => \N__26585\,
            lcout => \tok.A_stk.tail_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28529\,
            ce => \N__26060\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i59_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26586\,
            in1 => \N__25576\,
            in2 => \_gnd_net_\,
            in3 => \N__25568\,
            lcout => \tok.A_stk.tail_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28529\,
            ce => \N__26060\,
            sr => \_gnd_net_\
        );

    \tok.i4_4_lut_adj_31_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__29733\,
            in1 => \N__25328\,
            in2 => \N__27196\,
            in3 => \N__27290\,
            lcout => \tok.n20_adj_648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i4_1_lut_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29732\,
            lcout => \tok.n299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29734\,
            in1 => \N__25282\,
            in2 => \_gnd_net_\,
            in3 => \N__25504\,
            lcout => \tok.S_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28534\,
            ce => \N__26074\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.head_i0_i5_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27291\,
            in1 => \_gnd_net_\,
            in2 => \N__25513\,
            in3 => \N__25394\,
            lcout => \tok.S_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28534\,
            ce => \N__26074\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i3_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26589\,
            in1 => \N__26645\,
            in2 => \_gnd_net_\,
            in3 => \N__25329\,
            lcout => \tok.A_stk.tail_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28534\,
            ce => \N__26074\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i19_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26636\,
            in1 => \_gnd_net_\,
            in2 => \N__25286\,
            in3 => \N__26587\,
            lcout => \tok.A_stk.tail_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28534\,
            ce => \N__26074\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i35_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__26588\,
            in1 => \N__26644\,
            in2 => \_gnd_net_\,
            in3 => \N__26092\,
            lcout => \tok.A_stk.tail_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28534\,
            ce => \N__26074\,
            sr => \_gnd_net_\
        );

    \tok.A_stk.tail_i0_i51_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26635\,
            in1 => \N__26627\,
            in2 => \_gnd_net_\,
            in3 => \N__26590\,
            lcout => \tok.A_stk.tail_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28534\,
            ce => \N__26074\,
            sr => \_gnd_net_\
        );

    \tok.i5240_3_lut_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__27886\,
            in1 => \N__26795\,
            in2 => \_gnd_net_\,
            in3 => \N__25742\,
            lcout => \tok.n5412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_112_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__27654\,
            in1 => \N__25817\,
            in2 => \N__25764\,
            in3 => \N__26764\,
            lcout => OPEN,
            ltout => \tok.n13_adj_772_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_113_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__25811\,
            in1 => \N__25799\,
            in2 => \N__25784\,
            in3 => \N__25781\,
            lcout => OPEN,
            ltout => \tok.n22_adj_773_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i15_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__28626\,
            in1 => \N__28850\,
            in2 => \N__25775\,
            in3 => \N__28667\,
            lcout => \tok.A_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28540\,
            ce => \N__28301\,
            sr => \N__28233\
        );

    \tok.A_i6_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110001011100"
        )
    port map (
            in0 => \N__26796\,
            in1 => \N__27180\,
            in2 => \N__28638\,
            in3 => \N__27002\,
            lcout => \tok.A_low_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28540\,
            ce => \N__28301\,
            sr => \N__28233\
        );

    \tok.i2_3_lut_adj_189_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__27885\,
            in1 => \N__27292\,
            in2 => \_gnd_net_\,
            in3 => \N__27653\,
            lcout => \tok.n14_adj_856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.uart.rx_data_i0_i5_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25693\,
            in1 => \N__25616\,
            in2 => \_gnd_net_\,
            in3 => \N__27124\,
            lcout => uart_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_adj_192_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__27195\,
            in1 => \N__27957\,
            in2 => \N__27125\,
            in3 => \N__28788\,
            lcout => \tok.n18_adj_860\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i8_4_lut_adj_190_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__27113\,
            in1 => \N__26995\,
            in2 => \N__27107\,
            in3 => \N__27077\,
            lcout => OPEN,
            ltout => \tok.n20_adj_857_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_adj_193_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27071\,
            in1 => \N__27056\,
            in2 => \N__27044\,
            in3 => \N__27041\,
            lcout => OPEN,
            ltout => \tok.n22_adj_861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5564_4_lut_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27035\,
            in1 => \N__27026\,
            in2 => \N__27011\,
            in3 => \N__27008\,
            lcout => \tok.n5556\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i3_3_lut_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__26996\,
            in1 => \N__26891\,
            in2 => \_gnd_net_\,
            in3 => \N__26882\,
            lcout => \tok.n15_adj_670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5244_3_lut_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__27884\,
            in1 => \_gnd_net_\,
            in2 => \N__26829\,
            in3 => \N__29411\,
            lcout => \tok.n5416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_43_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__27656\,
            in1 => \N__26780\,
            in2 => \N__29441\,
            in3 => \N__26753\,
            lcout => OPEN,
            ltout => \tok.n13_adj_674_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i10_4_lut_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__26660\,
            in1 => \N__27893\,
            in2 => \N__26654\,
            in3 => \N__26651\,
            lcout => OPEN,
            ltout => \tok.n22_adj_676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.A_i9_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__28648\,
            in1 => \N__28072\,
            in2 => \N__28547\,
            in3 => \N__27977\,
            lcout => \tok.A_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__28543\,
            ce => \N__28292\,
            sr => \N__28231\
        );

    \tok.i5496_4_lut_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__28071\,
            in1 => \N__28784\,
            in2 => \N__27986\,
            in3 => \N__29477\,
            lcout => \tok.n5542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i2_3_lut_adj_41_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__27785\,
            in1 => \N__27971\,
            in2 => \_gnd_net_\,
            in3 => \N__27958\,
            lcout => \tok.n14_adj_668\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i45_3_lut_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27883\,
            in1 => \N__27784\,
            in2 => \_gnd_net_\,
            in3 => \N__27655\,
            lcout => \tok.n5372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_52_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__28935\,
            in1 => \N__28785\,
            in2 => \N__27554\,
            in3 => \N__29565\,
            lcout => \tok.n8_adj_689\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i1_4_lut_adj_61_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110011"
        )
    port map (
            in0 => \N__28786\,
            in1 => \N__27297\,
            in2 => \N__27448\,
            in3 => \N__28937\,
            lcout => \tok.n8_adj_702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i5_1_lut_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29564\,
            lcout => \tok.n298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i6_1_lut_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27296\,
            lcout => \tok.n297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5197_2_lut_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__28936\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30032\,
            lcout => \tok.n5366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5225_2_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29703\,
            in2 => \_gnd_net_\,
            in3 => \N__28938\,
            lcout => OPEN,
            ltout => \tok.n5396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_4_lut_adj_183_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111101111"
        )
    port map (
            in0 => \N__29353\,
            in1 => \N__29566\,
            in2 => \N__29480\,
            in3 => \N__29179\,
            lcout => \tok.n18_adj_677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.inv_106_i9_1_lut_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29407\,
            lcout => \tok.n294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.or_101_i15_2_lut_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29354\,
            in2 => \_gnd_net_\,
            in3 => \N__29278\,
            lcout => OPEN,
            ltout => \tok.n202_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i6_4_lut_4_lut_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__29180\,
            in1 => \N__29066\,
            in2 => \N__28982\,
            in3 => \N__28977\,
            lcout => OPEN,
            ltout => \tok.n18_adj_774_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tok.i5455_4_lut_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__28874\,
            in1 => \N__28858\,
            in2 => \N__28793\,
            in3 => \N__28787\,
            lcout => \tok.n5518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
