// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Dec 31 2020 10:49:39

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    tx,
    rx,
    reset);

    output tx;
    input rx;
    input reset;

    wire N__30609;
    wire N__30608;
    wire N__30607;
    wire N__30600;
    wire N__30599;
    wire N__30598;
    wire N__30591;
    wire N__30590;
    wire N__30589;
    wire N__30572;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30545;
    wire N__30542;
    wire N__30539;
    wire N__30538;
    wire N__30537;
    wire N__30536;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30505;
    wire N__30500;
    wire N__30497;
    wire N__30494;
    wire N__30493;
    wire N__30490;
    wire N__30489;
    wire N__30488;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30452;
    wire N__30449;
    wire N__30448;
    wire N__30447;
    wire N__30446;
    wire N__30445;
    wire N__30444;
    wire N__30443;
    wire N__30442;
    wire N__30441;
    wire N__30438;
    wire N__30433;
    wire N__30424;
    wire N__30423;
    wire N__30420;
    wire N__30419;
    wire N__30418;
    wire N__30417;
    wire N__30416;
    wire N__30413;
    wire N__30412;
    wire N__30411;
    wire N__30410;
    wire N__30405;
    wire N__30402;
    wire N__30395;
    wire N__30394;
    wire N__30393;
    wire N__30392;
    wire N__30391;
    wire N__30390;
    wire N__30389;
    wire N__30386;
    wire N__30385;
    wire N__30384;
    wire N__30383;
    wire N__30382;
    wire N__30381;
    wire N__30380;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30363;
    wire N__30356;
    wire N__30353;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30345;
    wire N__30340;
    wire N__30333;
    wire N__30324;
    wire N__30323;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30291;
    wire N__30290;
    wire N__30289;
    wire N__30288;
    wire N__30287;
    wire N__30286;
    wire N__30283;
    wire N__30282;
    wire N__30281;
    wire N__30280;
    wire N__30279;
    wire N__30276;
    wire N__30271;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30253;
    wire N__30250;
    wire N__30245;
    wire N__30238;
    wire N__30231;
    wire N__30220;
    wire N__30213;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30164;
    wire N__30163;
    wire N__30162;
    wire N__30161;
    wire N__30160;
    wire N__30159;
    wire N__30158;
    wire N__30157;
    wire N__30156;
    wire N__30155;
    wire N__30154;
    wire N__30153;
    wire N__30152;
    wire N__30151;
    wire N__30150;
    wire N__30149;
    wire N__30148;
    wire N__30147;
    wire N__30146;
    wire N__30145;
    wire N__30138;
    wire N__30137;
    wire N__30136;
    wire N__30135;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30121;
    wire N__30114;
    wire N__30113;
    wire N__30112;
    wire N__30111;
    wire N__30110;
    wire N__30109;
    wire N__30108;
    wire N__30107;
    wire N__30106;
    wire N__30105;
    wire N__30104;
    wire N__30103;
    wire N__30102;
    wire N__30099;
    wire N__30094;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30045;
    wire N__30044;
    wire N__30041;
    wire N__30040;
    wire N__30037;
    wire N__30030;
    wire N__30021;
    wire N__30020;
    wire N__30015;
    wire N__30010;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29975;
    wire N__29974;
    wire N__29973;
    wire N__29970;
    wire N__29969;
    wire N__29968;
    wire N__29967;
    wire N__29966;
    wire N__29965;
    wire N__29964;
    wire N__29963;
    wire N__29962;
    wire N__29959;
    wire N__29954;
    wire N__29951;
    wire N__29944;
    wire N__29931;
    wire N__29928;
    wire N__29921;
    wire N__29914;
    wire N__29911;
    wire N__29900;
    wire N__29893;
    wire N__29876;
    wire N__29873;
    wire N__29872;
    wire N__29871;
    wire N__29870;
    wire N__29869;
    wire N__29868;
    wire N__29867;
    wire N__29866;
    wire N__29865;
    wire N__29864;
    wire N__29863;
    wire N__29862;
    wire N__29861;
    wire N__29860;
    wire N__29859;
    wire N__29858;
    wire N__29857;
    wire N__29856;
    wire N__29855;
    wire N__29854;
    wire N__29853;
    wire N__29852;
    wire N__29851;
    wire N__29850;
    wire N__29849;
    wire N__29848;
    wire N__29847;
    wire N__29844;
    wire N__29837;
    wire N__29832;
    wire N__29825;
    wire N__29824;
    wire N__29821;
    wire N__29820;
    wire N__29819;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29803;
    wire N__29802;
    wire N__29801;
    wire N__29800;
    wire N__29799;
    wire N__29794;
    wire N__29791;
    wire N__29786;
    wire N__29783;
    wire N__29782;
    wire N__29779;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29757;
    wire N__29754;
    wire N__29747;
    wire N__29738;
    wire N__29733;
    wire N__29728;
    wire N__29725;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29697;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29685;
    wire N__29684;
    wire N__29683;
    wire N__29682;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29678;
    wire N__29677;
    wire N__29676;
    wire N__29675;
    wire N__29674;
    wire N__29671;
    wire N__29666;
    wire N__29663;
    wire N__29648;
    wire N__29643;
    wire N__29636;
    wire N__29621;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29575;
    wire N__29574;
    wire N__29573;
    wire N__29572;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29549;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29519;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29487;
    wire N__29480;
    wire N__29473;
    wire N__29470;
    wire N__29465;
    wire N__29462;
    wire N__29461;
    wire N__29460;
    wire N__29459;
    wire N__29458;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29446;
    wire N__29445;
    wire N__29444;
    wire N__29441;
    wire N__29440;
    wire N__29437;
    wire N__29436;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29398;
    wire N__29395;
    wire N__29394;
    wire N__29393;
    wire N__29392;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29371;
    wire N__29368;
    wire N__29363;
    wire N__29358;
    wire N__29353;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29326;
    wire N__29323;
    wire N__29322;
    wire N__29321;
    wire N__29318;
    wire N__29317;
    wire N__29306;
    wire N__29305;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29294;
    wire N__29293;
    wire N__29292;
    wire N__29291;
    wire N__29286;
    wire N__29285;
    wire N__29284;
    wire N__29283;
    wire N__29282;
    wire N__29281;
    wire N__29280;
    wire N__29279;
    wire N__29278;
    wire N__29275;
    wire N__29268;
    wire N__29267;
    wire N__29266;
    wire N__29265;
    wire N__29262;
    wire N__29261;
    wire N__29260;
    wire N__29259;
    wire N__29258;
    wire N__29255;
    wire N__29252;
    wire N__29251;
    wire N__29248;
    wire N__29247;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29226;
    wire N__29223;
    wire N__29222;
    wire N__29221;
    wire N__29218;
    wire N__29209;
    wire N__29204;
    wire N__29199;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29181;
    wire N__29170;
    wire N__29165;
    wire N__29162;
    wire N__29155;
    wire N__29150;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29138;
    wire N__29135;
    wire N__29126;
    wire N__29123;
    wire N__29122;
    wire N__29121;
    wire N__29118;
    wire N__29113;
    wire N__29108;
    wire N__29107;
    wire N__29106;
    wire N__29105;
    wire N__29104;
    wire N__29103;
    wire N__29102;
    wire N__29101;
    wire N__29096;
    wire N__29085;
    wire N__29082;
    wire N__29081;
    wire N__29080;
    wire N__29079;
    wire N__29078;
    wire N__29077;
    wire N__29072;
    wire N__29069;
    wire N__29064;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29046;
    wire N__29043;
    wire N__29036;
    wire N__29035;
    wire N__29034;
    wire N__29033;
    wire N__29032;
    wire N__29031;
    wire N__29030;
    wire N__29029;
    wire N__29028;
    wire N__29027;
    wire N__29026;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29010;
    wire N__29009;
    wire N__29008;
    wire N__29007;
    wire N__29000;
    wire N__28999;
    wire N__28998;
    wire N__28991;
    wire N__28990;
    wire N__28989;
    wire N__28986;
    wire N__28981;
    wire N__28974;
    wire N__28973;
    wire N__28972;
    wire N__28971;
    wire N__28968;
    wire N__28963;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28945;
    wire N__28942;
    wire N__28941;
    wire N__28940;
    wire N__28939;
    wire N__28936;
    wire N__28935;
    wire N__28934;
    wire N__28931;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28907;
    wire N__28906;
    wire N__28905;
    wire N__28904;
    wire N__28903;
    wire N__28900;
    wire N__28895;
    wire N__28892;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28876;
    wire N__28869;
    wire N__28866;
    wire N__28859;
    wire N__28850;
    wire N__28835;
    wire N__28834;
    wire N__28833;
    wire N__28832;
    wire N__28831;
    wire N__28830;
    wire N__28829;
    wire N__28828;
    wire N__28823;
    wire N__28822;
    wire N__28821;
    wire N__28816;
    wire N__28813;
    wire N__28812;
    wire N__28809;
    wire N__28808;
    wire N__28807;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28793;
    wire N__28790;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28775;
    wire N__28774;
    wire N__28773;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28757;
    wire N__28752;
    wire N__28747;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28728;
    wire N__28723;
    wire N__28720;
    wire N__28713;
    wire N__28700;
    wire N__28699;
    wire N__28698;
    wire N__28697;
    wire N__28694;
    wire N__28693;
    wire N__28692;
    wire N__28691;
    wire N__28690;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28679;
    wire N__28678;
    wire N__28671;
    wire N__28668;
    wire N__28663;
    wire N__28662;
    wire N__28659;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28638;
    wire N__28635;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28627;
    wire N__28626;
    wire N__28625;
    wire N__28622;
    wire N__28617;
    wire N__28608;
    wire N__28605;
    wire N__28600;
    wire N__28595;
    wire N__28594;
    wire N__28591;
    wire N__28590;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28574;
    wire N__28567;
    wire N__28556;
    wire N__28555;
    wire N__28554;
    wire N__28551;
    wire N__28550;
    wire N__28549;
    wire N__28548;
    wire N__28545;
    wire N__28544;
    wire N__28543;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28532;
    wire N__28531;
    wire N__28530;
    wire N__28529;
    wire N__28528;
    wire N__28525;
    wire N__28524;
    wire N__28523;
    wire N__28518;
    wire N__28517;
    wire N__28514;
    wire N__28513;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28505;
    wire N__28504;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28481;
    wire N__28478;
    wire N__28473;
    wire N__28470;
    wire N__28465;
    wire N__28460;
    wire N__28459;
    wire N__28454;
    wire N__28451;
    wire N__28450;
    wire N__28449;
    wire N__28446;
    wire N__28439;
    wire N__28436;
    wire N__28431;
    wire N__28428;
    wire N__28417;
    wire N__28416;
    wire N__28413;
    wire N__28408;
    wire N__28403;
    wire N__28402;
    wire N__28401;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28383;
    wire N__28380;
    wire N__28373;
    wire N__28366;
    wire N__28349;
    wire N__28348;
    wire N__28345;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28337;
    wire N__28334;
    wire N__28329;
    wire N__28326;
    wire N__28325;
    wire N__28324;
    wire N__28323;
    wire N__28316;
    wire N__28313;
    wire N__28308;
    wire N__28303;
    wire N__28300;
    wire N__28299;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28270;
    wire N__28269;
    wire N__28268;
    wire N__28265;
    wire N__28264;
    wire N__28261;
    wire N__28260;
    wire N__28259;
    wire N__28256;
    wire N__28255;
    wire N__28254;
    wire N__28253;
    wire N__28252;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28219;
    wire N__28218;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28184;
    wire N__28179;
    wire N__28176;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28148;
    wire N__28145;
    wire N__28142;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28117;
    wire N__28116;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28104;
    wire N__28103;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28088;
    wire N__28079;
    wire N__28076;
    wire N__28075;
    wire N__28074;
    wire N__28073;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28058;
    wire N__28057;
    wire N__28056;
    wire N__28055;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28040;
    wire N__28037;
    wire N__28032;
    wire N__28019;
    wire N__28018;
    wire N__28017;
    wire N__28016;
    wire N__28015;
    wire N__28014;
    wire N__28013;
    wire N__28012;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__28001;
    wire N__28000;
    wire N__27999;
    wire N__27994;
    wire N__27993;
    wire N__27992;
    wire N__27989;
    wire N__27988;
    wire N__27987;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27979;
    wire N__27976;
    wire N__27969;
    wire N__27966;
    wire N__27963;
    wire N__27960;
    wire N__27957;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27939;
    wire N__27936;
    wire N__27931;
    wire N__27930;
    wire N__27929;
    wire N__27928;
    wire N__27927;
    wire N__27926;
    wire N__27925;
    wire N__27924;
    wire N__27923;
    wire N__27920;
    wire N__27915;
    wire N__27908;
    wire N__27905;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27884;
    wire N__27881;
    wire N__27880;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27869;
    wire N__27868;
    wire N__27865;
    wire N__27860;
    wire N__27857;
    wire N__27848;
    wire N__27841;
    wire N__27834;
    wire N__27819;
    wire N__27806;
    wire N__27805;
    wire N__27804;
    wire N__27801;
    wire N__27796;
    wire N__27795;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27781;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27763;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27749;
    wire N__27746;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27691;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27676;
    wire N__27671;
    wire N__27668;
    wire N__27667;
    wire N__27666;
    wire N__27665;
    wire N__27664;
    wire N__27663;
    wire N__27662;
    wire N__27661;
    wire N__27660;
    wire N__27659;
    wire N__27658;
    wire N__27657;
    wire N__27656;
    wire N__27655;
    wire N__27654;
    wire N__27653;
    wire N__27646;
    wire N__27637;
    wire N__27626;
    wire N__27617;
    wire N__27614;
    wire N__27607;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27571;
    wire N__27570;
    wire N__27567;
    wire N__27562;
    wire N__27557;
    wire N__27556;
    wire N__27555;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27539;
    wire N__27538;
    wire N__27533;
    wire N__27530;
    wire N__27529;
    wire N__27528;
    wire N__27525;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27448;
    wire N__27447;
    wire N__27446;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27435;
    wire N__27434;
    wire N__27433;
    wire N__27430;
    wire N__27429;
    wire N__27428;
    wire N__27427;
    wire N__27424;
    wire N__27423;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27411;
    wire N__27408;
    wire N__27403;
    wire N__27400;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27378;
    wire N__27375;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27346;
    wire N__27341;
    wire N__27334;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27268;
    wire N__27267;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27245;
    wire N__27244;
    wire N__27243;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27232;
    wire N__27229;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27218;
    wire N__27217;
    wire N__27216;
    wire N__27215;
    wire N__27212;
    wire N__27211;
    wire N__27210;
    wire N__27209;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27192;
    wire N__27189;
    wire N__27188;
    wire N__27181;
    wire N__27178;
    wire N__27169;
    wire N__27168;
    wire N__27163;
    wire N__27160;
    wire N__27155;
    wire N__27148;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27073;
    wire N__27072;
    wire N__27071;
    wire N__27068;
    wire N__27067;
    wire N__27064;
    wire N__27063;
    wire N__27062;
    wire N__27061;
    wire N__27058;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27050;
    wire N__27047;
    wire N__27046;
    wire N__27045;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27001;
    wire N__26998;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26963;
    wire N__26958;
    wire N__26955;
    wire N__26942;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26934;
    wire N__26933;
    wire N__26930;
    wire N__26929;
    wire N__26928;
    wire N__26927;
    wire N__26926;
    wire N__26925;
    wire N__26922;
    wire N__26921;
    wire N__26920;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26900;
    wire N__26899;
    wire N__26894;
    wire N__26891;
    wire N__26886;
    wire N__26883;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26871;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26850;
    wire N__26847;
    wire N__26840;
    wire N__26835;
    wire N__26832;
    wire N__26819;
    wire N__26816;
    wire N__26815;
    wire N__26814;
    wire N__26813;
    wire N__26812;
    wire N__26811;
    wire N__26810;
    wire N__26805;
    wire N__26804;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26796;
    wire N__26795;
    wire N__26792;
    wire N__26791;
    wire N__26790;
    wire N__26789;
    wire N__26784;
    wire N__26781;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26754;
    wire N__26749;
    wire N__26742;
    wire N__26739;
    wire N__26734;
    wire N__26731;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26717;
    wire N__26714;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26696;
    wire N__26695;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26684;
    wire N__26683;
    wire N__26682;
    wire N__26679;
    wire N__26674;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26659;
    wire N__26656;
    wire N__26651;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26639;
    wire N__26636;
    wire N__26627;
    wire N__26624;
    wire N__26623;
    wire N__26622;
    wire N__26619;
    wire N__26618;
    wire N__26617;
    wire N__26616;
    wire N__26615;
    wire N__26610;
    wire N__26605;
    wire N__26604;
    wire N__26603;
    wire N__26602;
    wire N__26601;
    wire N__26600;
    wire N__26599;
    wire N__26598;
    wire N__26597;
    wire N__26592;
    wire N__26589;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26563;
    wire N__26562;
    wire N__26559;
    wire N__26554;
    wire N__26549;
    wire N__26544;
    wire N__26539;
    wire N__26536;
    wire N__26529;
    wire N__26526;
    wire N__26521;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26498;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26486;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26456;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26417;
    wire N__26416;
    wire N__26411;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26388;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26363;
    wire N__26360;
    wire N__26359;
    wire N__26358;
    wire N__26353;
    wire N__26352;
    wire N__26349;
    wire N__26348;
    wire N__26347;
    wire N__26346;
    wire N__26345;
    wire N__26342;
    wire N__26337;
    wire N__26332;
    wire N__26331;
    wire N__26330;
    wire N__26325;
    wire N__26324;
    wire N__26323;
    wire N__26322;
    wire N__26317;
    wire N__26314;
    wire N__26309;
    wire N__26306;
    wire N__26305;
    wire N__26304;
    wire N__26303;
    wire N__26296;
    wire N__26291;
    wire N__26286;
    wire N__26279;
    wire N__26270;
    wire N__26269;
    wire N__26268;
    wire N__26267;
    wire N__26266;
    wire N__26265;
    wire N__26264;
    wire N__26263;
    wire N__26262;
    wire N__26261;
    wire N__26260;
    wire N__26259;
    wire N__26258;
    wire N__26257;
    wire N__26256;
    wire N__26255;
    wire N__26254;
    wire N__26253;
    wire N__26252;
    wire N__26251;
    wire N__26250;
    wire N__26249;
    wire N__26248;
    wire N__26247;
    wire N__26246;
    wire N__26245;
    wire N__26244;
    wire N__26243;
    wire N__26242;
    wire N__26241;
    wire N__26240;
    wire N__26239;
    wire N__26238;
    wire N__26237;
    wire N__26236;
    wire N__26235;
    wire N__26234;
    wire N__26233;
    wire N__26232;
    wire N__26231;
    wire N__26230;
    wire N__26229;
    wire N__26228;
    wire N__26227;
    wire N__26226;
    wire N__26225;
    wire N__26224;
    wire N__26223;
    wire N__26222;
    wire N__26221;
    wire N__26220;
    wire N__26219;
    wire N__26218;
    wire N__26217;
    wire N__26216;
    wire N__26215;
    wire N__26214;
    wire N__26213;
    wire N__26212;
    wire N__26211;
    wire N__26210;
    wire N__26209;
    wire N__26208;
    wire N__26207;
    wire N__26206;
    wire N__26205;
    wire N__26204;
    wire N__26203;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26199;
    wire N__26198;
    wire N__26197;
    wire N__26196;
    wire N__26195;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26032;
    wire N__26031;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26019;
    wire N__26016;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26000;
    wire N__25997;
    wire N__25996;
    wire N__25995;
    wire N__25994;
    wire N__25991;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25983;
    wire N__25980;
    wire N__25979;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25954;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25938;
    wire N__25933;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25909;
    wire N__25908;
    wire N__25905;
    wire N__25900;
    wire N__25899;
    wire N__25898;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25884;
    wire N__25881;
    wire N__25874;
    wire N__25873;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25825;
    wire N__25822;
    wire N__25821;
    wire N__25820;
    wire N__25817;
    wire N__25816;
    wire N__25813;
    wire N__25806;
    wire N__25803;
    wire N__25796;
    wire N__25793;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25733;
    wire N__25732;
    wire N__25731;
    wire N__25730;
    wire N__25729;
    wire N__25728;
    wire N__25727;
    wire N__25726;
    wire N__25725;
    wire N__25724;
    wire N__25723;
    wire N__25722;
    wire N__25721;
    wire N__25720;
    wire N__25719;
    wire N__25718;
    wire N__25717;
    wire N__25716;
    wire N__25715;
    wire N__25714;
    wire N__25713;
    wire N__25712;
    wire N__25711;
    wire N__25710;
    wire N__25709;
    wire N__25708;
    wire N__25707;
    wire N__25706;
    wire N__25705;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25697;
    wire N__25696;
    wire N__25695;
    wire N__25678;
    wire N__25661;
    wire N__25660;
    wire N__25643;
    wire N__25642;
    wire N__25641;
    wire N__25640;
    wire N__25639;
    wire N__25638;
    wire N__25637;
    wire N__25636;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25622;
    wire N__25621;
    wire N__25620;
    wire N__25619;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25598;
    wire N__25597;
    wire N__25596;
    wire N__25595;
    wire N__25594;
    wire N__25593;
    wire N__25592;
    wire N__25591;
    wire N__25590;
    wire N__25589;
    wire N__25588;
    wire N__25587;
    wire N__25586;
    wire N__25585;
    wire N__25584;
    wire N__25583;
    wire N__25582;
    wire N__25581;
    wire N__25578;
    wire N__25561;
    wire N__25544;
    wire N__25537;
    wire N__25530;
    wire N__25513;
    wire N__25496;
    wire N__25493;
    wire N__25488;
    wire N__25485;
    wire N__25472;
    wire N__25471;
    wire N__25468;
    wire N__25467;
    wire N__25466;
    wire N__25465;
    wire N__25464;
    wire N__25463;
    wire N__25462;
    wire N__25461;
    wire N__25460;
    wire N__25459;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25428;
    wire N__25427;
    wire N__25426;
    wire N__25423;
    wire N__25422;
    wire N__25421;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25389;
    wire N__25386;
    wire N__25377;
    wire N__25364;
    wire N__25363;
    wire N__25360;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25352;
    wire N__25349;
    wire N__25344;
    wire N__25341;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25297;
    wire N__25296;
    wire N__25295;
    wire N__25292;
    wire N__25285;
    wire N__25280;
    wire N__25277;
    wire N__25276;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25265;
    wire N__25262;
    wire N__25261;
    wire N__25260;
    wire N__25259;
    wire N__25252;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25225;
    wire N__25222;
    wire N__25217;
    wire N__25208;
    wire N__25205;
    wire N__25204;
    wire N__25203;
    wire N__25202;
    wire N__25195;
    wire N__25192;
    wire N__25191;
    wire N__25190;
    wire N__25189;
    wire N__25184;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25160;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25133;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25111;
    wire N__25108;
    wire N__25107;
    wire N__25106;
    wire N__25105;
    wire N__25102;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25078;
    wire N__25075;
    wire N__25074;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25062;
    wire N__25059;
    wire N__25054;
    wire N__25043;
    wire N__25042;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25034;
    wire N__25031;
    wire N__25026;
    wire N__25023;
    wire N__25016;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25004;
    wire N__25003;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24974;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24941;
    wire N__24940;
    wire N__24935;
    wire N__24932;
    wire N__24931;
    wire N__24926;
    wire N__24923;
    wire N__24922;
    wire N__24917;
    wire N__24914;
    wire N__24913;
    wire N__24908;
    wire N__24905;
    wire N__24904;
    wire N__24899;
    wire N__24896;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24884;
    wire N__24883;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24868;
    wire N__24865;
    wire N__24862;
    wire N__24857;
    wire N__24856;
    wire N__24855;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24847;
    wire N__24846;
    wire N__24845;
    wire N__24844;
    wire N__24843;
    wire N__24840;
    wire N__24839;
    wire N__24836;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24798;
    wire N__24795;
    wire N__24794;
    wire N__24791;
    wire N__24786;
    wire N__24785;
    wire N__24782;
    wire N__24775;
    wire N__24770;
    wire N__24767;
    wire N__24762;
    wire N__24759;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24737;
    wire N__24736;
    wire N__24735;
    wire N__24730;
    wire N__24729;
    wire N__24728;
    wire N__24727;
    wire N__24726;
    wire N__24725;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24713;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24705;
    wire N__24704;
    wire N__24703;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24672;
    wire N__24667;
    wire N__24660;
    wire N__24659;
    wire N__24652;
    wire N__24645;
    wire N__24642;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24622;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24595;
    wire N__24590;
    wire N__24589;
    wire N__24586;
    wire N__24585;
    wire N__24584;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24567;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24553;
    wire N__24550;
    wire N__24547;
    wire N__24542;
    wire N__24541;
    wire N__24536;
    wire N__24533;
    wire N__24532;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24520;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24508;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24496;
    wire N__24495;
    wire N__24494;
    wire N__24493;
    wire N__24492;
    wire N__24491;
    wire N__24486;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24474;
    wire N__24473;
    wire N__24472;
    wire N__24471;
    wire N__24470;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24456;
    wire N__24451;
    wire N__24448;
    wire N__24443;
    wire N__24438;
    wire N__24435;
    wire N__24428;
    wire N__24425;
    wire N__24420;
    wire N__24415;
    wire N__24408;
    wire N__24403;
    wire N__24400;
    wire N__24395;
    wire N__24394;
    wire N__24393;
    wire N__24390;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24376;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24368;
    wire N__24367;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24315;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24247;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24187;
    wire N__24186;
    wire N__24185;
    wire N__24182;
    wire N__24181;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24173;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24149;
    wire N__24146;
    wire N__24141;
    wire N__24140;
    wire N__24137;
    wire N__24132;
    wire N__24131;
    wire N__24130;
    wire N__24129;
    wire N__24122;
    wire N__24119;
    wire N__24118;
    wire N__24113;
    wire N__24110;
    wire N__24105;
    wire N__24102;
    wire N__24097;
    wire N__24094;
    wire N__24089;
    wire N__24074;
    wire N__24073;
    wire N__24070;
    wire N__24069;
    wire N__24068;
    wire N__24067;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24031;
    wire N__24022;
    wire N__24019;
    wire N__24014;
    wire N__24013;
    wire N__24010;
    wire N__24009;
    wire N__24008;
    wire N__24005;
    wire N__24004;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23984;
    wire N__23983;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23952;
    wire N__23947;
    wire N__23942;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23899;
    wire N__23898;
    wire N__23897;
    wire N__23896;
    wire N__23895;
    wire N__23894;
    wire N__23893;
    wire N__23890;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23876;
    wire N__23875;
    wire N__23872;
    wire N__23871;
    wire N__23870;
    wire N__23869;
    wire N__23868;
    wire N__23867;
    wire N__23866;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23847;
    wire N__23838;
    wire N__23833;
    wire N__23828;
    wire N__23825;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23802;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23773;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23746;
    wire N__23745;
    wire N__23744;
    wire N__23741;
    wire N__23736;
    wire N__23733;
    wire N__23728;
    wire N__23725;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23692;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23620;
    wire N__23619;
    wire N__23616;
    wire N__23615;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23563;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23521;
    wire N__23520;
    wire N__23519;
    wire N__23518;
    wire N__23517;
    wire N__23516;
    wire N__23507;
    wire N__23506;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23499;
    wire N__23498;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23373;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23361;
    wire N__23356;
    wire N__23353;
    wire N__23348;
    wire N__23345;
    wire N__23344;
    wire N__23341;
    wire N__23338;
    wire N__23335;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23312;
    wire N__23311;
    wire N__23308;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23278;
    wire N__23275;
    wire N__23270;
    wire N__23267;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23255;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23243;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23231;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23210;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23198;
    wire N__23197;
    wire N__23192;
    wire N__23189;
    wire N__23188;
    wire N__23183;
    wire N__23180;
    wire N__23179;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23156;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23141;
    wire N__23138;
    wire N__23137;
    wire N__23132;
    wire N__23129;
    wire N__23128;
    wire N__23123;
    wire N__23120;
    wire N__23119;
    wire N__23114;
    wire N__23111;
    wire N__23110;
    wire N__23107;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23099;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23081;
    wire N__23078;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23056;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23005;
    wire N__23004;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22996;
    wire N__22995;
    wire N__22994;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22980;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22969;
    wire N__22966;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22932;
    wire N__22925;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22856;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22820;
    wire N__22819;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22720;
    wire N__22719;
    wire N__22718;
    wire N__22717;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22705;
    wire N__22702;
    wire N__22701;
    wire N__22698;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22680;
    wire N__22677;
    wire N__22672;
    wire N__22665;
    wire N__22658;
    wire N__22657;
    wire N__22656;
    wire N__22655;
    wire N__22652;
    wire N__22651;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22640;
    wire N__22637;
    wire N__22636;
    wire N__22633;
    wire N__22632;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22593;
    wire N__22590;
    wire N__22589;
    wire N__22588;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22566;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22550;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22528;
    wire N__22527;
    wire N__22526;
    wire N__22523;
    wire N__22522;
    wire N__22521;
    wire N__22520;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22508;
    wire N__22507;
    wire N__22504;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22493;
    wire N__22492;
    wire N__22491;
    wire N__22490;
    wire N__22489;
    wire N__22486;
    wire N__22481;
    wire N__22474;
    wire N__22469;
    wire N__22466;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22451;
    wire N__22450;
    wire N__22443;
    wire N__22440;
    wire N__22435;
    wire N__22430;
    wire N__22427;
    wire N__22422;
    wire N__22417;
    wire N__22414;
    wire N__22403;
    wire N__22402;
    wire N__22401;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22393;
    wire N__22390;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22376;
    wire N__22375;
    wire N__22374;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22366;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22350;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22338;
    wire N__22335;
    wire N__22334;
    wire N__22333;
    wire N__22332;
    wire N__22329;
    wire N__22322;
    wire N__22317;
    wire N__22312;
    wire N__22309;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22283;
    wire N__22282;
    wire N__22281;
    wire N__22278;
    wire N__22277;
    wire N__22274;
    wire N__22273;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22262;
    wire N__22261;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22240;
    wire N__22239;
    wire N__22238;
    wire N__22237;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22205;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22177;
    wire N__22176;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22138;
    wire N__22137;
    wire N__22134;
    wire N__22129;
    wire N__22124;
    wire N__22123;
    wire N__22122;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22114;
    wire N__22113;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22102;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22053;
    wire N__22046;
    wire N__22043;
    wire N__22038;
    wire N__22035;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21985;
    wire N__21982;
    wire N__21981;
    wire N__21978;
    wire N__21977;
    wire N__21976;
    wire N__21973;
    wire N__21972;
    wire N__21971;
    wire N__21968;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21957;
    wire N__21954;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21942;
    wire N__21939;
    wire N__21938;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21924;
    wire N__21921;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21893;
    wire N__21890;
    wire N__21885;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21850;
    wire N__21847;
    wire N__21846;
    wire N__21845;
    wire N__21842;
    wire N__21841;
    wire N__21840;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21832;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21824;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21813;
    wire N__21808;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21796;
    wire N__21795;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21743;
    wire N__21736;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21700;
    wire N__21699;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21691;
    wire N__21690;
    wire N__21689;
    wire N__21686;
    wire N__21685;
    wire N__21682;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21625;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21572;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21550;
    wire N__21547;
    wire N__21546;
    wire N__21545;
    wire N__21544;
    wire N__21541;
    wire N__21540;
    wire N__21539;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21492;
    wire N__21491;
    wire N__21484;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21436;
    wire N__21435;
    wire N__21434;
    wire N__21431;
    wire N__21430;
    wire N__21429;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21411;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21403;
    wire N__21402;
    wire N__21401;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21375;
    wire N__21370;
    wire N__21363;
    wire N__21358;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21326;
    wire N__21323;
    wire N__21322;
    wire N__21321;
    wire N__21320;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21303;
    wire N__21300;
    wire N__21299;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21270;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21258;
    wire N__21253;
    wire N__21250;
    wire N__21245;
    wire N__21240;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21207;
    wire N__21202;
    wire N__21199;
    wire N__21194;
    wire N__21193;
    wire N__21190;
    wire N__21185;
    wire N__21182;
    wire N__21181;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21173;
    wire N__21170;
    wire N__21169;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21096;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21055;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21034;
    wire N__21033;
    wire N__21032;
    wire N__21031;
    wire N__21030;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21001;
    wire N__20994;
    wire N__20987;
    wire N__20982;
    wire N__20977;
    wire N__20966;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20958;
    wire N__20955;
    wire N__20954;
    wire N__20953;
    wire N__20952;
    wire N__20949;
    wire N__20948;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20926;
    wire N__20923;
    wire N__20918;
    wire N__20913;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20869;
    wire N__20868;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20857;
    wire N__20854;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20843;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20792;
    wire N__20789;
    wire N__20784;
    wire N__20781;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20761;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20753;
    wire N__20752;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20732;
    wire N__20729;
    wire N__20724;
    wire N__20723;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20696;
    wire N__20693;
    wire N__20684;
    wire N__20681;
    wire N__20680;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20653;
    wire N__20652;
    wire N__20647;
    wire N__20644;
    wire N__20643;
    wire N__20642;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20627;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20611;
    wire N__20608;
    wire N__20597;
    wire N__20596;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20588;
    wire N__20587;
    wire N__20584;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20564;
    wire N__20563;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20513;
    wire N__20510;
    wire N__20509;
    wire N__20508;
    wire N__20507;
    wire N__20506;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20457;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20401;
    wire N__20400;
    wire N__20399;
    wire N__20396;
    wire N__20395;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20369;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20328;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20314;
    wire N__20313;
    wire N__20312;
    wire N__20311;
    wire N__20310;
    wire N__20309;
    wire N__20306;
    wire N__20305;
    wire N__20302;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20246;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20230;
    wire N__20225;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20170;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20155;
    wire N__20154;
    wire N__20151;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20113;
    wire N__20106;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20087;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20068;
    wire N__20065;
    wire N__20064;
    wire N__20061;
    wire N__20060;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20043;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20028;
    wire N__20025;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20006;
    wire N__20003;
    wire N__19998;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19977;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19951;
    wire N__19950;
    wire N__19949;
    wire N__19948;
    wire N__19947;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19906;
    wire N__19901;
    wire N__19898;
    wire N__19893;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19869;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19825;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19817;
    wire N__19814;
    wire N__19813;
    wire N__19812;
    wire N__19811;
    wire N__19808;
    wire N__19807;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19779;
    wire N__19776;
    wire N__19775;
    wire N__19774;
    wire N__19771;
    wire N__19766;
    wire N__19763;
    wire N__19762;
    wire N__19761;
    wire N__19758;
    wire N__19757;
    wire N__19754;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19732;
    wire N__19729;
    wire N__19722;
    wire N__19717;
    wire N__19714;
    wire N__19709;
    wire N__19704;
    wire N__19691;
    wire N__19690;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19679;
    wire N__19678;
    wire N__19675;
    wire N__19674;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19660;
    wire N__19657;
    wire N__19652;
    wire N__19649;
    wire N__19648;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19636;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19599;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19563;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19555;
    wire N__19554;
    wire N__19553;
    wire N__19550;
    wire N__19549;
    wire N__19546;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19492;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19469;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19433;
    wire N__19432;
    wire N__19431;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19409;
    wire N__19408;
    wire N__19407;
    wire N__19406;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19378;
    wire N__19377;
    wire N__19372;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19349;
    wire N__19346;
    wire N__19345;
    wire N__19344;
    wire N__19343;
    wire N__19340;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19313;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19299;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19283;
    wire N__19280;
    wire N__19279;
    wire N__19278;
    wire N__19277;
    wire N__19276;
    wire N__19275;
    wire N__19270;
    wire N__19261;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19232;
    wire N__19229;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19215;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19167;
    wire N__19164;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19144;
    wire N__19143;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19135;
    wire N__19132;
    wire N__19131;
    wire N__19130;
    wire N__19127;
    wire N__19122;
    wire N__19119;
    wire N__19118;
    wire N__19115;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19100;
    wire N__19097;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19086;
    wire N__19083;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19022;
    wire N__19017;
    wire N__19012;
    wire N__19007;
    wire N__19006;
    wire N__19005;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18991;
    wire N__18990;
    wire N__18989;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18973;
    wire N__18972;
    wire N__18971;
    wire N__18970;
    wire N__18969;
    wire N__18964;
    wire N__18955;
    wire N__18954;
    wire N__18949;
    wire N__18946;
    wire N__18941;
    wire N__18940;
    wire N__18937;
    wire N__18934;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18913;
    wire N__18912;
    wire N__18911;
    wire N__18908;
    wire N__18901;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18880;
    wire N__18879;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18867;
    wire N__18860;
    wire N__18857;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18845;
    wire N__18842;
    wire N__18841;
    wire N__18840;
    wire N__18837;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18815;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18803;
    wire N__18802;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18766;
    wire N__18765;
    wire N__18764;
    wire N__18761;
    wire N__18756;
    wire N__18753;
    wire N__18746;
    wire N__18745;
    wire N__18744;
    wire N__18743;
    wire N__18740;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18722;
    wire N__18719;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18673;
    wire N__18672;
    wire N__18671;
    wire N__18668;
    wire N__18661;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18643;
    wire N__18642;
    wire N__18641;
    wire N__18638;
    wire N__18631;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18604;
    wire N__18603;
    wire N__18602;
    wire N__18599;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18587;
    wire N__18584;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18524;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18512;
    wire N__18511;
    wire N__18508;
    wire N__18505;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18482;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18408;
    wire N__18407;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18340;
    wire N__18335;
    wire N__18334;
    wire N__18333;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18263;
    wire N__18262;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18213;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18175;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18160;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18136;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18097;
    wire N__18092;
    wire N__18089;
    wire N__18084;
    wire N__18081;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18067;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18055;
    wire N__18052;
    wire N__18049;
    wire N__18046;
    wire N__18045;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17923;
    wire N__17922;
    wire N__17921;
    wire N__17916;
    wire N__17913;
    wire N__17910;
    wire N__17909;
    wire N__17908;
    wire N__17905;
    wire N__17904;
    wire N__17899;
    wire N__17894;
    wire N__17893;
    wire N__17892;
    wire N__17891;
    wire N__17890;
    wire N__17889;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17881;
    wire N__17880;
    wire N__17875;
    wire N__17870;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17854;
    wire N__17849;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17818;
    wire N__17815;
    wire N__17812;
    wire N__17809;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17797;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17786;
    wire N__17785;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17749;
    wire N__17748;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17738;
    wire N__17737;
    wire N__17736;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17716;
    wire N__17715;
    wire N__17710;
    wire N__17703;
    wire N__17700;
    wire N__17693;
    wire N__17692;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17644;
    wire N__17643;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17631;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17617;
    wire N__17614;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17521;
    wire N__17520;
    wire N__17519;
    wire N__17518;
    wire N__17517;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17509;
    wire N__17508;
    wire N__17505;
    wire N__17502;
    wire N__17501;
    wire N__17500;
    wire N__17499;
    wire N__17498;
    wire N__17497;
    wire N__17490;
    wire N__17489;
    wire N__17488;
    wire N__17483;
    wire N__17480;
    wire N__17475;
    wire N__17472;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17442;
    wire N__17439;
    wire N__17436;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17416;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17389;
    wire N__17386;
    wire N__17385;
    wire N__17382;
    wire N__17381;
    wire N__17380;
    wire N__17379;
    wire N__17378;
    wire N__17375;
    wire N__17374;
    wire N__17371;
    wire N__17370;
    wire N__17369;
    wire N__17368;
    wire N__17361;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17349;
    wire N__17348;
    wire N__17347;
    wire N__17346;
    wire N__17345;
    wire N__17344;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17304;
    wire N__17297;
    wire N__17294;
    wire N__17289;
    wire N__17286;
    wire N__17279;
    wire N__17276;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17268;
    wire N__17267;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17228;
    wire N__17225;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17200;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17173;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17156;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17113;
    wire N__17112;
    wire N__17111;
    wire N__17110;
    wire N__17109;
    wire N__17108;
    wire N__17105;
    wire N__17100;
    wire N__17091;
    wire N__17090;
    wire N__17089;
    wire N__17088;
    wire N__17087;
    wire N__17086;
    wire N__17079;
    wire N__17074;
    wire N__17067;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17008;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16981;
    wire N__16976;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16964;
    wire N__16961;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16953;
    wire N__16948;
    wire N__16945;
    wire N__16944;
    wire N__16943;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16929;
    wire N__16928;
    wire N__16927;
    wire N__16926;
    wire N__16923;
    wire N__16922;
    wire N__16917;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16899;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16794;
    wire N__16789;
    wire N__16788;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16774;
    wire N__16771;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16708;
    wire N__16705;
    wire N__16702;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16685;
    wire N__16682;
    wire N__16681;
    wire N__16680;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16615;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16597;
    wire N__16594;
    wire N__16591;
    wire N__16588;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16559;
    wire N__16558;
    wire N__16553;
    wire N__16550;
    wire N__16549;
    wire N__16546;
    wire N__16543;
    wire N__16540;
    wire N__16537;
    wire N__16532;
    wire N__16531;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16471;
    wire N__16470;
    wire N__16469;
    wire N__16468;
    wire N__16467;
    wire N__16466;
    wire N__16465;
    wire N__16456;
    wire N__16449;
    wire N__16448;
    wire N__16447;
    wire N__16444;
    wire N__16439;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16427;
    wire N__16424;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16387;
    wire N__16386;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16367;
    wire N__16364;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16348;
    wire N__16345;
    wire N__16342;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16304;
    wire N__16301;
    wire N__16298;
    wire N__16295;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16265;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16199;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16051;
    wire N__16050;
    wire N__16049;
    wire N__16048;
    wire N__16047;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16039;
    wire N__16034;
    wire N__16025;
    wire N__16020;
    wire N__16015;
    wire N__16010;
    wire N__16009;
    wire N__16008;
    wire N__16003;
    wire N__16002;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15990;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15961;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15943;
    wire N__15942;
    wire N__15941;
    wire N__15940;
    wire N__15939;
    wire N__15936;
    wire N__15931;
    wire N__15928;
    wire N__15921;
    wire N__15914;
    wire N__15911;
    wire N__15910;
    wire N__15909;
    wire N__15902;
    wire N__15899;
    wire N__15898;
    wire N__15897;
    wire N__15896;
    wire N__15895;
    wire N__15894;
    wire N__15891;
    wire N__15890;
    wire N__15889;
    wire N__15886;
    wire N__15879;
    wire N__15870;
    wire N__15863;
    wire N__15860;
    wire N__15859;
    wire N__15858;
    wire N__15853;
    wire N__15850;
    wire N__15845;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15823;
    wire N__15820;
    wire N__15819;
    wire N__15818;
    wire N__15817;
    wire N__15814;
    wire N__15813;
    wire N__15808;
    wire N__15803;
    wire N__15798;
    wire N__15791;
    wire N__15788;
    wire N__15787;
    wire N__15786;
    wire N__15785;
    wire N__15784;
    wire N__15783;
    wire N__15778;
    wire N__15771;
    wire N__15768;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15745;
    wire N__15744;
    wire N__15743;
    wire N__15742;
    wire N__15741;
    wire N__15740;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15732;
    wire N__15731;
    wire N__15728;
    wire N__15725;
    wire N__15724;
    wire N__15721;
    wire N__15720;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15682;
    wire N__15681;
    wire N__15678;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15658;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15627;
    wire N__15624;
    wire N__15615;
    wire N__15602;
    wire N__15599;
    wire N__15598;
    wire N__15597;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15578;
    wire N__15577;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15553;
    wire N__15548;
    wire N__15545;
    wire N__15544;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15532;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15520;
    wire N__15515;
    wire N__15512;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15500;
    wire N__15499;
    wire N__15494;
    wire N__15491;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15479;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15322;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15125;
    wire N__15122;
    wire N__15121;
    wire N__15118;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15085;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15043;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14918;
    wire N__14915;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14903;
    wire N__14900;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14737;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14729;
    wire N__14728;
    wire N__14727;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14717;
    wire N__14714;
    wire N__14713;
    wire N__14712;
    wire N__14709;
    wire N__14708;
    wire N__14707;
    wire N__14704;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14682;
    wire N__14681;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14664;
    wire N__14661;
    wire N__14656;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14634;
    wire N__14631;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14606;
    wire N__14597;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14558;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14546;
    wire N__14543;
    wire N__14542;
    wire N__14541;
    wire N__14540;
    wire N__14539;
    wire N__14538;
    wire N__14537;
    wire N__14536;
    wire N__14535;
    wire N__14534;
    wire N__14533;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14529;
    wire N__14528;
    wire N__14527;
    wire N__14526;
    wire N__14525;
    wire N__14524;
    wire N__14523;
    wire N__14522;
    wire N__14521;
    wire N__14520;
    wire N__14519;
    wire N__14518;
    wire N__14517;
    wire N__14516;
    wire N__14515;
    wire N__14514;
    wire N__14513;
    wire N__14512;
    wire N__14511;
    wire N__14510;
    wire N__14509;
    wire N__14508;
    wire N__14507;
    wire N__14506;
    wire N__14491;
    wire N__14490;
    wire N__14489;
    wire N__14488;
    wire N__14487;
    wire N__14486;
    wire N__14485;
    wire N__14484;
    wire N__14469;
    wire N__14468;
    wire N__14467;
    wire N__14466;
    wire N__14465;
    wire N__14464;
    wire N__14463;
    wire N__14462;
    wire N__14461;
    wire N__14460;
    wire N__14459;
    wire N__14458;
    wire N__14457;
    wire N__14456;
    wire N__14455;
    wire N__14454;
    wire N__14451;
    wire N__14448;
    wire N__14447;
    wire N__14446;
    wire N__14445;
    wire N__14444;
    wire N__14431;
    wire N__14430;
    wire N__14429;
    wire N__14428;
    wire N__14427;
    wire N__14426;
    wire N__14425;
    wire N__14424;
    wire N__14423;
    wire N__14422;
    wire N__14421;
    wire N__14420;
    wire N__14419;
    wire N__14418;
    wire N__14417;
    wire N__14416;
    wire N__14415;
    wire N__14414;
    wire N__14413;
    wire N__14412;
    wire N__14411;
    wire N__14410;
    wire N__14409;
    wire N__14408;
    wire N__14407;
    wire N__14406;
    wire N__14405;
    wire N__14404;
    wire N__14403;
    wire N__14388;
    wire N__14387;
    wire N__14386;
    wire N__14385;
    wire N__14384;
    wire N__14383;
    wire N__14382;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14360;
    wire N__14357;
    wire N__14342;
    wire N__14339;
    wire N__14338;
    wire N__14337;
    wire N__14336;
    wire N__14335;
    wire N__14334;
    wire N__14333;
    wire N__14330;
    wire N__14315;
    wire N__14300;
    wire N__14295;
    wire N__14286;
    wire N__14283;
    wire N__14268;
    wire N__14253;
    wire N__14252;
    wire N__14251;
    wire N__14250;
    wire N__14249;
    wire N__14248;
    wire N__14247;
    wire N__14246;
    wire N__14245;
    wire N__14244;
    wire N__14243;
    wire N__14242;
    wire N__14241;
    wire N__14240;
    wire N__14239;
    wire N__14238;
    wire N__14237;
    wire N__14236;
    wire N__14235;
    wire N__14234;
    wire N__14233;
    wire N__14232;
    wire N__14217;
    wire N__14202;
    wire N__14199;
    wire N__14184;
    wire N__14179;
    wire N__14174;
    wire N__14171;
    wire N__14168;
    wire N__14155;
    wire N__14148;
    wire N__14137;
    wire N__14136;
    wire N__14135;
    wire N__14134;
    wire N__14119;
    wire N__14104;
    wire N__14089;
    wire N__14082;
    wire N__14075;
    wire N__14070;
    wire N__14063;
    wire N__14056;
    wire N__14039;
    wire N__14038;
    wire N__14035;
    wire N__14030;
    wire N__14027;
    wire N__14026;
    wire N__14021;
    wire N__14018;
    wire N__14017;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14005;
    wire N__14000;
    wire N__13997;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13985;
    wire N__13982;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13964;
    wire N__13961;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13949;
    wire N__13946;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13934;
    wire N__13933;
    wire N__13932;
    wire N__13931;
    wire N__13930;
    wire N__13929;
    wire N__13928;
    wire N__13927;
    wire N__13926;
    wire N__13925;
    wire N__13924;
    wire N__13923;
    wire N__13922;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13911;
    wire N__13910;
    wire N__13909;
    wire N__13908;
    wire N__13907;
    wire N__13906;
    wire N__13905;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13894;
    wire N__13893;
    wire N__13892;
    wire N__13891;
    wire N__13890;
    wire N__13889;
    wire N__13888;
    wire N__13887;
    wire N__13886;
    wire N__13885;
    wire N__13884;
    wire N__13883;
    wire N__13882;
    wire N__13881;
    wire N__13880;
    wire N__13879;
    wire N__13878;
    wire N__13877;
    wire N__13876;
    wire N__13875;
    wire N__13874;
    wire N__13873;
    wire N__13872;
    wire N__13871;
    wire N__13870;
    wire N__13867;
    wire N__13864;
    wire N__13861;
    wire N__13860;
    wire N__13859;
    wire N__13858;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13847;
    wire N__13846;
    wire N__13843;
    wire N__13842;
    wire N__13841;
    wire N__13840;
    wire N__13839;
    wire N__13838;
    wire N__13837;
    wire N__13836;
    wire N__13821;
    wire N__13818;
    wire N__13817;
    wire N__13816;
    wire N__13815;
    wire N__13814;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13803;
    wire N__13802;
    wire N__13801;
    wire N__13800;
    wire N__13785;
    wire N__13784;
    wire N__13783;
    wire N__13782;
    wire N__13781;
    wire N__13780;
    wire N__13779;
    wire N__13772;
    wire N__13771;
    wire N__13770;
    wire N__13769;
    wire N__13768;
    wire N__13767;
    wire N__13764;
    wire N__13761;
    wire N__13758;
    wire N__13757;
    wire N__13756;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13747;
    wire N__13746;
    wire N__13745;
    wire N__13730;
    wire N__13729;
    wire N__13728;
    wire N__13727;
    wire N__13726;
    wire N__13725;
    wire N__13724;
    wire N__13723;
    wire N__13722;
    wire N__13721;
    wire N__13720;
    wire N__13719;
    wire N__13716;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13705;
    wire N__13704;
    wire N__13703;
    wire N__13696;
    wire N__13683;
    wire N__13670;
    wire N__13667;
    wire N__13660;
    wire N__13651;
    wire N__13646;
    wire N__13645;
    wire N__13644;
    wire N__13643;
    wire N__13642;
    wire N__13641;
    wire N__13640;
    wire N__13639;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13619;
    wire N__13610;
    wire N__13607;
    wire N__13594;
    wire N__13591;
    wire N__13582;
    wire N__13567;
    wire N__13554;
    wire N__13551;
    wire N__13548;
    wire N__13545;
    wire N__13542;
    wire N__13539;
    wire N__13538;
    wire N__13537;
    wire N__13536;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13526;
    wire N__13525;
    wire N__13524;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13513;
    wire N__13512;
    wire N__13511;
    wire N__13508;
    wire N__13507;
    wire N__13506;
    wire N__13505;
    wire N__13504;
    wire N__13503;
    wire N__13502;
    wire N__13501;
    wire N__13500;
    wire N__13497;
    wire N__13482;
    wire N__13473;
    wire N__13466;
    wire N__13463;
    wire N__13448;
    wire N__13443;
    wire N__13436;
    wire N__13433;
    wire N__13426;
    wire N__13421;
    wire N__13406;
    wire N__13393;
    wire N__13378;
    wire N__13373;
    wire N__13358;
    wire N__13351;
    wire N__13348;
    wire N__13339;
    wire N__13332;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13273;
    wire N__13268;
    wire N__13265;
    wire N__13264;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13130;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13037;
    wire N__13034;
    wire N__13031;
    wire N__13028;
    wire N__13025;
    wire N__13022;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13009;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12967;
    wire N__12964;
    wire N__12961;
    wire N__12958;
    wire N__12953;
    wire N__12950;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12940;
    wire N__12937;
    wire N__12934;
    wire N__12931;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12919;
    wire N__12916;
    wire N__12913;
    wire N__12910;
    wire N__12907;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12895;
    wire N__12890;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12877;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12865;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12847;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12835;
    wire N__12830;
    wire N__12827;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12817;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12805;
    wire N__12802;
    wire N__12799;
    wire N__12796;
    wire N__12791;
    wire N__12790;
    wire N__12785;
    wire N__12782;
    wire N__12781;
    wire N__12778;
    wire N__12775;
    wire N__12770;
    wire N__12767;
    wire N__12766;
    wire N__12761;
    wire N__12758;
    wire N__12757;
    wire N__12752;
    wire N__12749;
    wire N__12748;
    wire N__12743;
    wire N__12740;
    wire N__12739;
    wire N__12736;
    wire N__12733;
    wire N__12730;
    wire N__12725;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12713;
    wire N__12712;
    wire N__12707;
    wire N__12704;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12689;
    wire N__12688;
    wire N__12683;
    wire N__12680;
    wire N__12679;
    wire N__12676;
    wire N__12673;
    wire N__12668;
    wire N__12667;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12653;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12643;
    wire N__12640;
    wire N__12635;
    wire N__12634;
    wire N__12631;
    wire N__12628;
    wire N__12623;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12608;
    wire N__12607;
    wire N__12604;
    wire N__12601;
    wire N__12596;
    wire N__12593;
    wire N__12592;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12580;
    wire N__12577;
    wire N__12572;
    wire N__12569;
    wire N__12568;
    wire N__12563;
    wire N__12560;
    wire N__12559;
    wire N__12554;
    wire N__12551;
    wire N__12550;
    wire N__12545;
    wire N__12542;
    wire N__12541;
    wire N__12538;
    wire N__12535;
    wire N__12530;
    wire N__12529;
    wire N__12524;
    wire N__12521;
    wire N__12520;
    wire N__12515;
    wire N__12512;
    wire N__12511;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12499;
    wire N__12496;
    wire N__12493;
    wire N__12490;
    wire N__12485;
    wire N__12484;
    wire N__12481;
    wire N__12478;
    wire N__12473;
    wire N__12470;
    wire N__12469;
    wire N__12466;
    wire N__12463;
    wire N__12458;
    wire N__12455;
    wire N__12454;
    wire N__12451;
    wire N__12448;
    wire N__12443;
    wire N__12442;
    wire N__12439;
    wire N__12434;
    wire N__12431;
    wire N__12430;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12364;
    wire N__12361;
    wire N__12358;
    wire N__12355;
    wire N__12352;
    wire N__12347;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12332;
    wire N__12329;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12271;
    wire N__12270;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12256;
    wire N__12255;
    wire N__12252;
    wire N__12247;
    wire N__12242;
    wire N__12241;
    wire N__12240;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12232;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12210;
    wire N__12207;
    wire N__12206;
    wire N__12203;
    wire N__12198;
    wire N__12195;
    wire N__12192;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12154;
    wire N__12153;
    wire N__12152;
    wire N__12151;
    wire N__12144;
    wire N__12139;
    wire N__12136;
    wire N__12131;
    wire N__12130;
    wire N__12129;
    wire N__12128;
    wire N__12121;
    wire N__12118;
    wire N__12115;
    wire N__12110;
    wire N__12109;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12097;
    wire N__12092;
    wire N__12089;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12077;
    wire N__12074;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12062;
    wire N__12061;
    wire N__12058;
    wire N__12055;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12037;
    wire N__12034;
    wire N__12031;
    wire N__12026;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12014;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11957;
    wire N__11954;
    wire N__11953;
    wire N__11950;
    wire N__11947;
    wire N__11942;
    wire N__11939;
    wire N__11938;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11926;
    wire N__11921;
    wire N__11918;
    wire N__11917;
    wire N__11912;
    wire N__11909;
    wire N__11908;
    wire N__11905;
    wire N__11900;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11881;
    wire N__11876;
    wire N__11873;
    wire N__11872;
    wire N__11867;
    wire N__11864;
    wire N__11863;
    wire N__11858;
    wire N__11855;
    wire N__11854;
    wire N__11851;
    wire N__11846;
    wire N__11843;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11831;
    wire N__11828;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11813;
    wire N__11810;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11789;
    wire N__11788;
    wire N__11783;
    wire N__11780;
    wire N__11779;
    wire N__11774;
    wire N__11771;
    wire N__11770;
    wire N__11767;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11744;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11729;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11717;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11705;
    wire N__11702;
    wire N__11701;
    wire N__11696;
    wire N__11693;
    wire N__11692;
    wire N__11687;
    wire N__11684;
    wire N__11683;
    wire N__11678;
    wire N__11675;
    wire N__11674;
    wire N__11671;
    wire N__11666;
    wire N__11663;
    wire N__11662;
    wire N__11657;
    wire N__11654;
    wire N__11653;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11630;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11609;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11560;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11488;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11470;
    wire N__11469;
    wire N__11468;
    wire N__11465;
    wire N__11462;
    wire N__11457;
    wire N__11450;
    wire N__11449;
    wire N__11448;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11435;
    wire N__11430;
    wire N__11423;
    wire N__11422;
    wire N__11421;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11409;
    wire N__11402;
    wire N__11401;
    wire N__11400;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11388;
    wire N__11381;
    wire N__11380;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11363;
    wire N__11360;
    wire N__11359;
    wire N__11358;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11346;
    wire N__11339;
    wire N__11336;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11324;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11316;
    wire N__11313;
    wire N__11308;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11272;
    wire N__11267;
    wire N__11264;
    wire N__11263;
    wire N__11262;
    wire N__11259;
    wire N__11252;
    wire N__11249;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11231;
    wire N__11228;
    wire N__11227;
    wire N__11222;
    wire N__11219;
    wire N__11218;
    wire N__11213;
    wire N__11210;
    wire N__11209;
    wire N__11204;
    wire N__11201;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11189;
    wire N__11186;
    wire N__11185;
    wire N__11182;
    wire N__11177;
    wire N__11174;
    wire N__11173;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11144;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11126;
    wire N__11123;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11108;
    wire N__11105;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11093;
    wire N__11090;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11075;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11063;
    wire N__11060;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11026;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10970;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10958;
    wire N__10955;
    wire N__10954;
    wire N__10951;
    wire N__10948;
    wire N__10943;
    wire N__10942;
    wire N__10937;
    wire N__10934;
    wire N__10933;
    wire N__10928;
    wire N__10925;
    wire N__10924;
    wire N__10921;
    wire N__10918;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10906;
    wire N__10901;
    wire N__10898;
    wire N__10897;
    wire N__10892;
    wire N__10889;
    wire N__10888;
    wire N__10883;
    wire N__10880;
    wire N__10879;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10867;
    wire N__10864;
    wire N__10861;
    wire N__10856;
    wire N__10853;
    wire N__10852;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10840;
    wire N__10835;
    wire N__10832;
    wire N__10831;
    wire N__10826;
    wire N__10823;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10777;
    wire N__10772;
    wire N__10769;
    wire N__10768;
    wire N__10765;
    wire N__10762;
    wire N__10759;
    wire N__10754;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10684;
    wire N__10681;
    wire N__10678;
    wire N__10673;
    wire N__10672;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10658;
    wire N__10657;
    wire N__10654;
    wire N__10651;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10612;
    wire N__10609;
    wire N__10606;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10562;
    wire N__10559;
    wire N__10558;
    wire N__10555;
    wire N__10552;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10528;
    wire N__10525;
    wire N__10522;
    wire N__10519;
    wire N__10514;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10499;
    wire N__10496;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10481;
    wire N__10480;
    wire N__10477;
    wire N__10474;
    wire N__10471;
    wire N__10466;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10451;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10441;
    wire N__10436;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10421;
    wire N__10420;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10406;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10378;
    wire N__10373;
    wire N__10370;
    wire N__10369;
    wire N__10366;
    wire N__10361;
    wire N__10358;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10313;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10294;
    wire N__10289;
    wire N__10286;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10268;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10256;
    wire N__10253;
    wire N__10252;
    wire N__10247;
    wire N__10244;
    wire N__10243;
    wire N__10238;
    wire N__10235;
    wire N__10234;
    wire N__10229;
    wire N__10226;
    wire N__10225;
    wire N__10220;
    wire N__10217;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10198;
    wire N__10193;
    wire N__10190;
    wire N__10189;
    wire N__10184;
    wire N__10181;
    wire N__10180;
    wire N__10177;
    wire N__10174;
    wire N__10169;
    wire N__10168;
    wire N__10163;
    wire N__10160;
    wire N__10159;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10136;
    wire N__10135;
    wire N__10130;
    wire VCCG0;
    wire \tok.A_stk.tail_89 ;
    wire \tok.A_stk.tail_73 ;
    wire \tok.A_stk.tail_57 ;
    wire \tok.A_stk.tail_41 ;
    wire \tok.A_stk.tail_25 ;
    wire \tok.A_stk.tail_9 ;
    wire \tok.A_stk.tail_87 ;
    wire \tok.A_stk.tail_71 ;
    wire \tok.A_stk.tail_55 ;
    wire \tok.A_stk.tail_39 ;
    wire \tok.A_stk.tail_23 ;
    wire \tok.A_stk.tail_7 ;
    wire tail_123;
    wire tail_107;
    wire \tok.A_stk.tail_91 ;
    wire \tok.A_stk.tail_75 ;
    wire \tok.A_stk.tail_59 ;
    wire \tok.A_stk.tail_43 ;
    wire \tok.A_stk.tail_27 ;
    wire \tok.A_stk.tail_11 ;
    wire bfn_1_5_0_;
    wire \tok.uart.n3955 ;
    wire \tok.uart.n3956 ;
    wire \tok.uart.n3957 ;
    wire \tok.uart.n3958 ;
    wire \tok.uart.n3959 ;
    wire \tok.uart.n3960 ;
    wire \tok.uart.n3961 ;
    wire \tok.uart.n3962 ;
    wire bfn_1_6_0_;
    wire \tok.uart.txclkcounter_3 ;
    wire \tok.uart.txclkcounter_5 ;
    wire \tok.uart.txclkcounter_0 ;
    wire \tok.uart.txclkcounter_2 ;
    wire \tok.uart.txclkcounter_6 ;
    wire \tok.uart.txclkcounter_1 ;
    wire \tok.uart.txclkcounter_7 ;
    wire \tok.uart.txclkcounter_8 ;
    wire \tok.uart.txclkcounter_4 ;
    wire \tok.uart.n14_cascade_ ;
    wire \tok.uart.n15_adj_640 ;
    wire txtick_cascade_;
    wire \tok.uart.n1081 ;
    wire \tok.uart.rxclkcounter_0 ;
    wire bfn_1_8_0_;
    wire \tok.uart.rxclkcounter_1 ;
    wire \tok.uart.n3968 ;
    wire \tok.uart.n3969 ;
    wire \tok.uart.rxclkcounter_3 ;
    wire \tok.uart.n3970 ;
    wire \tok.uart.rxclkcounter_4 ;
    wire \tok.uart.n3971 ;
    wire \tok.uart.n3972 ;
    wire \tok.uart.n3973 ;
    wire \tok.table_wr_data_8 ;
    wire \tok.table_wr_data_15 ;
    wire \tok.table_wr_data_14 ;
    wire \tok.table_wr_data_13 ;
    wire \tok.uart.n12 ;
    wire \tok.uart.rxclkcounter_6 ;
    wire \tok.uart.rxclkcounter_5 ;
    wire \tok.uart.rxclkcounter_2 ;
    wire n795_cascade_;
    wire \tok.table_wr_data_9 ;
    wire bfn_1_10_0_;
    wire \tok.uart.n3963 ;
    wire \tok.uart.n3964 ;
    wire \tok.uart.n3965 ;
    wire \tok.uart.n3966 ;
    wire \tok.uart.n3967 ;
    wire n940;
    wire \tok.A_stk.tail_16 ;
    wire \tok.A_stk.tail_32 ;
    wire \tok.A_stk.tail_48 ;
    wire \tok.A_stk.tail_64 ;
    wire \tok.A_stk.tail_80 ;
    wire \tok.A_stk.tail_0 ;
    wire \tok.A_stk.tail_94 ;
    wire \tok.A_stk.tail_78 ;
    wire \tok.A_stk.tail_62 ;
    wire \tok.A_stk.tail_46 ;
    wire \tok.A_stk.tail_30 ;
    wire \tok.A_stk.tail_14 ;
    wire \tok.A_stk.tail_88 ;
    wire \tok.A_stk.tail_72 ;
    wire \tok.A_stk.tail_56 ;
    wire \tok.A_stk.tail_40 ;
    wire \tok.A_stk.tail_24 ;
    wire \tok.A_stk.tail_8 ;
    wire tail_96;
    wire tail_112;
    wire tail_105;
    wire tail_121;
    wire tail_104;
    wire tail_120;
    wire tail_103;
    wire tail_119;
    wire \tok.table_wr_data_12 ;
    wire tail_122;
    wire tail_106;
    wire \tok.A_stk.tail_90 ;
    wire \tok.A_stk.tail_74 ;
    wire \tok.A_stk.tail_58 ;
    wire \tok.A_stk.tail_42 ;
    wire \tok.A_stk.tail_26 ;
    wire \tok.A_stk.tail_10 ;
    wire \tok.n2_adj_763 ;
    wire \tok.n13_adj_765_cascade_ ;
    wire \tok.n18_adj_767_cascade_ ;
    wire \tok.n20_adj_770_cascade_ ;
    wire \tok.A_15_N_113_7_cascade_ ;
    wire \tok.A_15_N_84_7 ;
    wire \tok.A_15_N_113_7 ;
    wire \tok.uart.sentbits_3 ;
    wire \tok.uart.sentbits_2 ;
    wire \tok.uart.n3994_cascade_ ;
    wire n795;
    wire \tok.uart.n4506_cascade_ ;
    wire \tok.uart.rxclkcounter_6__N_477 ;
    wire \tok.uart.n4438 ;
    wire \tok.uart.n2 ;
    wire \tok.n16_adj_769 ;
    wire \tok.uart.bytephase_1 ;
    wire \tok.uart.bytephase_5 ;
    wire \tok.uart.bytephase_3 ;
    wire \tok.uart.bytephase_0 ;
    wire \tok.uart.bytephase_2 ;
    wire \tok.uart.n13_cascade_ ;
    wire \tok.uart.bytephase_4 ;
    wire bytephase_5__N_510;
    wire rx_c;
    wire capture_9;
    wire \tok.n4508_cascade_ ;
    wire \tok.n4680 ;
    wire \tok.n16_adj_660_cascade_ ;
    wire \tok.n4 ;
    wire \tok.n206_cascade_ ;
    wire \tok.n204_cascade_ ;
    wire \tok.n16_adj_699_cascade_ ;
    wire \tok.n4667 ;
    wire \tok.A_stk.tail_18 ;
    wire \tok.A_stk.tail_34 ;
    wire \tok.A_stk.tail_50 ;
    wire \tok.A_stk.tail_66 ;
    wire \tok.A_stk.tail_82 ;
    wire \tok.A_stk.tail_2 ;
    wire tail_110;
    wire tail_126;
    wire tail_98;
    wire tail_114;
    wire tail_125;
    wire tail_109;
    wire \tok.A_stk.tail_93 ;
    wire \tok.A_stk.tail_77 ;
    wire \tok.A_stk.tail_61 ;
    wire \tok.A_stk.tail_45 ;
    wire \tok.A_stk.tail_29 ;
    wire \tok.A_stk.tail_13 ;
    wire tail_118;
    wire tail_102;
    wire \tok.A_stk.tail_86 ;
    wire \tok.A_stk.tail_70 ;
    wire \tok.A_stk.tail_54 ;
    wire \tok.A_stk.tail_38 ;
    wire \tok.A_stk.tail_22 ;
    wire \tok.A_stk.tail_6 ;
    wire \tok.n20_adj_803_cascade_ ;
    wire \tok.key_rd_5 ;
    wire \tok.key_rd_3 ;
    wire \tok.key_rd_8 ;
    wire \tok.n28 ;
    wire \tok.n25_cascade_ ;
    wire \tok.n26 ;
    wire \tok.key_rd_14 ;
    wire \tok.key_rd_11 ;
    wire \tok.table_wr_data_11 ;
    wire \tok.key_rd_15 ;
    wire \tok.key_rd_9 ;
    wire \tok.table_wr_data_7 ;
    wire \tok.table_wr_data_4 ;
    wire \tok.table_wr_data_1 ;
    wire \tok.n15_adj_771 ;
    wire \tok.uart.n6_cascade_ ;
    wire n23_cascade_;
    wire \tok.uart.sentbits_0 ;
    wire \tok.uart.sentbits_1 ;
    wire \tok.uart.n978 ;
    wire \tok.uart.n1083 ;
    wire capture_7;
    wire capture_6;
    wire txtick;
    wire bfn_4_11_0_;
    wire \tok.n3910 ;
    wire \tok.n300 ;
    wire \tok.n3911 ;
    wire \tok.n3912 ;
    wire \tok.n3913 ;
    wire \tok.n3914 ;
    wire \tok.n3915 ;
    wire \tok.n295 ;
    wire \tok.n6_adj_768 ;
    wire \tok.n3916 ;
    wire \tok.n3917 ;
    wire bfn_4_12_0_;
    wire \tok.n3918 ;
    wire \tok.n3919 ;
    wire \tok.n291 ;
    wire \tok.n3920 ;
    wire \tok.n290 ;
    wire \tok.n6_adj_701 ;
    wire \tok.n3921 ;
    wire \tok.n3922 ;
    wire \tok.n288 ;
    wire \tok.n3923 ;
    wire GNDG0;
    wire \tok.n3924 ;
    wire \tok.n3924_THRU_CRY_0_THRU_CO ;
    wire bfn_4_13_0_;
    wire \tok.n292 ;
    wire \tok.n287 ;
    wire tail_124;
    wire tail_108;
    wire \tok.A_stk.tail_92 ;
    wire \tok.A_stk.tail_76 ;
    wire \tok.A_stk.tail_60 ;
    wire \tok.A_stk.tail_44 ;
    wire \tok.A_stk.tail_28 ;
    wire \tok.A_stk.tail_12 ;
    wire \tok.A_stk.tail_17 ;
    wire \tok.A_stk.tail_33 ;
    wire \tok.A_stk.tail_49 ;
    wire \tok.A_stk.tail_65 ;
    wire \tok.A_stk.tail_81 ;
    wire \tok.A_stk.tail_1 ;
    wire tail_115;
    wire \tok.A_stk.tail_51 ;
    wire tail_117;
    wire tail_101;
    wire \tok.A_stk.tail_67 ;
    wire tail_99;
    wire \tok.A_stk.tail_83 ;
    wire \tok.A_stk.tail_35 ;
    wire \tok.A_stk.tail_3 ;
    wire \tok.A_stk.tail_19 ;
    wire \tok.A_stk.tail_85 ;
    wire \tok.A_stk.tail_69 ;
    wire \tok.A_stk.tail_53 ;
    wire \tok.A_stk.tail_37 ;
    wire \tok.A_stk.tail_21 ;
    wire \tok.A_stk.tail_5 ;
    wire tail_116;
    wire tail_100;
    wire \tok.A_stk.tail_84 ;
    wire \tok.A_stk.tail_68 ;
    wire \tok.A_stk.tail_52 ;
    wire \tok.A_stk.tail_36 ;
    wire \tok.A_stk.tail_20 ;
    wire \tok.A_stk.tail_4 ;
    wire \tok.n23_adj_677 ;
    wire \tok.n24 ;
    wire \tok.n26_adj_805 ;
    wire \tok.n30_adj_824_cascade_ ;
    wire \tok.found_slot_N_145 ;
    wire \tok.n4642_cascade_ ;
    wire \tok.key_rd_13 ;
    wire \tok.n14_adj_804 ;
    wire \tok.n27_adj_734 ;
    wire \tok.key_rd_12 ;
    wire \tok.key_rd_10 ;
    wire \tok.n21_adj_714 ;
    wire \tok.key_rd_2 ;
    wire \tok.key_rd_7 ;
    wire \tok.n22 ;
    wire bfn_5_8_0_;
    wire \tok.n3940 ;
    wire \tok.n3941 ;
    wire \tok.n3942 ;
    wire \tok.n3943 ;
    wire \tok.n3944 ;
    wire \tok.n3945 ;
    wire \tok.n10_adj_764 ;
    wire \tok.n3946 ;
    wire \tok.n3947 ;
    wire bfn_5_9_0_;
    wire \tok.n3948 ;
    wire \tok.n3949 ;
    wire \tok.n3950 ;
    wire \tok.n3951 ;
    wire \tok.n3952 ;
    wire \tok.n3953 ;
    wire \tok.n3954 ;
    wire \tok.n2_adj_739_cascade_ ;
    wire \tok.n6_adj_753 ;
    wire \tok.n14_adj_741_cascade_ ;
    wire \tok.n13_adj_748 ;
    wire \tok.n4656 ;
    wire \tok.n20_adj_754_cascade_ ;
    wire \tok.n9_adj_749 ;
    wire \tok.table_rd_15 ;
    wire \tok.n16_adj_751 ;
    wire \tok.n17_adj_774 ;
    wire \tok.n10_adj_705 ;
    wire \tok.n6_adj_692 ;
    wire \tok.n13_adj_688_cascade_ ;
    wire \tok.n12_adj_687 ;
    wire \tok.n4674 ;
    wire \tok.n20_adj_693_cascade_ ;
    wire \tok.n6_adj_667 ;
    wire \tok.n294 ;
    wire \tok.table_wr_data_3 ;
    wire \tok.n298 ;
    wire \tok.n289 ;
    wire \tok.n6_adj_814 ;
    wire \tok.n34_cascade_ ;
    wire \tok.n13 ;
    wire \tok.n2_adj_685_cascade_ ;
    wire \tok.n14_adj_686 ;
    wire sender_1;
    wire tx_c;
    wire reset_c;
    wire \tok.A_stk.tail_63 ;
    wire \tok.A_stk.tail_47 ;
    wire \tok.A_stk.tail_31 ;
    wire \tok.A_stk.tail_15 ;
    wire \tok.A_stk.tail_79 ;
    wire \tok.A_stk.tail_95 ;
    wire tail_111;
    wire tail_127;
    wire tail_97;
    wire tail_113;
    wire n29;
    wire n29_cascade_;
    wire \tok.A_stk.rd_15__N_301 ;
    wire \tok.n83_adj_735_cascade_ ;
    wire \tok.n7_cascade_ ;
    wire \tok.n4516 ;
    wire capture_0;
    wire \tok.n17 ;
    wire \tok.n4_adj_654_cascade_ ;
    wire n786;
    wire \tok.n83_adj_716_cascade_ ;
    wire \tok.n12_adj_740_cascade_ ;
    wire \tok.n12_adj_801_cascade_ ;
    wire \tok.n284 ;
    wire \tok.n284_cascade_ ;
    wire \tok.n182_cascade_ ;
    wire \tok.n12_adj_766 ;
    wire \tok.n24_adj_854 ;
    wire \tok.n21_adj_857 ;
    wire \tok.n30_adj_862_cascade_ ;
    wire \tok.n19_adj_860_cascade_ ;
    wire \tok.n17_adj_861 ;
    wire \tok.n29_adj_864 ;
    wire capture_8;
    wire uart_rx_data_7;
    wire \tok.table_wr_data_10 ;
    wire \tok.n293 ;
    wire \tok.n2634 ;
    wire \tok.write_slot ;
    wire \tok.table_wr_data_5 ;
    wire \tok.key_rd_4 ;
    wire \tok.key_rd_1 ;
    wire \tok.n18_adj_756 ;
    wire \tok.key_rd_0 ;
    wire \tok.key_rd_6 ;
    wire \tok.n4645 ;
    wire \tok.n13_adj_657 ;
    wire \tok.n10_adj_656 ;
    wire \tok.table_rd_9 ;
    wire \tok.n30_cascade_ ;
    wire \tok.n12_adj_659 ;
    wire \tok.uart.n922 ;
    wire \tok.n301 ;
    wire \tok.n15_cascade_ ;
    wire \tok.n183 ;
    wire \tok.table_rd_6 ;
    wire \tok.n16_adj_778_cascade_ ;
    wire \tok.n6_adj_780 ;
    wire \tok.table_rd_13 ;
    wire \tok.table_rd_10 ;
    wire \tok.n10_adj_671 ;
    wire \tok.n14_adj_669_cascade_ ;
    wire \tok.table_rd_11 ;
    wire \tok.n16_adj_691 ;
    wire \tok.n4653 ;
    wire \tok.n4671 ;
    wire \tok.n18_adj_672 ;
    wire \tok.n6_adj_676 ;
    wire \tok.n20_adj_674_cascade_ ;
    wire \tok.n16_adj_673 ;
    wire \tok.n4676_cascade_ ;
    wire \tok.n12_adj_744 ;
    wire \tok.n4524 ;
    wire \tok.n12_adj_670 ;
    wire \tok.n2_adj_720_cascade_ ;
    wire \tok.n14_adj_722 ;
    wire \tok.n6_adj_731 ;
    wire \tok.n13_adj_726_cascade_ ;
    wire \tok.n12_adj_723 ;
    wire \tok.n4661 ;
    wire \tok.n20_adj_732_cascade_ ;
    wire \tok.n4658 ;
    wire \tok.n9_adj_728 ;
    wire \tok.n184 ;
    wire uart_rx_data_5;
    wire \tok.n12_adj_815_cascade_ ;
    wire \tok.n16_adj_820 ;
    wire \tok.n20_adj_822_cascade_ ;
    wire \tok.A_15_N_113_5_cascade_ ;
    wire \tok.n297 ;
    wire \tok.n208 ;
    wire \tok.n20_adj_858 ;
    wire \tok.n299 ;
    wire \tok.n27_adj_644_cascade_ ;
    wire \tok.tail_9 ;
    wire \tok.C_stk.tail_17 ;
    wire \tok.tail_25 ;
    wire \tok.C_stk.tail_33 ;
    wire \tok.tail_57 ;
    wire \tok.tail_41 ;
    wire \tok.tail_49 ;
    wire \tok.tail_58 ;
    wire \tok.n875_cascade_ ;
    wire \tok.n2562 ;
    wire \tok.n2503 ;
    wire \tok.n2562_cascade_ ;
    wire \tok.n4474_cascade_ ;
    wire \tok.n875 ;
    wire \tok.n20_adj_772_cascade_ ;
    wire \tok.n63 ;
    wire \tok.A_stk_delta_1__N_4_cascade_ ;
    wire \tok.n61 ;
    wire \tok.n4_adj_809_cascade_ ;
    wire \tok.depth_3_cascade_ ;
    wire \tok.depth_1 ;
    wire \tok.n4554_cascade_ ;
    wire \tok.n237 ;
    wire \tok.n6_adj_832 ;
    wire \tok.n4504 ;
    wire \tok.n4432_cascade_ ;
    wire \tok.A_stk_delta_1__N_4 ;
    wire \tok.n1_adj_802_cascade_ ;
    wire \tok.n189 ;
    wire \tok.n62 ;
    wire \tok.n189_cascade_ ;
    wire \tok.n4_adj_809 ;
    wire \tok.n27_adj_793_cascade_ ;
    wire \tok.n25_adj_794 ;
    wire \tok.n26_adj_792 ;
    wire \tok.n28_adj_791 ;
    wire \tok.n18_adj_859 ;
    wire \tok.n22_adj_855 ;
    wire \tok.n880 ;
    wire \tok.n23_cascade_ ;
    wire \tok.n23_adj_856 ;
    wire \tok.n64 ;
    wire \tok.n1_adj_802 ;
    wire \tok.depth_2 ;
    wire \tok.depth_0_cascade_ ;
    wire \tok.n6_adj_853 ;
    wire \tok.A__15__N_129_cascade_ ;
    wire \tok.n27_adj_867_cascade_ ;
    wire \tok.n1 ;
    wire \tok.n14_adj_678_cascade_ ;
    wire \tok.n2 ;
    wire \tok.n19_cascade_ ;
    wire \tok.n6_adj_684 ;
    wire \tok.n22_adj_683_cascade_ ;
    wire \tok.n4544 ;
    wire \tok.A_15_N_113_0_cascade_ ;
    wire \tok.n4520 ;
    wire \tok.n46_cascade_ ;
    wire \tok.A_15_N_113_1 ;
    wire \tok.A_15_N_113_1_cascade_ ;
    wire \tok.A_1_cascade_ ;
    wire \tok.uart.sender_3 ;
    wire \tok.A_0 ;
    wire sender_2;
    wire \tok.A_2 ;
    wire \tok.uart.sender_4 ;
    wire \tok.n10_adj_783 ;
    wire \tok.n14_adj_779_cascade_ ;
    wire \tok.n20_adj_781 ;
    wire \tok.n22_adj_784_cascade_ ;
    wire \tok.A_15_N_113_6_cascade_ ;
    wire \tok.A_6_cascade_ ;
    wire \tok.uart.sender_9 ;
    wire \tok.uart.sender_8 ;
    wire \tok.A_5 ;
    wire \tok.uart.sender_7 ;
    wire \tok.uart.sender_6 ;
    wire n23;
    wire \tok.uart.sender_5 ;
    wire \tok.uart.n964 ;
    wire \tok.n16_adj_706 ;
    wire \tok.n14_adj_707 ;
    wire \tok.n20_adj_708_cascade_ ;
    wire \tok.n22_adj_709_cascade_ ;
    wire \tok.A_15_N_113_5 ;
    wire \tok.n10_adj_806 ;
    wire \tok.n13_adj_813_cascade_ ;
    wire \tok.n18_adj_819 ;
    wire \tok.n15_adj_823 ;
    wire \tok.n27_adj_863_cascade_ ;
    wire \tok.n27_adj_865_cascade_ ;
    wire \tok.n27_adj_664 ;
    wire \tok.n27_adj_866 ;
    wire \tok.tail_50 ;
    wire \tok.C_stk.tail_34 ;
    wire \tok.tail_42 ;
    wire \tok.tail_28 ;
    wire \tok.n127_cascade_ ;
    wire \tok.n4446 ;
    wire \tok.n4394_cascade_ ;
    wire \tok.n28_adj_834_cascade_ ;
    wire \tok.n4604_cascade_ ;
    wire \tok.n34_adj_719 ;
    wire \tok.n4610_cascade_ ;
    wire \tok.n37 ;
    wire \tok.table_rd_7 ;
    wire \tok.n83_adj_796_cascade_ ;
    wire capture_3;
    wire \tok.n847 ;
    wire \tok.n31 ;
    wire \tok.C_stk.n4906_cascade_ ;
    wire \tok.ram.n4699_cascade_ ;
    wire \tok.n4649 ;
    wire \tok.n1_adj_760_cascade_ ;
    wire \tok.n13_adj_761_cascade_ ;
    wire \tok.tc_7 ;
    wire \tok.C_stk.tail_1 ;
    wire \tok.C_stk.n4870_cascade_ ;
    wire \tok.ram.n4714_cascade_ ;
    wire \tok.c_stk_r_1 ;
    wire \tok.n4690 ;
    wire \tok.n1_adj_717_cascade_ ;
    wire \tok.n5_adj_718_cascade_ ;
    wire n92_cascade_;
    wire \tok.tc_1 ;
    wire \tok.n28_adj_821 ;
    wire \tok.n10_adj_786 ;
    wire \tok.n6_adj_848_cascade_ ;
    wire \tok.n32_cascade_ ;
    wire uart_rx_data_1;
    wire \tok.table_wr_data_6 ;
    wire capture_2;
    wire n4005;
    wire \tok.table_wr_data_2 ;
    wire \tok.n18_adj_844_cascade_ ;
    wire \tok.n16_adj_845 ;
    wire \tok.n20_adj_846_cascade_ ;
    wire \tok.A_15_N_113_2 ;
    wire \tok.n15_adj_847 ;
    wire uart_rx_data_2;
    wire \tok.n12_adj_843 ;
    wire capture_1;
    wire uart_rx_data_0;
    wire \tok.table_rd_14 ;
    wire \tok.n16_adj_730 ;
    wire \tok.n400 ;
    wire \tok.table_wr_data_0 ;
    wire \tok.n2614 ;
    wire \tok.n2614_cascade_ ;
    wire \tok.n2616_cascade_ ;
    wire \tok.n10_adj_849 ;
    wire \tok.n12_adj_851 ;
    wire \tok.table_rd_1 ;
    wire \tok.n8_adj_850 ;
    wire \tok.A_4 ;
    wire \tok.n4051 ;
    wire \tok.A_15_N_113_4 ;
    wire \tok.A_15_N_113_4_cascade_ ;
    wire \tok.A_15_N_113_0 ;
    wire \tok.A_15_N_113_6 ;
    wire \tok.n23 ;
    wire \tok.n950 ;
    wire \tok.A__15__N_129 ;
    wire \tok.A_15_N_113_3 ;
    wire \tok.A_3 ;
    wire \tok.n4528_cascade_ ;
    wire \tok.n892_cascade_ ;
    wire \tok.n10_adj_818 ;
    wire \tok.n13_adj_842 ;
    wire \tok.n8_adj_666 ;
    wire \tok.n8_adj_777 ;
    wire \tok.n4502_cascade_ ;
    wire \tok.n12_adj_830 ;
    wire \tok.n4607 ;
    wire \tok.n9_adj_689 ;
    wire \tok.n181_cascade_ ;
    wire \tok.n12_cascade_ ;
    wire \tok.n6_adj_653 ;
    wire \tok.n20_cascade_ ;
    wire \tok.n16 ;
    wire \tok.n4684 ;
    wire \tok.n892 ;
    wire \tok.n177_cascade_ ;
    wire \tok.n12_adj_696_cascade_ ;
    wire \tok.n20_adj_700 ;
    wire \tok.n52 ;
    wire \tok.n33_adj_663 ;
    wire bfn_8_13_0_;
    wire \tok.n50 ;
    wire \tok.n33_adj_841 ;
    wire \tok.n3888 ;
    wire \tok.n49 ;
    wire \tok.n33_adj_665 ;
    wire \tok.n3889 ;
    wire \tok.n47 ;
    wire \tok.n33_adj_755 ;
    wire \tok.n3890 ;
    wire \tok.n45 ;
    wire \tok.n33_adj_852 ;
    wire \tok.n3891 ;
    wire \tok.n44 ;
    wire \tok.n3892 ;
    wire \tok.n3893 ;
    wire \tok.n39 ;
    wire \tok.n3894 ;
    wire \tok.n33_adj_643 ;
    wire \tok.C_stk.tail_20 ;
    wire \tok.tail_26 ;
    wire \tok.tail_12 ;
    wire \tok.C_stk.tail_36 ;
    wire \tok.tail_56 ;
    wire \tok.tail_40 ;
    wire \tok.tail_48 ;
    wire \tok.n83_adj_704 ;
    wire \tok.n4694_cascade_ ;
    wire \tok.n13_adj_713_cascade_ ;
    wire \tok.C_stk.n4894_cascade_ ;
    wire \tok.c_stk_r_0 ;
    wire \tok.ram.n4717_cascade_ ;
    wire \tok.n1_adj_712 ;
    wire \tok.C_stk.tail_7 ;
    wire \tok.C_stk.n4912_cascade_ ;
    wire \tok.tc_6 ;
    wire \tok.c_stk_r_7 ;
    wire \tok.ram.n4696_cascade_ ;
    wire \tok.n4602 ;
    wire \tok.n1_adj_798_cascade_ ;
    wire \tok.n13_adj_799 ;
    wire \tok.tc_0 ;
    wire \tok.tc_plus_1_0 ;
    wire bfn_9_5_0_;
    wire \tok.tc_plus_1_1 ;
    wire \tok.n3895 ;
    wire \tok.n3896 ;
    wire \tok.n3897 ;
    wire \tok.n3898 ;
    wire \tok.n3899 ;
    wire \tok.tc_plus_1_6 ;
    wire \tok.n3900 ;
    wire \tok.n3901 ;
    wire \tok.tc_plus_1_7 ;
    wire n92_adj_872;
    wire c_stk_w_7_N_18_7;
    wire n92_adj_871;
    wire c_stk_w_7_N_18_6;
    wire n92;
    wire c_stk_w_7_N_18_1;
    wire n10_adj_875;
    wire c_stk_w_7_N_18_0;
    wire \tok.found_slot ;
    wire \tok.n5_adj_655_cascade_ ;
    wire \tok.uart_tx_busy ;
    wire \tok.uart_rx_valid ;
    wire \tok.uart_stall_cascade_ ;
    wire \tok.n2732 ;
    wire \tok.n2732_cascade_ ;
    wire \tok.n43 ;
    wire \tok.n5_adj_655 ;
    wire \tok.reset_N_2 ;
    wire \tok.uart_stall ;
    wire \tok.n2724 ;
    wire \tok.n4431 ;
    wire \tok.n5_adj_682 ;
    wire bfn_9_8_0_;
    wire \tok.S_1 ;
    wire \tok.n4_adj_790 ;
    wire \tok.n3925 ;
    wire \tok.S_2 ;
    wire \tok.n5_adj_789 ;
    wire \tok.n3926 ;
    wire \tok.n3927 ;
    wire \tok.n3928 ;
    wire \tok.S_5 ;
    wire \tok.n5_adj_775 ;
    wire \tok.n3929 ;
    wire \tok.n5_adj_773 ;
    wire \tok.n3930 ;
    wire \tok.A_low_7 ;
    wire \tok.S_7 ;
    wire \tok.n5_adj_752 ;
    wire \tok.n3931 ;
    wire \tok.n3932 ;
    wire \tok.S_8 ;
    wire bfn_9_9_0_;
    wire \tok.S_9 ;
    wire \tok.n21 ;
    wire \tok.n3933 ;
    wire \tok.n58 ;
    wire \tok.S_10 ;
    wire \tok.n5_adj_668 ;
    wire \tok.n3934 ;
    wire \tok.S_11 ;
    wire \tok.n5_adj_690 ;
    wire \tok.n3935 ;
    wire \tok.S_12 ;
    wire \tok.n3936 ;
    wire \tok.n55 ;
    wire \tok.S_13 ;
    wire \tok.n3937 ;
    wire \tok.S_14 ;
    wire \tok.n5_adj_729 ;
    wire \tok.n3938 ;
    wire \tok.S_15 ;
    wire \tok.n53 ;
    wire \tok.n3939 ;
    wire \tok.n5_adj_750 ;
    wire \tok.n6_adj_812 ;
    wire \tok.n9_adj_836 ;
    wire \tok.n5_adj_837_cascade_ ;
    wire \tok.S_3 ;
    wire \tok.n23_adj_788 ;
    wire \tok.n10_adj_838_cascade_ ;
    wire \tok.n12_adj_840 ;
    wire \tok.n57 ;
    wire \tok.n6_adj_835 ;
    wire uart_rx_data_6;
    wire \tok.n109_cascade_ ;
    wire \tok.S_6 ;
    wire \tok.n18_adj_782 ;
    wire capture_4;
    wire uart_rx_data_3;
    wire bfn_9_11_0_;
    wire \tok.n13_adj_816 ;
    wire \tok.n3902 ;
    wire \tok.n2_adj_811 ;
    wire \tok.n3903 ;
    wire \tok.n26_adj_808 ;
    wire \tok.n3904 ;
    wire \tok.n3905 ;
    wire \tok.n3906 ;
    wire \tok.A_low_2 ;
    wire \tok.n210 ;
    wire \tok.n3907 ;
    wire \tok.A_low_3 ;
    wire \tok.n209 ;
    wire \tok.n3908 ;
    wire \tok.n3909 ;
    wire CONSTANT_ONE_NET;
    wire bfn_9_12_0_;
    wire \tok.n2598 ;
    wire \tok.n211 ;
    wire \tok.n2_adj_810 ;
    wire \tok.n5_adj_710 ;
    wire \tok.n6_adj_711 ;
    wire \tok.n4664 ;
    wire \tok.n4663 ;
    wire \tok.n33 ;
    wire \tok.n27 ;
    wire \tok.n296 ;
    wire \tok.n191 ;
    wire \tok.n59 ;
    wire \tok.n2_adj_703 ;
    wire \tok.stall ;
    wire \tok.A_low_5 ;
    wire \tok.search_clk ;
    wire \tok.n33_adj_817 ;
    wire \tok.n27_adj_868 ;
    wire \tok.n82 ;
    wire capture_5;
    wire rx_data_7__N_511;
    wire \tok.n9_adj_807 ;
    wire uart_rx_data_4;
    wire \tok.n3_adj_826 ;
    wire \tok.n6_adj_827_cascade_ ;
    wire \tok.n36 ;
    wire \tok.n33_adj_828_cascade_ ;
    wire \tok.n11_adj_831 ;
    wire \tok.n56 ;
    wire \tok.n2514 ;
    wire \tok.C_stk.tail_0 ;
    wire \tok.tail_8 ;
    wire \tok.tail_15 ;
    wire \tok.C_stk.tail_23 ;
    wire \tok.tail_31 ;
    wire \tok.C_stk.tail_39 ;
    wire \tok.tail_47 ;
    wire \tok.C_stk.tail_16 ;
    wire \tok.C_stk.tail_32 ;
    wire \tok.tail_24 ;
    wire \tok.tail_30 ;
    wire \tok.C_stk.tail_38 ;
    wire \tok.tail_46 ;
    wire \tok.c_stk_r_6 ;
    wire \tok.tail_44 ;
    wire \tok.C_stk.tail_18 ;
    wire \tok.n240 ;
    wire \tok.tail_55 ;
    wire \tok.tail_63 ;
    wire \tok.tail_54 ;
    wire \tok.tail_62 ;
    wire \tok.tail_52 ;
    wire \tok.tail_60 ;
    wire \tok.C_stk.n4900_cascade_ ;
    wire \tok.table_rd_5 ;
    wire \tok.n83_adj_742_cascade_ ;
    wire \tok.n4651_cascade_ ;
    wire \tok.ram.n4702_cascade_ ;
    wire \tok.n1_adj_757 ;
    wire \tok.tc_plus_1_5 ;
    wire \tok.n13_adj_758 ;
    wire n10_adj_873;
    wire n10_adj_873_cascade_;
    wire c_stk_w_7_N_18_5;
    wire \tok.tc_5 ;
    wire n10_adj_874;
    wire n10_adj_874_cascade_;
    wire \tok.tc_2 ;
    wire \tok.tc_plus_1_3 ;
    wire n92_adj_870;
    wire n92_adj_870_cascade_;
    wire c_stk_w_7_N_18_3;
    wire \tok.tc_3 ;
    wire stall_;
    wire \tok.tc_4 ;
    wire \tok.n9_adj_797 ;
    wire \tok.n11_adj_647 ;
    wire \tok.n4575_cascade_ ;
    wire \tok.n83_cascade_ ;
    wire \tok.n40 ;
    wire \tok.n4571_cascade_ ;
    wire \tok.n4393 ;
    wire \tok.n4460_cascade_ ;
    wire \tok.n2726 ;
    wire \tok.S_4 ;
    wire \tok.n13_adj_787 ;
    wire \tok.n10_adj_829_cascade_ ;
    wire \tok.n13_adj_833 ;
    wire \tok.n2746 ;
    wire \tok.n8_adj_839 ;
    wire \tok.table_rd_0 ;
    wire \tok.n18_adj_681 ;
    wire \tok.A_low_1 ;
    wire \tok.n101 ;
    wire \tok.n54 ;
    wire \tok.n244_cascade_ ;
    wire \tok.n17_adj_785 ;
    wire \tok.n60 ;
    wire \tok.n83 ;
    wire \tok.n3 ;
    wire \tok.n4478 ;
    wire \tok.c_stk_r_5 ;
    wire \tok.C_stk.tail_5 ;
    wire \tok.tail_13 ;
    wire \tok.C_stk.tail_21 ;
    wire \tok.tail_29 ;
    wire \tok.C_stk.tail_37 ;
    wire \tok.tail_61 ;
    wire \tok.tail_45 ;
    wire \tok.tail_53 ;
    wire \tok.C_stk.tail_22 ;
    wire \tok.C_stk.tail_6 ;
    wire \tok.tail_14 ;
    wire \tok.tail_11 ;
    wire \tok.C_stk.tail_19 ;
    wire \tok.tail_27 ;
    wire \tok.C_stk.tail_35 ;
    wire \tok.tail_59 ;
    wire \tok.tail_43 ;
    wire \tok.tail_51 ;
    wire \tok.tail_10 ;
    wire \tok.C_stk_delta_1 ;
    wire \tok.rd_7__N_374 ;
    wire c_stk_w_7_N_18_4;
    wire \tok.C_stk.tail_4 ;
    wire \tok.C_stk.n4888_cascade_ ;
    wire \tok.ram.n4705_cascade_ ;
    wire \tok.n1_adj_745_cascade_ ;
    wire \tok.tc_plus_1_4 ;
    wire \tok.n802 ;
    wire \tok.n13_adj_746_cascade_ ;
    wire \tok.n86 ;
    wire n10;
    wire \tok.C_stk.tail_3 ;
    wire \tok.C_stk.n4882 ;
    wire \tok.n602 ;
    wire c_stk_w_7_N_18_2;
    wire \tok.C_stk.tail_2 ;
    wire \tok.C_stk.n4876_cascade_ ;
    wire \tok.C_stk.n600 ;
    wire clk;
    wire \tok.tc_plus_1_2 ;
    wire \tok.tc__7__N_134 ;
    wire \tok.ram.n4711_cascade_ ;
    wire \tok.n1_adj_724_cascade_ ;
    wire \tok.n13_adj_725 ;
    wire \tok.n101_adj_776 ;
    wire \tok.ram.n4708 ;
    wire \tok.n1_adj_736 ;
    wire \tok.n5_adj_737 ;
    wire \tok.c_stk_r_2 ;
    wire \tok.table_rd_2 ;
    wire \tok.n83_adj_721_cascade_ ;
    wire \tok.n4692 ;
    wire \tok.ram.n14_adj_631_cascade_ ;
    wire \tok.n2635 ;
    wire \tok.n4_adj_795 ;
    wire \tok.n41_cascade_ ;
    wire \tok.n884 ;
    wire \tok.n14_adj_702 ;
    wire \tok.n15_adj_662 ;
    wire \tok.n4464 ;
    wire \tok.n4573 ;
    wire \tok.n9_adj_645 ;
    wire \tok.n11 ;
    wire \tok.n6_cascade_ ;
    wire \tok.n14 ;
    wire \tok.n4422_cascade_ ;
    wire \tok.n11_adj_648 ;
    wire \tok.n4558 ;
    wire \tok.n14_adj_650 ;
    wire \tok.n51_cascade_ ;
    wire \tok.n4424 ;
    wire \tok.n48 ;
    wire \tok.table_rd_12 ;
    wire \tok.n5_adj_694 ;
    wire \tok.n10_adj_697 ;
    wire \tok.n14_adj_695_cascade_ ;
    wire \tok.A_low_4 ;
    wire \tok.n18_adj_698 ;
    wire \tok.n2177 ;
    wire \tok.n14_adj_825 ;
    wire \tok.n2177_cascade_ ;
    wire \tok.n10_adj_646 ;
    wire \tok.n132 ;
    wire \tok.table_rd_8 ;
    wire \tok.n132_cascade_ ;
    wire \tok.n5 ;
    wire \tok.n10_adj_652 ;
    wire \tok.n14_adj_651 ;
    wire \tok.n109 ;
    wire \tok.A_low_0 ;
    wire \tok.n18 ;
    wire \tok.A_low_6 ;
    wire \tok.n179 ;
    wire \tok.n10_adj_675 ;
    wire \tok.n9 ;
    wire \tok.n10_adj_675_cascade_ ;
    wire \tok.n2586 ;
    wire \tok.T_3 ;
    wire \tok.n2178 ;
    wire \tok.n41 ;
    wire \tok.n4484 ;
    wire \tok.n40_adj_661 ;
    wire \tok.n42 ;
    wire \tok.n4688 ;
    wire \tok.n10 ;
    wire \tok.n14_adj_658_cascade_ ;
    wire \tok.n399 ;
    wire \tok.table_rd_4 ;
    wire \tok.c_stk_r_4 ;
    wire \tok.n83_adj_743 ;
    wire \tok.c_stk_r_3 ;
    wire \tok.T_1 ;
    wire \tok.table_rd_3 ;
    wire \tok.T_0 ;
    wire \tok.n83_adj_733_cascade_ ;
    wire \tok.T_2 ;
    wire \tok.n4627 ;
    wire \tok.n883 ;
    wire \tok.n10_adj_679 ;
    wire \tok.S_0 ;
    wire \tok.n2616 ;
    wire \tok.n15_adj_680 ;
    wire \tok.n14_adj_658 ;
    wire \tok.n11_adj_649 ;
    wire \tok.write_flag ;
    wire \tok.T_4 ;
    wire \tok.T_7 ;
    wire \tok.T_5 ;
    wire \tok.T_6 ;
    wire \tok.n8 ;
    wire _gnd_net_;

    defparam \tok.vals.mem1_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .WRITE_MODE=0;
    defparam \tok.vals.mem1_physical .READ_MODE=0;
    defparam \tok.vals.mem1_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.vals.mem1_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \tok.vals.mem1_physical  (
            .RDATA({\tok.table_rd_15 ,\tok.table_rd_14 ,\tok.table_rd_13 ,\tok.table_rd_12 ,\tok.table_rd_11 ,\tok.table_rd_10 ,\tok.table_rd_9 ,\tok.table_rd_8 ,\tok.table_rd_7 ,\tok.table_rd_6 ,\tok.table_rd_5 ,\tok.table_rd_4 ,\tok.table_rd_3 ,\tok.table_rd_2 ,\tok.table_rd_1 ,\tok.table_rd_0 }),
            .RADDR({dangling_wire_0,dangling_wire_1,dangling_wire_2,N__18058,N__19219,N__18127,N__18209,N__18286,N__18352,N__18427,N__17809}),
            .WADDR({dangling_wire_3,dangling_wire_4,dangling_wire_5,N__18055,N__19216,N__18124,N__18206,N__18283,N__18355,N__18424,N__17806}),
            .MASK({dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .WDATA({N__10730,N__10718,N__10703,N__11000,N__12050,N__14888,N__10643,N__10739,N__12014,N__17000,N__14822,N__12005,N__13238,N__16892,N__11993,N__17054}),
            .RCLKE(),
            .RCLK(N__26234),
            .RE(N__21681),
            .WCLKE(),
            .WCLK(N__26233),
            .WE(N__14846));
    defparam \tok.keys.mem0_physical .WRITE_MODE=0;
    defparam \tok.keys.mem0_physical .READ_MODE=0;
    defparam \tok.keys.mem0_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.keys.mem0_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \tok.keys.mem0_physical  (
            .RDATA({\tok.key_rd_15 ,\tok.key_rd_14 ,\tok.key_rd_13 ,\tok.key_rd_12 ,\tok.key_rd_11 ,\tok.key_rd_10 ,\tok.key_rd_9 ,\tok.key_rd_8 ,\tok.key_rd_7 ,\tok.key_rd_6 ,\tok.key_rd_5 ,\tok.key_rd_4 ,\tok.key_rd_3 ,\tok.key_rd_2 ,\tok.key_rd_1 ,\tok.key_rd_0 }),
            .RADDR({dangling_wire_22,dangling_wire_23,dangling_wire_24,N__18068,N__19229,N__18137,N__18221,N__18296,N__18364,N__18437,N__17819}),
            .WADDR({dangling_wire_25,dangling_wire_26,dangling_wire_27,N__18067,N__19228,N__18136,N__18220,N__18295,N__18365,N__18436,N__17818}),
            .MASK({dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .WDATA({N__20314,N__24004,N__20681,N__22995,N__21436,N__21067,N__22640,N__24839,N__19762,N__28269,N__22400,N__27447,N__21850,N__21988,N__24187,N__26941}),
            .RCLKE(),
            .RCLK(N__26221),
            .RE(N__21698),
            .WCLKE(),
            .WCLK(N__26222),
            .WE(N__14845));
    defparam \tok.ram.mem2_physical .INIT_0=256'b0000000000000000000001000000010000000101010000000000010100000100000001000000000000000100000001000000010100010101000001010000010000000100000000000000010000000100000001010001010000000101000001000000010000000000000001000000010000000101000100010000010100000100;
    defparam \tok.ram.mem2_physical .WRITE_MODE=1;
    defparam \tok.ram.mem2_physical .READ_MODE=1;
    defparam \tok.ram.mem2_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \tok.ram.mem2_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \tok.ram.mem2_physical  (
            .RDATA({dangling_wire_44,\tok.T_7 ,dangling_wire_45,\tok.T_6 ,dangling_wire_46,\tok.T_5 ,dangling_wire_47,\tok.T_4 ,dangling_wire_48,\tok.T_3 ,dangling_wire_49,\tok.T_2 ,dangling_wire_50,\tok.T_1 ,dangling_wire_51,\tok.T_0 }),
            .RADDR({dangling_wire_52,dangling_wire_53,dangling_wire_54,N__16844,N__18548,N__23663,N__23447,N__23534,N__23639,N__16745,N__18692}),
            .WADDR({dangling_wire_55,dangling_wire_56,dangling_wire_57,N__19690,N__21322,N__19952,N__24395,N__21551,N__20068,N__20171,N__29575}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,N__19824,dangling_wire_75,N__28268,dangling_wire_76,N__22401,dangling_wire_77,N__27452,dangling_wire_78,N__21845,dangling_wire_79,N__21985,dangling_wire_80,N__24181,dangling_wire_81,N__26934}),
            .RCLKE(),
            .RCLK(N__26258),
            .RE(N__21699),
            .WCLKE(),
            .WCLK(N__26259),
            .WE(N__29101));
    defparam rx_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_pad_iopad.PULLUP=1'b0;
    IO_PAD rx_pad_iopad (
            .OE(N__30609),
            .DIN(N__30608),
            .DOUT(N__30607),
            .PACKAGEPIN(rx));
    defparam rx_pad_preio.PIN_TYPE=6'b000001;
    defparam rx_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_pad_preio (
            .PADOEN(N__30609),
            .PADOUT(N__30608),
            .PADIN(N__30607),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(rx_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam tx_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_pad_iopad.PULLUP=1'b0;
    IO_PAD tx_pad_iopad (
            .OE(N__30600),
            .DIN(N__30599),
            .DOUT(N__30598),
            .PACKAGEPIN(tx));
    defparam tx_pad_preio.PIN_TYPE=6'b011001;
    defparam tx_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_pad_preio (
            .PADOEN(N__30600),
            .PADOUT(N__30599),
            .PADIN(N__30598),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13289),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam reset_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam reset_pad_iopad.PULLUP=1'b0;
    IO_PAD reset_pad_iopad (
            .OE(N__30591),
            .DIN(N__30590),
            .DOUT(N__30589),
            .PACKAGEPIN(reset));
    defparam reset_pad_preio.PIN_TYPE=6'b000001;
    defparam reset_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO reset_pad_preio (
            .PADOEN(N__30591),
            .PADOUT(N__30590),
            .PADIN(N__30589),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(reset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__7643 (
            .O(N__30572),
            .I(N__30568));
    InMux I__7642 (
            .O(N__30571),
            .I(N__30565));
    LocalMux I__7641 (
            .O(N__30568),
            .I(N__30562));
    LocalMux I__7640 (
            .O(N__30565),
            .I(N__30559));
    Span4Mux_v I__7639 (
            .O(N__30562),
            .I(N__30556));
    Span4Mux_v I__7638 (
            .O(N__30559),
            .I(N__30553));
    Span4Mux_h I__7637 (
            .O(N__30556),
            .I(N__30550));
    Sp12to4 I__7636 (
            .O(N__30553),
            .I(N__30545));
    Sp12to4 I__7635 (
            .O(N__30550),
            .I(N__30545));
    Span12Mux_s10_h I__7634 (
            .O(N__30545),
            .I(N__30542));
    Odrv12 I__7633 (
            .O(N__30542),
            .I(\tok.table_rd_4 ));
    CascadeMux I__7632 (
            .O(N__30539),
            .I(N__30532));
    InMux I__7631 (
            .O(N__30538),
            .I(N__30529));
    InMux I__7630 (
            .O(N__30537),
            .I(N__30526));
    InMux I__7629 (
            .O(N__30536),
            .I(N__30519));
    InMux I__7628 (
            .O(N__30535),
            .I(N__30519));
    InMux I__7627 (
            .O(N__30532),
            .I(N__30519));
    LocalMux I__7626 (
            .O(N__30529),
            .I(N__30516));
    LocalMux I__7625 (
            .O(N__30526),
            .I(N__30513));
    LocalMux I__7624 (
            .O(N__30519),
            .I(N__30510));
    Span4Mux_h I__7623 (
            .O(N__30516),
            .I(N__30505));
    Span4Mux_v I__7622 (
            .O(N__30513),
            .I(N__30505));
    Odrv4 I__7621 (
            .O(N__30510),
            .I(\tok.c_stk_r_4 ));
    Odrv4 I__7620 (
            .O(N__30505),
            .I(\tok.c_stk_r_4 ));
    InMux I__7619 (
            .O(N__30500),
            .I(N__30497));
    LocalMux I__7618 (
            .O(N__30497),
            .I(\tok.n83_adj_743 ));
    InMux I__7617 (
            .O(N__30494),
            .I(N__30490));
    CascadeMux I__7616 (
            .O(N__30493),
            .I(N__30484));
    LocalMux I__7615 (
            .O(N__30490),
            .I(N__30481));
    CascadeMux I__7614 (
            .O(N__30489),
            .I(N__30478));
    InMux I__7613 (
            .O(N__30488),
            .I(N__30475));
    InMux I__7612 (
            .O(N__30487),
            .I(N__30472));
    InMux I__7611 (
            .O(N__30484),
            .I(N__30469));
    Span4Mux_v I__7610 (
            .O(N__30481),
            .I(N__30466));
    InMux I__7609 (
            .O(N__30478),
            .I(N__30463));
    LocalMux I__7608 (
            .O(N__30475),
            .I(\tok.c_stk_r_3 ));
    LocalMux I__7607 (
            .O(N__30472),
            .I(\tok.c_stk_r_3 ));
    LocalMux I__7606 (
            .O(N__30469),
            .I(\tok.c_stk_r_3 ));
    Odrv4 I__7605 (
            .O(N__30466),
            .I(\tok.c_stk_r_3 ));
    LocalMux I__7604 (
            .O(N__30463),
            .I(\tok.c_stk_r_3 ));
    CascadeMux I__7603 (
            .O(N__30452),
            .I(N__30449));
    InMux I__7602 (
            .O(N__30449),
            .I(N__30438));
    InMux I__7601 (
            .O(N__30448),
            .I(N__30433));
    InMux I__7600 (
            .O(N__30447),
            .I(N__30433));
    InMux I__7599 (
            .O(N__30446),
            .I(N__30424));
    InMux I__7598 (
            .O(N__30445),
            .I(N__30424));
    InMux I__7597 (
            .O(N__30444),
            .I(N__30424));
    InMux I__7596 (
            .O(N__30443),
            .I(N__30424));
    CascadeMux I__7595 (
            .O(N__30442),
            .I(N__30420));
    InMux I__7594 (
            .O(N__30441),
            .I(N__30413));
    LocalMux I__7593 (
            .O(N__30438),
            .I(N__30405));
    LocalMux I__7592 (
            .O(N__30433),
            .I(N__30405));
    LocalMux I__7591 (
            .O(N__30424),
            .I(N__30402));
    InMux I__7590 (
            .O(N__30423),
            .I(N__30395));
    InMux I__7589 (
            .O(N__30420),
            .I(N__30395));
    InMux I__7588 (
            .O(N__30419),
            .I(N__30395));
    CascadeMux I__7587 (
            .O(N__30418),
            .I(N__30386));
    InMux I__7586 (
            .O(N__30417),
            .I(N__30375));
    InMux I__7585 (
            .O(N__30416),
            .I(N__30375));
    LocalMux I__7584 (
            .O(N__30413),
            .I(N__30372));
    InMux I__7583 (
            .O(N__30412),
            .I(N__30369));
    InMux I__7582 (
            .O(N__30411),
            .I(N__30366));
    InMux I__7581 (
            .O(N__30410),
            .I(N__30363));
    Span4Mux_h I__7580 (
            .O(N__30405),
            .I(N__30356));
    Span4Mux_s3_v I__7579 (
            .O(N__30402),
            .I(N__30356));
    LocalMux I__7578 (
            .O(N__30395),
            .I(N__30356));
    InMux I__7577 (
            .O(N__30394),
            .I(N__30353));
    InMux I__7576 (
            .O(N__30393),
            .I(N__30349));
    InMux I__7575 (
            .O(N__30392),
            .I(N__30346));
    InMux I__7574 (
            .O(N__30391),
            .I(N__30340));
    InMux I__7573 (
            .O(N__30390),
            .I(N__30340));
    InMux I__7572 (
            .O(N__30389),
            .I(N__30333));
    InMux I__7571 (
            .O(N__30386),
            .I(N__30333));
    InMux I__7570 (
            .O(N__30385),
            .I(N__30333));
    InMux I__7569 (
            .O(N__30384),
            .I(N__30324));
    InMux I__7568 (
            .O(N__30383),
            .I(N__30324));
    InMux I__7567 (
            .O(N__30382),
            .I(N__30324));
    InMux I__7566 (
            .O(N__30381),
            .I(N__30324));
    InMux I__7565 (
            .O(N__30380),
            .I(N__30319));
    LocalMux I__7564 (
            .O(N__30375),
            .I(N__30316));
    Span4Mux_v I__7563 (
            .O(N__30372),
            .I(N__30313));
    LocalMux I__7562 (
            .O(N__30369),
            .I(N__30310));
    LocalMux I__7561 (
            .O(N__30366),
            .I(N__30301));
    LocalMux I__7560 (
            .O(N__30363),
            .I(N__30301));
    Span4Mux_h I__7559 (
            .O(N__30356),
            .I(N__30301));
    LocalMux I__7558 (
            .O(N__30353),
            .I(N__30301));
    InMux I__7557 (
            .O(N__30352),
            .I(N__30298));
    LocalMux I__7556 (
            .O(N__30349),
            .I(N__30295));
    LocalMux I__7555 (
            .O(N__30346),
            .I(N__30292));
    CascadeMux I__7554 (
            .O(N__30345),
            .I(N__30283));
    LocalMux I__7553 (
            .O(N__30340),
            .I(N__30276));
    LocalMux I__7552 (
            .O(N__30333),
            .I(N__30271));
    LocalMux I__7551 (
            .O(N__30324),
            .I(N__30271));
    InMux I__7550 (
            .O(N__30323),
            .I(N__30266));
    InMux I__7549 (
            .O(N__30322),
            .I(N__30266));
    LocalMux I__7548 (
            .O(N__30319),
            .I(N__30263));
    Span4Mux_v I__7547 (
            .O(N__30316),
            .I(N__30260));
    Span4Mux_h I__7546 (
            .O(N__30313),
            .I(N__30253));
    Span4Mux_v I__7545 (
            .O(N__30310),
            .I(N__30253));
    Span4Mux_v I__7544 (
            .O(N__30301),
            .I(N__30253));
    LocalMux I__7543 (
            .O(N__30298),
            .I(N__30250));
    Span4Mux_v I__7542 (
            .O(N__30295),
            .I(N__30245));
    Span4Mux_s2_h I__7541 (
            .O(N__30292),
            .I(N__30245));
    InMux I__7540 (
            .O(N__30291),
            .I(N__30238));
    InMux I__7539 (
            .O(N__30290),
            .I(N__30238));
    InMux I__7538 (
            .O(N__30289),
            .I(N__30238));
    InMux I__7537 (
            .O(N__30288),
            .I(N__30231));
    InMux I__7536 (
            .O(N__30287),
            .I(N__30231));
    InMux I__7535 (
            .O(N__30286),
            .I(N__30231));
    InMux I__7534 (
            .O(N__30283),
            .I(N__30220));
    InMux I__7533 (
            .O(N__30282),
            .I(N__30220));
    InMux I__7532 (
            .O(N__30281),
            .I(N__30220));
    InMux I__7531 (
            .O(N__30280),
            .I(N__30220));
    InMux I__7530 (
            .O(N__30279),
            .I(N__30220));
    Span4Mux_h I__7529 (
            .O(N__30276),
            .I(N__30213));
    Span4Mux_s3_h I__7528 (
            .O(N__30271),
            .I(N__30213));
    LocalMux I__7527 (
            .O(N__30266),
            .I(N__30213));
    Odrv4 I__7526 (
            .O(N__30263),
            .I(\tok.T_1 ));
    Odrv4 I__7525 (
            .O(N__30260),
            .I(\tok.T_1 ));
    Odrv4 I__7524 (
            .O(N__30253),
            .I(\tok.T_1 ));
    Odrv4 I__7523 (
            .O(N__30250),
            .I(\tok.T_1 ));
    Odrv4 I__7522 (
            .O(N__30245),
            .I(\tok.T_1 ));
    LocalMux I__7521 (
            .O(N__30238),
            .I(\tok.T_1 ));
    LocalMux I__7520 (
            .O(N__30231),
            .I(\tok.T_1 ));
    LocalMux I__7519 (
            .O(N__30220),
            .I(\tok.T_1 ));
    Odrv4 I__7518 (
            .O(N__30213),
            .I(\tok.T_1 ));
    CascadeMux I__7517 (
            .O(N__30194),
            .I(N__30191));
    InMux I__7516 (
            .O(N__30191),
            .I(N__30188));
    LocalMux I__7515 (
            .O(N__30188),
            .I(N__30185));
    Span4Mux_v I__7514 (
            .O(N__30185),
            .I(N__30181));
    InMux I__7513 (
            .O(N__30184),
            .I(N__30178));
    Span4Mux_h I__7512 (
            .O(N__30181),
            .I(N__30175));
    LocalMux I__7511 (
            .O(N__30178),
            .I(N__30172));
    Span4Mux_h I__7510 (
            .O(N__30175),
            .I(N__30169));
    Odrv12 I__7509 (
            .O(N__30172),
            .I(\tok.table_rd_3 ));
    Odrv4 I__7508 (
            .O(N__30169),
            .I(\tok.table_rd_3 ));
    InMux I__7507 (
            .O(N__30164),
            .I(N__30138));
    InMux I__7506 (
            .O(N__30163),
            .I(N__30138));
    InMux I__7505 (
            .O(N__30162),
            .I(N__30138));
    InMux I__7504 (
            .O(N__30161),
            .I(N__30131));
    InMux I__7503 (
            .O(N__30160),
            .I(N__30128));
    InMux I__7502 (
            .O(N__30159),
            .I(N__30121));
    InMux I__7501 (
            .O(N__30158),
            .I(N__30121));
    InMux I__7500 (
            .O(N__30157),
            .I(N__30121));
    InMux I__7499 (
            .O(N__30156),
            .I(N__30114));
    InMux I__7498 (
            .O(N__30155),
            .I(N__30114));
    InMux I__7497 (
            .O(N__30154),
            .I(N__30114));
    InMux I__7496 (
            .O(N__30153),
            .I(N__30099));
    InMux I__7495 (
            .O(N__30152),
            .I(N__30094));
    InMux I__7494 (
            .O(N__30151),
            .I(N__30094));
    InMux I__7493 (
            .O(N__30150),
            .I(N__30089));
    InMux I__7492 (
            .O(N__30149),
            .I(N__30089));
    InMux I__7491 (
            .O(N__30148),
            .I(N__30086));
    InMux I__7490 (
            .O(N__30147),
            .I(N__30083));
    InMux I__7489 (
            .O(N__30146),
            .I(N__30078));
    InMux I__7488 (
            .O(N__30145),
            .I(N__30078));
    LocalMux I__7487 (
            .O(N__30138),
            .I(N__30075));
    InMux I__7486 (
            .O(N__30137),
            .I(N__30072));
    InMux I__7485 (
            .O(N__30136),
            .I(N__30069));
    InMux I__7484 (
            .O(N__30135),
            .I(N__30066));
    InMux I__7483 (
            .O(N__30134),
            .I(N__30063));
    LocalMux I__7482 (
            .O(N__30131),
            .I(N__30056));
    LocalMux I__7481 (
            .O(N__30128),
            .I(N__30056));
    LocalMux I__7480 (
            .O(N__30121),
            .I(N__30056));
    LocalMux I__7479 (
            .O(N__30114),
            .I(N__30053));
    InMux I__7478 (
            .O(N__30113),
            .I(N__30050));
    InMux I__7477 (
            .O(N__30112),
            .I(N__30045));
    InMux I__7476 (
            .O(N__30111),
            .I(N__30045));
    InMux I__7475 (
            .O(N__30110),
            .I(N__30041));
    InMux I__7474 (
            .O(N__30109),
            .I(N__30037));
    InMux I__7473 (
            .O(N__30108),
            .I(N__30030));
    InMux I__7472 (
            .O(N__30107),
            .I(N__30030));
    InMux I__7471 (
            .O(N__30106),
            .I(N__30030));
    InMux I__7470 (
            .O(N__30105),
            .I(N__30021));
    InMux I__7469 (
            .O(N__30104),
            .I(N__30021));
    InMux I__7468 (
            .O(N__30103),
            .I(N__30021));
    InMux I__7467 (
            .O(N__30102),
            .I(N__30021));
    LocalMux I__7466 (
            .O(N__30099),
            .I(N__30015));
    LocalMux I__7465 (
            .O(N__30094),
            .I(N__30015));
    LocalMux I__7464 (
            .O(N__30089),
            .I(N__30010));
    LocalMux I__7463 (
            .O(N__30086),
            .I(N__30010));
    LocalMux I__7462 (
            .O(N__30083),
            .I(N__30001));
    LocalMux I__7461 (
            .O(N__30078),
            .I(N__30001));
    Span4Mux_v I__7460 (
            .O(N__30075),
            .I(N__30001));
    LocalMux I__7459 (
            .O(N__30072),
            .I(N__30001));
    LocalMux I__7458 (
            .O(N__30069),
            .I(N__29998));
    LocalMux I__7457 (
            .O(N__30066),
            .I(N__29995));
    LocalMux I__7456 (
            .O(N__30063),
            .I(N__29988));
    Span4Mux_s3_v I__7455 (
            .O(N__30056),
            .I(N__29988));
    Span4Mux_h I__7454 (
            .O(N__30053),
            .I(N__29988));
    LocalMux I__7453 (
            .O(N__30050),
            .I(N__29985));
    LocalMux I__7452 (
            .O(N__30045),
            .I(N__29982));
    InMux I__7451 (
            .O(N__30044),
            .I(N__29979));
    LocalMux I__7450 (
            .O(N__30041),
            .I(N__29976));
    CascadeMux I__7449 (
            .O(N__30040),
            .I(N__29970));
    LocalMux I__7448 (
            .O(N__30037),
            .I(N__29959));
    LocalMux I__7447 (
            .O(N__30030),
            .I(N__29954));
    LocalMux I__7446 (
            .O(N__30021),
            .I(N__29954));
    InMux I__7445 (
            .O(N__30020),
            .I(N__29951));
    Span4Mux_s3_h I__7444 (
            .O(N__30015),
            .I(N__29944));
    Span4Mux_h I__7443 (
            .O(N__30010),
            .I(N__29944));
    Span4Mux_h I__7442 (
            .O(N__30001),
            .I(N__29944));
    Span4Mux_v I__7441 (
            .O(N__29998),
            .I(N__29931));
    Span4Mux_h I__7440 (
            .O(N__29995),
            .I(N__29931));
    Span4Mux_v I__7439 (
            .O(N__29988),
            .I(N__29931));
    Span4Mux_v I__7438 (
            .O(N__29985),
            .I(N__29931));
    Span4Mux_v I__7437 (
            .O(N__29982),
            .I(N__29931));
    LocalMux I__7436 (
            .O(N__29979),
            .I(N__29931));
    Span4Mux_s2_h I__7435 (
            .O(N__29976),
            .I(N__29928));
    InMux I__7434 (
            .O(N__29975),
            .I(N__29921));
    InMux I__7433 (
            .O(N__29974),
            .I(N__29921));
    InMux I__7432 (
            .O(N__29973),
            .I(N__29921));
    InMux I__7431 (
            .O(N__29970),
            .I(N__29914));
    InMux I__7430 (
            .O(N__29969),
            .I(N__29914));
    InMux I__7429 (
            .O(N__29968),
            .I(N__29914));
    InMux I__7428 (
            .O(N__29967),
            .I(N__29911));
    InMux I__7427 (
            .O(N__29966),
            .I(N__29900));
    InMux I__7426 (
            .O(N__29965),
            .I(N__29900));
    InMux I__7425 (
            .O(N__29964),
            .I(N__29900));
    InMux I__7424 (
            .O(N__29963),
            .I(N__29900));
    InMux I__7423 (
            .O(N__29962),
            .I(N__29900));
    Span4Mux_s3_h I__7422 (
            .O(N__29959),
            .I(N__29893));
    Span4Mux_s3_h I__7421 (
            .O(N__29954),
            .I(N__29893));
    LocalMux I__7420 (
            .O(N__29951),
            .I(N__29893));
    Odrv4 I__7419 (
            .O(N__29944),
            .I(\tok.T_0 ));
    Odrv4 I__7418 (
            .O(N__29931),
            .I(\tok.T_0 ));
    Odrv4 I__7417 (
            .O(N__29928),
            .I(\tok.T_0 ));
    LocalMux I__7416 (
            .O(N__29921),
            .I(\tok.T_0 ));
    LocalMux I__7415 (
            .O(N__29914),
            .I(\tok.T_0 ));
    LocalMux I__7414 (
            .O(N__29911),
            .I(\tok.T_0 ));
    LocalMux I__7413 (
            .O(N__29900),
            .I(\tok.T_0 ));
    Odrv4 I__7412 (
            .O(N__29893),
            .I(\tok.T_0 ));
    CascadeMux I__7411 (
            .O(N__29876),
            .I(\tok.n83_adj_733_cascade_ ));
    InMux I__7410 (
            .O(N__29873),
            .I(N__29844));
    InMux I__7409 (
            .O(N__29872),
            .I(N__29837));
    InMux I__7408 (
            .O(N__29871),
            .I(N__29837));
    InMux I__7407 (
            .O(N__29870),
            .I(N__29837));
    InMux I__7406 (
            .O(N__29869),
            .I(N__29832));
    InMux I__7405 (
            .O(N__29868),
            .I(N__29832));
    InMux I__7404 (
            .O(N__29867),
            .I(N__29825));
    InMux I__7403 (
            .O(N__29866),
            .I(N__29825));
    InMux I__7402 (
            .O(N__29865),
            .I(N__29825));
    CascadeMux I__7401 (
            .O(N__29864),
            .I(N__29821));
    InMux I__7400 (
            .O(N__29863),
            .I(N__29814));
    InMux I__7399 (
            .O(N__29862),
            .I(N__29814));
    InMux I__7398 (
            .O(N__29861),
            .I(N__29811));
    InMux I__7397 (
            .O(N__29860),
            .I(N__29808));
    InMux I__7396 (
            .O(N__29859),
            .I(N__29803));
    InMux I__7395 (
            .O(N__29858),
            .I(N__29803));
    InMux I__7394 (
            .O(N__29857),
            .I(N__29794));
    InMux I__7393 (
            .O(N__29856),
            .I(N__29794));
    InMux I__7392 (
            .O(N__29855),
            .I(N__29791));
    InMux I__7391 (
            .O(N__29854),
            .I(N__29786));
    InMux I__7390 (
            .O(N__29853),
            .I(N__29786));
    InMux I__7389 (
            .O(N__29852),
            .I(N__29783));
    InMux I__7388 (
            .O(N__29851),
            .I(N__29779));
    InMux I__7387 (
            .O(N__29850),
            .I(N__29774));
    InMux I__7386 (
            .O(N__29849),
            .I(N__29774));
    InMux I__7385 (
            .O(N__29848),
            .I(N__29771));
    InMux I__7384 (
            .O(N__29847),
            .I(N__29768));
    LocalMux I__7383 (
            .O(N__29844),
            .I(N__29765));
    LocalMux I__7382 (
            .O(N__29837),
            .I(N__29762));
    LocalMux I__7381 (
            .O(N__29832),
            .I(N__29757));
    LocalMux I__7380 (
            .O(N__29825),
            .I(N__29757));
    InMux I__7379 (
            .O(N__29824),
            .I(N__29754));
    InMux I__7378 (
            .O(N__29821),
            .I(N__29747));
    InMux I__7377 (
            .O(N__29820),
            .I(N__29747));
    InMux I__7376 (
            .O(N__29819),
            .I(N__29747));
    LocalMux I__7375 (
            .O(N__29814),
            .I(N__29738));
    LocalMux I__7374 (
            .O(N__29811),
            .I(N__29738));
    LocalMux I__7373 (
            .O(N__29808),
            .I(N__29738));
    LocalMux I__7372 (
            .O(N__29803),
            .I(N__29738));
    InMux I__7371 (
            .O(N__29802),
            .I(N__29733));
    InMux I__7370 (
            .O(N__29801),
            .I(N__29733));
    InMux I__7369 (
            .O(N__29800),
            .I(N__29728));
    InMux I__7368 (
            .O(N__29799),
            .I(N__29728));
    LocalMux I__7367 (
            .O(N__29794),
            .I(N__29725));
    LocalMux I__7366 (
            .O(N__29791),
            .I(N__29718));
    LocalMux I__7365 (
            .O(N__29786),
            .I(N__29718));
    LocalMux I__7364 (
            .O(N__29783),
            .I(N__29718));
    InMux I__7363 (
            .O(N__29782),
            .I(N__29715));
    LocalMux I__7362 (
            .O(N__29779),
            .I(N__29712));
    LocalMux I__7361 (
            .O(N__29774),
            .I(N__29709));
    LocalMux I__7360 (
            .O(N__29771),
            .I(N__29706));
    LocalMux I__7359 (
            .O(N__29768),
            .I(N__29697));
    Span4Mux_h I__7358 (
            .O(N__29765),
            .I(N__29697));
    Span4Mux_s3_v I__7357 (
            .O(N__29762),
            .I(N__29697));
    Span4Mux_h I__7356 (
            .O(N__29757),
            .I(N__29697));
    LocalMux I__7355 (
            .O(N__29754),
            .I(N__29692));
    LocalMux I__7354 (
            .O(N__29747),
            .I(N__29692));
    Span4Mux_v I__7353 (
            .O(N__29738),
            .I(N__29689));
    LocalMux I__7352 (
            .O(N__29733),
            .I(N__29686));
    LocalMux I__7351 (
            .O(N__29728),
            .I(N__29671));
    Span4Mux_v I__7350 (
            .O(N__29725),
            .I(N__29666));
    Span4Mux_h I__7349 (
            .O(N__29718),
            .I(N__29666));
    LocalMux I__7348 (
            .O(N__29715),
            .I(N__29663));
    Span4Mux_v I__7347 (
            .O(N__29712),
            .I(N__29648));
    Span4Mux_h I__7346 (
            .O(N__29709),
            .I(N__29648));
    Span4Mux_h I__7345 (
            .O(N__29706),
            .I(N__29648));
    Span4Mux_v I__7344 (
            .O(N__29697),
            .I(N__29648));
    Span4Mux_v I__7343 (
            .O(N__29692),
            .I(N__29648));
    Span4Mux_s0_h I__7342 (
            .O(N__29689),
            .I(N__29648));
    Span4Mux_v I__7341 (
            .O(N__29686),
            .I(N__29648));
    InMux I__7340 (
            .O(N__29685),
            .I(N__29643));
    InMux I__7339 (
            .O(N__29684),
            .I(N__29643));
    InMux I__7338 (
            .O(N__29683),
            .I(N__29636));
    InMux I__7337 (
            .O(N__29682),
            .I(N__29636));
    InMux I__7336 (
            .O(N__29681),
            .I(N__29636));
    InMux I__7335 (
            .O(N__29680),
            .I(N__29621));
    InMux I__7334 (
            .O(N__29679),
            .I(N__29621));
    InMux I__7333 (
            .O(N__29678),
            .I(N__29621));
    InMux I__7332 (
            .O(N__29677),
            .I(N__29621));
    InMux I__7331 (
            .O(N__29676),
            .I(N__29621));
    InMux I__7330 (
            .O(N__29675),
            .I(N__29621));
    InMux I__7329 (
            .O(N__29674),
            .I(N__29621));
    Odrv4 I__7328 (
            .O(N__29671),
            .I(\tok.T_2 ));
    Odrv4 I__7327 (
            .O(N__29666),
            .I(\tok.T_2 ));
    Odrv4 I__7326 (
            .O(N__29663),
            .I(\tok.T_2 ));
    Odrv4 I__7325 (
            .O(N__29648),
            .I(\tok.T_2 ));
    LocalMux I__7324 (
            .O(N__29643),
            .I(\tok.T_2 ));
    LocalMux I__7323 (
            .O(N__29636),
            .I(\tok.T_2 ));
    LocalMux I__7322 (
            .O(N__29621),
            .I(\tok.T_2 ));
    CascadeMux I__7321 (
            .O(N__29606),
            .I(N__29603));
    InMux I__7320 (
            .O(N__29603),
            .I(N__29600));
    LocalMux I__7319 (
            .O(N__29600),
            .I(\tok.n4627 ));
    InMux I__7318 (
            .O(N__29597),
            .I(N__29594));
    LocalMux I__7317 (
            .O(N__29594),
            .I(\tok.n883 ));
    InMux I__7316 (
            .O(N__29591),
            .I(N__29588));
    LocalMux I__7315 (
            .O(N__29588),
            .I(N__29585));
    Sp12to4 I__7314 (
            .O(N__29585),
            .I(N__29582));
    Span12Mux_s7_v I__7313 (
            .O(N__29582),
            .I(N__29579));
    Odrv12 I__7312 (
            .O(N__29579),
            .I(\tok.n10_adj_679 ));
    CascadeMux I__7311 (
            .O(N__29576),
            .I(N__29568));
    CascadeMux I__7310 (
            .O(N__29575),
            .I(N__29565));
    CascadeMux I__7309 (
            .O(N__29574),
            .I(N__29562));
    InMux I__7308 (
            .O(N__29573),
            .I(N__29559));
    InMux I__7307 (
            .O(N__29572),
            .I(N__29556));
    CascadeMux I__7306 (
            .O(N__29571),
            .I(N__29553));
    InMux I__7305 (
            .O(N__29568),
            .I(N__29550));
    InMux I__7304 (
            .O(N__29565),
            .I(N__29545));
    InMux I__7303 (
            .O(N__29562),
            .I(N__29542));
    LocalMux I__7302 (
            .O(N__29559),
            .I(N__29539));
    LocalMux I__7301 (
            .O(N__29556),
            .I(N__29536));
    InMux I__7300 (
            .O(N__29553),
            .I(N__29533));
    LocalMux I__7299 (
            .O(N__29550),
            .I(N__29530));
    InMux I__7298 (
            .O(N__29549),
            .I(N__29527));
    InMux I__7297 (
            .O(N__29548),
            .I(N__29524));
    LocalMux I__7296 (
            .O(N__29545),
            .I(N__29519));
    LocalMux I__7295 (
            .O(N__29542),
            .I(N__29519));
    Span4Mux_v I__7294 (
            .O(N__29539),
            .I(N__29515));
    Span4Mux_v I__7293 (
            .O(N__29536),
            .I(N__29512));
    LocalMux I__7292 (
            .O(N__29533),
            .I(N__29509));
    Span4Mux_h I__7291 (
            .O(N__29530),
            .I(N__29506));
    LocalMux I__7290 (
            .O(N__29527),
            .I(N__29501));
    LocalMux I__7289 (
            .O(N__29524),
            .I(N__29501));
    Span4Mux_v I__7288 (
            .O(N__29519),
            .I(N__29498));
    InMux I__7287 (
            .O(N__29518),
            .I(N__29495));
    Span4Mux_h I__7286 (
            .O(N__29515),
            .I(N__29492));
    Span4Mux_h I__7285 (
            .O(N__29512),
            .I(N__29487));
    Span4Mux_v I__7284 (
            .O(N__29509),
            .I(N__29487));
    Span4Mux_v I__7283 (
            .O(N__29506),
            .I(N__29480));
    Span4Mux_v I__7282 (
            .O(N__29501),
            .I(N__29480));
    Span4Mux_h I__7281 (
            .O(N__29498),
            .I(N__29480));
    LocalMux I__7280 (
            .O(N__29495),
            .I(N__29473));
    Span4Mux_h I__7279 (
            .O(N__29492),
            .I(N__29473));
    Span4Mux_v I__7278 (
            .O(N__29487),
            .I(N__29473));
    Span4Mux_h I__7277 (
            .O(N__29480),
            .I(N__29470));
    Odrv4 I__7276 (
            .O(N__29473),
            .I(\tok.S_0 ));
    Odrv4 I__7275 (
            .O(N__29470),
            .I(\tok.S_0 ));
    InMux I__7274 (
            .O(N__29465),
            .I(N__29462));
    LocalMux I__7273 (
            .O(N__29462),
            .I(N__29454));
    InMux I__7272 (
            .O(N__29461),
            .I(N__29451));
    InMux I__7271 (
            .O(N__29460),
            .I(N__29446));
    InMux I__7270 (
            .O(N__29459),
            .I(N__29446));
    InMux I__7269 (
            .O(N__29458),
            .I(N__29441));
    InMux I__7268 (
            .O(N__29457),
            .I(N__29437));
    Span4Mux_h I__7267 (
            .O(N__29454),
            .I(N__29431));
    LocalMux I__7266 (
            .O(N__29451),
            .I(N__29431));
    LocalMux I__7265 (
            .O(N__29446),
            .I(N__29428));
    InMux I__7264 (
            .O(N__29445),
            .I(N__29425));
    InMux I__7263 (
            .O(N__29444),
            .I(N__29422));
    LocalMux I__7262 (
            .O(N__29441),
            .I(N__29418));
    InMux I__7261 (
            .O(N__29440),
            .I(N__29415));
    LocalMux I__7260 (
            .O(N__29437),
            .I(N__29412));
    InMux I__7259 (
            .O(N__29436),
            .I(N__29408));
    Span4Mux_v I__7258 (
            .O(N__29431),
            .I(N__29405));
    Span4Mux_h I__7257 (
            .O(N__29428),
            .I(N__29398));
    LocalMux I__7256 (
            .O(N__29425),
            .I(N__29398));
    LocalMux I__7255 (
            .O(N__29422),
            .I(N__29398));
    InMux I__7254 (
            .O(N__29421),
            .I(N__29395));
    Span4Mux_h I__7253 (
            .O(N__29418),
            .I(N__29387));
    LocalMux I__7252 (
            .O(N__29415),
            .I(N__29387));
    Span4Mux_s0_h I__7251 (
            .O(N__29412),
            .I(N__29384));
    InMux I__7250 (
            .O(N__29411),
            .I(N__29381));
    LocalMux I__7249 (
            .O(N__29408),
            .I(N__29378));
    Span4Mux_h I__7248 (
            .O(N__29405),
            .I(N__29371));
    Span4Mux_h I__7247 (
            .O(N__29398),
            .I(N__29371));
    LocalMux I__7246 (
            .O(N__29395),
            .I(N__29371));
    InMux I__7245 (
            .O(N__29394),
            .I(N__29368));
    InMux I__7244 (
            .O(N__29393),
            .I(N__29363));
    InMux I__7243 (
            .O(N__29392),
            .I(N__29363));
    Span4Mux_h I__7242 (
            .O(N__29387),
            .I(N__29358));
    Span4Mux_h I__7241 (
            .O(N__29384),
            .I(N__29358));
    LocalMux I__7240 (
            .O(N__29381),
            .I(N__29353));
    Span12Mux_s5_v I__7239 (
            .O(N__29378),
            .I(N__29353));
    Odrv4 I__7238 (
            .O(N__29371),
            .I(\tok.n2616 ));
    LocalMux I__7237 (
            .O(N__29368),
            .I(\tok.n2616 ));
    LocalMux I__7236 (
            .O(N__29363),
            .I(\tok.n2616 ));
    Odrv4 I__7235 (
            .O(N__29358),
            .I(\tok.n2616 ));
    Odrv12 I__7234 (
            .O(N__29353),
            .I(\tok.n2616 ));
    InMux I__7233 (
            .O(N__29342),
            .I(N__29339));
    LocalMux I__7232 (
            .O(N__29339),
            .I(N__29336));
    Span4Mux_h I__7231 (
            .O(N__29336),
            .I(N__29333));
    Span4Mux_h I__7230 (
            .O(N__29333),
            .I(N__29330));
    Odrv4 I__7229 (
            .O(N__29330),
            .I(\tok.n15_adj_680 ));
    CascadeMux I__7228 (
            .O(N__29327),
            .I(N__29323));
    CascadeMux I__7227 (
            .O(N__29326),
            .I(N__29318));
    InMux I__7226 (
            .O(N__29323),
            .I(N__29306));
    InMux I__7225 (
            .O(N__29322),
            .I(N__29306));
    InMux I__7224 (
            .O(N__29321),
            .I(N__29306));
    InMux I__7223 (
            .O(N__29318),
            .I(N__29306));
    InMux I__7222 (
            .O(N__29317),
            .I(N__29306));
    LocalMux I__7221 (
            .O(N__29306),
            .I(N__29301));
    InMux I__7220 (
            .O(N__29305),
            .I(N__29298));
    InMux I__7219 (
            .O(N__29304),
            .I(N__29295));
    Span4Mux_h I__7218 (
            .O(N__29301),
            .I(N__29286));
    LocalMux I__7217 (
            .O(N__29298),
            .I(N__29286));
    LocalMux I__7216 (
            .O(N__29295),
            .I(N__29275));
    InMux I__7215 (
            .O(N__29294),
            .I(N__29268));
    InMux I__7214 (
            .O(N__29293),
            .I(N__29268));
    InMux I__7213 (
            .O(N__29292),
            .I(N__29268));
    CascadeMux I__7212 (
            .O(N__29291),
            .I(N__29262));
    Span4Mux_v I__7211 (
            .O(N__29286),
            .I(N__29255));
    InMux I__7210 (
            .O(N__29285),
            .I(N__29252));
    CascadeMux I__7209 (
            .O(N__29284),
            .I(N__29248));
    InMux I__7208 (
            .O(N__29283),
            .I(N__29236));
    InMux I__7207 (
            .O(N__29282),
            .I(N__29236));
    InMux I__7206 (
            .O(N__29281),
            .I(N__29236));
    InMux I__7205 (
            .O(N__29280),
            .I(N__29236));
    InMux I__7204 (
            .O(N__29279),
            .I(N__29236));
    InMux I__7203 (
            .O(N__29278),
            .I(N__29233));
    Span4Mux_h I__7202 (
            .O(N__29275),
            .I(N__29230));
    LocalMux I__7201 (
            .O(N__29268),
            .I(N__29227));
    CascadeMux I__7200 (
            .O(N__29267),
            .I(N__29223));
    CascadeMux I__7199 (
            .O(N__29266),
            .I(N__29218));
    InMux I__7198 (
            .O(N__29265),
            .I(N__29209));
    InMux I__7197 (
            .O(N__29262),
            .I(N__29209));
    InMux I__7196 (
            .O(N__29261),
            .I(N__29209));
    InMux I__7195 (
            .O(N__29260),
            .I(N__29209));
    InMux I__7194 (
            .O(N__29259),
            .I(N__29204));
    InMux I__7193 (
            .O(N__29258),
            .I(N__29204));
    Span4Mux_h I__7192 (
            .O(N__29255),
            .I(N__29199));
    LocalMux I__7191 (
            .O(N__29252),
            .I(N__29199));
    InMux I__7190 (
            .O(N__29251),
            .I(N__29192));
    InMux I__7189 (
            .O(N__29248),
            .I(N__29192));
    InMux I__7188 (
            .O(N__29247),
            .I(N__29192));
    LocalMux I__7187 (
            .O(N__29236),
            .I(N__29189));
    LocalMux I__7186 (
            .O(N__29233),
            .I(N__29186));
    Span4Mux_h I__7185 (
            .O(N__29230),
            .I(N__29181));
    Span4Mux_h I__7184 (
            .O(N__29227),
            .I(N__29181));
    InMux I__7183 (
            .O(N__29226),
            .I(N__29170));
    InMux I__7182 (
            .O(N__29223),
            .I(N__29170));
    InMux I__7181 (
            .O(N__29222),
            .I(N__29170));
    InMux I__7180 (
            .O(N__29221),
            .I(N__29170));
    InMux I__7179 (
            .O(N__29218),
            .I(N__29170));
    LocalMux I__7178 (
            .O(N__29209),
            .I(N__29165));
    LocalMux I__7177 (
            .O(N__29204),
            .I(N__29165));
    Span4Mux_h I__7176 (
            .O(N__29199),
            .I(N__29162));
    LocalMux I__7175 (
            .O(N__29192),
            .I(N__29155));
    Span4Mux_h I__7174 (
            .O(N__29189),
            .I(N__29155));
    Span4Mux_v I__7173 (
            .O(N__29186),
            .I(N__29155));
    Sp12to4 I__7172 (
            .O(N__29181),
            .I(N__29150));
    LocalMux I__7171 (
            .O(N__29170),
            .I(N__29150));
    Span12Mux_h I__7170 (
            .O(N__29165),
            .I(N__29146));
    Span4Mux_v I__7169 (
            .O(N__29162),
            .I(N__29143));
    Sp12to4 I__7168 (
            .O(N__29155),
            .I(N__29138));
    Span12Mux_s7_v I__7167 (
            .O(N__29150),
            .I(N__29138));
    InMux I__7166 (
            .O(N__29149),
            .I(N__29135));
    Odrv12 I__7165 (
            .O(N__29146),
            .I(\tok.n14_adj_658 ));
    Odrv4 I__7164 (
            .O(N__29143),
            .I(\tok.n14_adj_658 ));
    Odrv12 I__7163 (
            .O(N__29138),
            .I(\tok.n14_adj_658 ));
    LocalMux I__7162 (
            .O(N__29135),
            .I(\tok.n14_adj_658 ));
    InMux I__7161 (
            .O(N__29126),
            .I(N__29123));
    LocalMux I__7160 (
            .O(N__29123),
            .I(N__29118));
    InMux I__7159 (
            .O(N__29122),
            .I(N__29113));
    InMux I__7158 (
            .O(N__29121),
            .I(N__29113));
    Odrv4 I__7157 (
            .O(N__29118),
            .I(\tok.n11_adj_649 ));
    LocalMux I__7156 (
            .O(N__29113),
            .I(\tok.n11_adj_649 ));
    InMux I__7155 (
            .O(N__29108),
            .I(N__29096));
    InMux I__7154 (
            .O(N__29107),
            .I(N__29096));
    InMux I__7153 (
            .O(N__29106),
            .I(N__29085));
    InMux I__7152 (
            .O(N__29105),
            .I(N__29085));
    InMux I__7151 (
            .O(N__29104),
            .I(N__29085));
    InMux I__7150 (
            .O(N__29103),
            .I(N__29085));
    InMux I__7149 (
            .O(N__29102),
            .I(N__29085));
    SRMux I__7148 (
            .O(N__29101),
            .I(N__29082));
    LocalMux I__7147 (
            .O(N__29096),
            .I(N__29072));
    LocalMux I__7146 (
            .O(N__29085),
            .I(N__29072));
    LocalMux I__7145 (
            .O(N__29082),
            .I(N__29069));
    InMux I__7144 (
            .O(N__29081),
            .I(N__29064));
    InMux I__7143 (
            .O(N__29080),
            .I(N__29064));
    InMux I__7142 (
            .O(N__29079),
            .I(N__29057));
    InMux I__7141 (
            .O(N__29078),
            .I(N__29057));
    InMux I__7140 (
            .O(N__29077),
            .I(N__29057));
    Span4Mux_h I__7139 (
            .O(N__29072),
            .I(N__29054));
    Span4Mux_h I__7138 (
            .O(N__29069),
            .I(N__29051));
    LocalMux I__7137 (
            .O(N__29064),
            .I(N__29046));
    LocalMux I__7136 (
            .O(N__29057),
            .I(N__29046));
    Span4Mux_h I__7135 (
            .O(N__29054),
            .I(N__29043));
    Odrv4 I__7134 (
            .O(N__29051),
            .I(\tok.write_flag ));
    Odrv12 I__7133 (
            .O(N__29046),
            .I(\tok.write_flag ));
    Odrv4 I__7132 (
            .O(N__29043),
            .I(\tok.write_flag ));
    InMux I__7131 (
            .O(N__29036),
            .I(N__29022));
    InMux I__7130 (
            .O(N__29035),
            .I(N__29019));
    InMux I__7129 (
            .O(N__29034),
            .I(N__29010));
    InMux I__7128 (
            .O(N__29033),
            .I(N__29010));
    InMux I__7127 (
            .O(N__29032),
            .I(N__29010));
    InMux I__7126 (
            .O(N__29031),
            .I(N__29010));
    InMux I__7125 (
            .O(N__29030),
            .I(N__29000));
    InMux I__7124 (
            .O(N__29029),
            .I(N__29000));
    InMux I__7123 (
            .O(N__29028),
            .I(N__29000));
    InMux I__7122 (
            .O(N__29027),
            .I(N__28991));
    InMux I__7121 (
            .O(N__29026),
            .I(N__28991));
    InMux I__7120 (
            .O(N__29025),
            .I(N__28991));
    LocalMux I__7119 (
            .O(N__29022),
            .I(N__28986));
    LocalMux I__7118 (
            .O(N__29019),
            .I(N__28981));
    LocalMux I__7117 (
            .O(N__29010),
            .I(N__28981));
    InMux I__7116 (
            .O(N__29009),
            .I(N__28974));
    InMux I__7115 (
            .O(N__29008),
            .I(N__28974));
    InMux I__7114 (
            .O(N__29007),
            .I(N__28974));
    LocalMux I__7113 (
            .O(N__29000),
            .I(N__28968));
    InMux I__7112 (
            .O(N__28999),
            .I(N__28963));
    InMux I__7111 (
            .O(N__28998),
            .I(N__28963));
    LocalMux I__7110 (
            .O(N__28991),
            .I(N__28959));
    InMux I__7109 (
            .O(N__28990),
            .I(N__28956));
    InMux I__7108 (
            .O(N__28989),
            .I(N__28953));
    Span4Mux_h I__7107 (
            .O(N__28986),
            .I(N__28950));
    Span4Mux_s2_v I__7106 (
            .O(N__28981),
            .I(N__28945));
    LocalMux I__7105 (
            .O(N__28974),
            .I(N__28945));
    InMux I__7104 (
            .O(N__28973),
            .I(N__28942));
    InMux I__7103 (
            .O(N__28972),
            .I(N__28936));
    InMux I__7102 (
            .O(N__28971),
            .I(N__28931));
    Span4Mux_v I__7101 (
            .O(N__28968),
            .I(N__28926));
    LocalMux I__7100 (
            .O(N__28963),
            .I(N__28926));
    InMux I__7099 (
            .O(N__28962),
            .I(N__28923));
    Span4Mux_h I__7098 (
            .O(N__28959),
            .I(N__28920));
    LocalMux I__7097 (
            .O(N__28956),
            .I(N__28917));
    LocalMux I__7096 (
            .O(N__28953),
            .I(N__28914));
    Span4Mux_h I__7095 (
            .O(N__28950),
            .I(N__28907));
    Span4Mux_v I__7094 (
            .O(N__28945),
            .I(N__28907));
    LocalMux I__7093 (
            .O(N__28942),
            .I(N__28907));
    InMux I__7092 (
            .O(N__28941),
            .I(N__28900));
    InMux I__7091 (
            .O(N__28940),
            .I(N__28895));
    InMux I__7090 (
            .O(N__28939),
            .I(N__28895));
    LocalMux I__7089 (
            .O(N__28936),
            .I(N__28892));
    InMux I__7088 (
            .O(N__28935),
            .I(N__28887));
    InMux I__7087 (
            .O(N__28934),
            .I(N__28887));
    LocalMux I__7086 (
            .O(N__28931),
            .I(N__28884));
    Span4Mux_h I__7085 (
            .O(N__28926),
            .I(N__28881));
    LocalMux I__7084 (
            .O(N__28923),
            .I(N__28876));
    Span4Mux_h I__7083 (
            .O(N__28920),
            .I(N__28876));
    Span4Mux_v I__7082 (
            .O(N__28917),
            .I(N__28869));
    Span4Mux_v I__7081 (
            .O(N__28914),
            .I(N__28869));
    Span4Mux_v I__7080 (
            .O(N__28907),
            .I(N__28869));
    InMux I__7079 (
            .O(N__28906),
            .I(N__28866));
    InMux I__7078 (
            .O(N__28905),
            .I(N__28859));
    InMux I__7077 (
            .O(N__28904),
            .I(N__28859));
    InMux I__7076 (
            .O(N__28903),
            .I(N__28859));
    LocalMux I__7075 (
            .O(N__28900),
            .I(N__28850));
    LocalMux I__7074 (
            .O(N__28895),
            .I(N__28850));
    Span12Mux_s6_v I__7073 (
            .O(N__28892),
            .I(N__28850));
    LocalMux I__7072 (
            .O(N__28887),
            .I(N__28850));
    Odrv4 I__7071 (
            .O(N__28884),
            .I(\tok.T_4 ));
    Odrv4 I__7070 (
            .O(N__28881),
            .I(\tok.T_4 ));
    Odrv4 I__7069 (
            .O(N__28876),
            .I(\tok.T_4 ));
    Odrv4 I__7068 (
            .O(N__28869),
            .I(\tok.T_4 ));
    LocalMux I__7067 (
            .O(N__28866),
            .I(\tok.T_4 ));
    LocalMux I__7066 (
            .O(N__28859),
            .I(\tok.T_4 ));
    Odrv12 I__7065 (
            .O(N__28850),
            .I(\tok.T_4 ));
    InMux I__7064 (
            .O(N__28835),
            .I(N__28823));
    InMux I__7063 (
            .O(N__28834),
            .I(N__28823));
    InMux I__7062 (
            .O(N__28833),
            .I(N__28816));
    InMux I__7061 (
            .O(N__28832),
            .I(N__28816));
    CascadeMux I__7060 (
            .O(N__28831),
            .I(N__28813));
    InMux I__7059 (
            .O(N__28830),
            .I(N__28809));
    InMux I__7058 (
            .O(N__28829),
            .I(N__28804));
    InMux I__7057 (
            .O(N__28828),
            .I(N__28801));
    LocalMux I__7056 (
            .O(N__28823),
            .I(N__28798));
    InMux I__7055 (
            .O(N__28822),
            .I(N__28793));
    InMux I__7054 (
            .O(N__28821),
            .I(N__28793));
    LocalMux I__7053 (
            .O(N__28816),
            .I(N__28790));
    InMux I__7052 (
            .O(N__28813),
            .I(N__28785));
    InMux I__7051 (
            .O(N__28812),
            .I(N__28785));
    LocalMux I__7050 (
            .O(N__28809),
            .I(N__28782));
    InMux I__7049 (
            .O(N__28808),
            .I(N__28779));
    CascadeMux I__7048 (
            .O(N__28807),
            .I(N__28776));
    LocalMux I__7047 (
            .O(N__28804),
            .I(N__28770));
    LocalMux I__7046 (
            .O(N__28801),
            .I(N__28767));
    Span4Mux_h I__7045 (
            .O(N__28798),
            .I(N__28764));
    LocalMux I__7044 (
            .O(N__28793),
            .I(N__28757));
    Span4Mux_v I__7043 (
            .O(N__28790),
            .I(N__28757));
    LocalMux I__7042 (
            .O(N__28785),
            .I(N__28757));
    Span4Mux_s3_h I__7041 (
            .O(N__28782),
            .I(N__28752));
    LocalMux I__7040 (
            .O(N__28779),
            .I(N__28752));
    InMux I__7039 (
            .O(N__28776),
            .I(N__28747));
    InMux I__7038 (
            .O(N__28775),
            .I(N__28747));
    CascadeMux I__7037 (
            .O(N__28774),
            .I(N__28743));
    CascadeMux I__7036 (
            .O(N__28773),
            .I(N__28740));
    Span4Mux_h I__7035 (
            .O(N__28770),
            .I(N__28736));
    Span4Mux_h I__7034 (
            .O(N__28767),
            .I(N__28733));
    Span4Mux_h I__7033 (
            .O(N__28764),
            .I(N__28728));
    Span4Mux_h I__7032 (
            .O(N__28757),
            .I(N__28728));
    Span4Mux_v I__7031 (
            .O(N__28752),
            .I(N__28723));
    LocalMux I__7030 (
            .O(N__28747),
            .I(N__28723));
    InMux I__7029 (
            .O(N__28746),
            .I(N__28720));
    InMux I__7028 (
            .O(N__28743),
            .I(N__28713));
    InMux I__7027 (
            .O(N__28740),
            .I(N__28713));
    InMux I__7026 (
            .O(N__28739),
            .I(N__28713));
    Odrv4 I__7025 (
            .O(N__28736),
            .I(\tok.T_7 ));
    Odrv4 I__7024 (
            .O(N__28733),
            .I(\tok.T_7 ));
    Odrv4 I__7023 (
            .O(N__28728),
            .I(\tok.T_7 ));
    Odrv4 I__7022 (
            .O(N__28723),
            .I(\tok.T_7 ));
    LocalMux I__7021 (
            .O(N__28720),
            .I(\tok.T_7 ));
    LocalMux I__7020 (
            .O(N__28713),
            .I(\tok.T_7 ));
    CascadeMux I__7019 (
            .O(N__28700),
            .I(N__28694));
    CascadeMux I__7018 (
            .O(N__28699),
            .I(N__28686));
    InMux I__7017 (
            .O(N__28698),
            .I(N__28683));
    InMux I__7016 (
            .O(N__28697),
            .I(N__28680));
    InMux I__7015 (
            .O(N__28694),
            .I(N__28671));
    InMux I__7014 (
            .O(N__28693),
            .I(N__28671));
    InMux I__7013 (
            .O(N__28692),
            .I(N__28671));
    InMux I__7012 (
            .O(N__28691),
            .I(N__28668));
    InMux I__7011 (
            .O(N__28690),
            .I(N__28663));
    InMux I__7010 (
            .O(N__28689),
            .I(N__28663));
    InMux I__7009 (
            .O(N__28686),
            .I(N__28659));
    LocalMux I__7008 (
            .O(N__28683),
            .I(N__28655));
    LocalMux I__7007 (
            .O(N__28680),
            .I(N__28652));
    InMux I__7006 (
            .O(N__28679),
            .I(N__28649));
    InMux I__7005 (
            .O(N__28678),
            .I(N__28646));
    LocalMux I__7004 (
            .O(N__28671),
            .I(N__28643));
    LocalMux I__7003 (
            .O(N__28668),
            .I(N__28638));
    LocalMux I__7002 (
            .O(N__28663),
            .I(N__28638));
    InMux I__7001 (
            .O(N__28662),
            .I(N__28635));
    LocalMux I__7000 (
            .O(N__28659),
            .I(N__28631));
    InMux I__6999 (
            .O(N__28658),
            .I(N__28628));
    Span4Mux_s3_v I__6998 (
            .O(N__28655),
            .I(N__28622));
    Span4Mux_s2_v I__6997 (
            .O(N__28652),
            .I(N__28617));
    LocalMux I__6996 (
            .O(N__28649),
            .I(N__28617));
    LocalMux I__6995 (
            .O(N__28646),
            .I(N__28608));
    Span4Mux_v I__6994 (
            .O(N__28643),
            .I(N__28608));
    Span4Mux_v I__6993 (
            .O(N__28638),
            .I(N__28608));
    LocalMux I__6992 (
            .O(N__28635),
            .I(N__28608));
    CascadeMux I__6991 (
            .O(N__28634),
            .I(N__28605));
    Span4Mux_s3_h I__6990 (
            .O(N__28631),
            .I(N__28600));
    LocalMux I__6989 (
            .O(N__28628),
            .I(N__28600));
    InMux I__6988 (
            .O(N__28627),
            .I(N__28595));
    InMux I__6987 (
            .O(N__28626),
            .I(N__28595));
    CascadeMux I__6986 (
            .O(N__28625),
            .I(N__28591));
    Span4Mux_v I__6985 (
            .O(N__28622),
            .I(N__28585));
    Span4Mux_v I__6984 (
            .O(N__28617),
            .I(N__28585));
    Span4Mux_h I__6983 (
            .O(N__28608),
            .I(N__28582));
    InMux I__6982 (
            .O(N__28605),
            .I(N__28579));
    Span4Mux_v I__6981 (
            .O(N__28600),
            .I(N__28574));
    LocalMux I__6980 (
            .O(N__28595),
            .I(N__28574));
    InMux I__6979 (
            .O(N__28594),
            .I(N__28567));
    InMux I__6978 (
            .O(N__28591),
            .I(N__28567));
    InMux I__6977 (
            .O(N__28590),
            .I(N__28567));
    Odrv4 I__6976 (
            .O(N__28585),
            .I(\tok.T_5 ));
    Odrv4 I__6975 (
            .O(N__28582),
            .I(\tok.T_5 ));
    LocalMux I__6974 (
            .O(N__28579),
            .I(\tok.T_5 ));
    Odrv4 I__6973 (
            .O(N__28574),
            .I(\tok.T_5 ));
    LocalMux I__6972 (
            .O(N__28567),
            .I(\tok.T_5 ));
    InMux I__6971 (
            .O(N__28556),
            .I(N__28551));
    CascadeMux I__6970 (
            .O(N__28555),
            .I(N__28545));
    InMux I__6969 (
            .O(N__28554),
            .I(N__28539));
    LocalMux I__6968 (
            .O(N__28551),
            .I(N__28536));
    InMux I__6967 (
            .O(N__28550),
            .I(N__28533));
    InMux I__6966 (
            .O(N__28549),
            .I(N__28525));
    InMux I__6965 (
            .O(N__28548),
            .I(N__28518));
    InMux I__6964 (
            .O(N__28545),
            .I(N__28518));
    CascadeMux I__6963 (
            .O(N__28544),
            .I(N__28514));
    InMux I__6962 (
            .O(N__28543),
            .I(N__28509));
    InMux I__6961 (
            .O(N__28542),
            .I(N__28506));
    LocalMux I__6960 (
            .O(N__28539),
            .I(N__28501));
    Span4Mux_v I__6959 (
            .O(N__28536),
            .I(N__28498));
    LocalMux I__6958 (
            .O(N__28533),
            .I(N__28495));
    InMux I__6957 (
            .O(N__28532),
            .I(N__28492));
    InMux I__6956 (
            .O(N__28531),
            .I(N__28489));
    InMux I__6955 (
            .O(N__28530),
            .I(N__28486));
    InMux I__6954 (
            .O(N__28529),
            .I(N__28481));
    InMux I__6953 (
            .O(N__28528),
            .I(N__28481));
    LocalMux I__6952 (
            .O(N__28525),
            .I(N__28478));
    InMux I__6951 (
            .O(N__28524),
            .I(N__28473));
    InMux I__6950 (
            .O(N__28523),
            .I(N__28473));
    LocalMux I__6949 (
            .O(N__28518),
            .I(N__28470));
    InMux I__6948 (
            .O(N__28517),
            .I(N__28465));
    InMux I__6947 (
            .O(N__28514),
            .I(N__28465));
    InMux I__6946 (
            .O(N__28513),
            .I(N__28460));
    InMux I__6945 (
            .O(N__28512),
            .I(N__28460));
    LocalMux I__6944 (
            .O(N__28509),
            .I(N__28454));
    LocalMux I__6943 (
            .O(N__28506),
            .I(N__28454));
    InMux I__6942 (
            .O(N__28505),
            .I(N__28451));
    InMux I__6941 (
            .O(N__28504),
            .I(N__28446));
    Span4Mux_v I__6940 (
            .O(N__28501),
            .I(N__28439));
    Span4Mux_s0_h I__6939 (
            .O(N__28498),
            .I(N__28439));
    Span4Mux_v I__6938 (
            .O(N__28495),
            .I(N__28439));
    LocalMux I__6937 (
            .O(N__28492),
            .I(N__28436));
    LocalMux I__6936 (
            .O(N__28489),
            .I(N__28431));
    LocalMux I__6935 (
            .O(N__28486),
            .I(N__28431));
    LocalMux I__6934 (
            .O(N__28481),
            .I(N__28428));
    Span4Mux_h I__6933 (
            .O(N__28478),
            .I(N__28417));
    LocalMux I__6932 (
            .O(N__28473),
            .I(N__28417));
    Span4Mux_h I__6931 (
            .O(N__28470),
            .I(N__28417));
    LocalMux I__6930 (
            .O(N__28465),
            .I(N__28417));
    LocalMux I__6929 (
            .O(N__28460),
            .I(N__28417));
    InMux I__6928 (
            .O(N__28459),
            .I(N__28413));
    Span4Mux_s3_h I__6927 (
            .O(N__28454),
            .I(N__28408));
    LocalMux I__6926 (
            .O(N__28451),
            .I(N__28408));
    InMux I__6925 (
            .O(N__28450),
            .I(N__28403));
    InMux I__6924 (
            .O(N__28449),
            .I(N__28403));
    LocalMux I__6923 (
            .O(N__28446),
            .I(N__28397));
    Sp12to4 I__6922 (
            .O(N__28439),
            .I(N__28394));
    Span4Mux_s2_h I__6921 (
            .O(N__28436),
            .I(N__28391));
    Span4Mux_h I__6920 (
            .O(N__28431),
            .I(N__28388));
    Span4Mux_v I__6919 (
            .O(N__28428),
            .I(N__28383));
    Span4Mux_v I__6918 (
            .O(N__28417),
            .I(N__28383));
    InMux I__6917 (
            .O(N__28416),
            .I(N__28380));
    LocalMux I__6916 (
            .O(N__28413),
            .I(N__28373));
    Span4Mux_v I__6915 (
            .O(N__28408),
            .I(N__28373));
    LocalMux I__6914 (
            .O(N__28403),
            .I(N__28373));
    InMux I__6913 (
            .O(N__28402),
            .I(N__28366));
    InMux I__6912 (
            .O(N__28401),
            .I(N__28366));
    InMux I__6911 (
            .O(N__28400),
            .I(N__28366));
    Odrv4 I__6910 (
            .O(N__28397),
            .I(\tok.T_6 ));
    Odrv12 I__6909 (
            .O(N__28394),
            .I(\tok.T_6 ));
    Odrv4 I__6908 (
            .O(N__28391),
            .I(\tok.T_6 ));
    Odrv4 I__6907 (
            .O(N__28388),
            .I(\tok.T_6 ));
    Odrv4 I__6906 (
            .O(N__28383),
            .I(\tok.T_6 ));
    LocalMux I__6905 (
            .O(N__28380),
            .I(\tok.T_6 ));
    Odrv4 I__6904 (
            .O(N__28373),
            .I(\tok.T_6 ));
    LocalMux I__6903 (
            .O(N__28366),
            .I(\tok.T_6 ));
    CascadeMux I__6902 (
            .O(N__28349),
            .I(N__28345));
    InMux I__6901 (
            .O(N__28348),
            .I(N__28341));
    InMux I__6900 (
            .O(N__28345),
            .I(N__28338));
    InMux I__6899 (
            .O(N__28344),
            .I(N__28334));
    LocalMux I__6898 (
            .O(N__28341),
            .I(N__28329));
    LocalMux I__6897 (
            .O(N__28338),
            .I(N__28329));
    InMux I__6896 (
            .O(N__28337),
            .I(N__28326));
    LocalMux I__6895 (
            .O(N__28334),
            .I(N__28316));
    Span4Mux_v I__6894 (
            .O(N__28329),
            .I(N__28316));
    LocalMux I__6893 (
            .O(N__28326),
            .I(N__28316));
    InMux I__6892 (
            .O(N__28325),
            .I(N__28313));
    InMux I__6891 (
            .O(N__28324),
            .I(N__28308));
    InMux I__6890 (
            .O(N__28323),
            .I(N__28308));
    Span4Mux_s3_v I__6889 (
            .O(N__28316),
            .I(N__28303));
    LocalMux I__6888 (
            .O(N__28313),
            .I(N__28303));
    LocalMux I__6887 (
            .O(N__28308),
            .I(N__28300));
    Span4Mux_h I__6886 (
            .O(N__28303),
            .I(N__28294));
    Span4Mux_s3_v I__6885 (
            .O(N__28300),
            .I(N__28294));
    InMux I__6884 (
            .O(N__28299),
            .I(N__28291));
    Span4Mux_h I__6883 (
            .O(N__28294),
            .I(N__28288));
    LocalMux I__6882 (
            .O(N__28291),
            .I(\tok.n8 ));
    Odrv4 I__6881 (
            .O(N__28288),
            .I(\tok.n8 ));
    InMux I__6880 (
            .O(N__28283),
            .I(N__28280));
    LocalMux I__6879 (
            .O(N__28280),
            .I(N__28277));
    Span4Mux_h I__6878 (
            .O(N__28277),
            .I(N__28274));
    Odrv4 I__6877 (
            .O(N__28274),
            .I(\tok.n18 ));
    InMux I__6876 (
            .O(N__28271),
            .I(N__28265));
    CascadeMux I__6875 (
            .O(N__28270),
            .I(N__28261));
    InMux I__6874 (
            .O(N__28269),
            .I(N__28256));
    InMux I__6873 (
            .O(N__28268),
            .I(N__28248));
    LocalMux I__6872 (
            .O(N__28265),
            .I(N__28245));
    InMux I__6871 (
            .O(N__28264),
            .I(N__28242));
    InMux I__6870 (
            .O(N__28261),
            .I(N__28239));
    InMux I__6869 (
            .O(N__28260),
            .I(N__28236));
    InMux I__6868 (
            .O(N__28259),
            .I(N__28233));
    LocalMux I__6867 (
            .O(N__28256),
            .I(N__28229));
    InMux I__6866 (
            .O(N__28255),
            .I(N__28226));
    InMux I__6865 (
            .O(N__28254),
            .I(N__28223));
    InMux I__6864 (
            .O(N__28253),
            .I(N__28220));
    InMux I__6863 (
            .O(N__28252),
            .I(N__28213));
    InMux I__6862 (
            .O(N__28251),
            .I(N__28213));
    LocalMux I__6861 (
            .O(N__28248),
            .I(N__28210));
    Span4Mux_v I__6860 (
            .O(N__28245),
            .I(N__28207));
    LocalMux I__6859 (
            .O(N__28242),
            .I(N__28202));
    LocalMux I__6858 (
            .O(N__28239),
            .I(N__28202));
    LocalMux I__6857 (
            .O(N__28236),
            .I(N__28199));
    LocalMux I__6856 (
            .O(N__28233),
            .I(N__28196));
    InMux I__6855 (
            .O(N__28232),
            .I(N__28193));
    Span4Mux_v I__6854 (
            .O(N__28229),
            .I(N__28184));
    LocalMux I__6853 (
            .O(N__28226),
            .I(N__28184));
    LocalMux I__6852 (
            .O(N__28223),
            .I(N__28184));
    LocalMux I__6851 (
            .O(N__28220),
            .I(N__28184));
    InMux I__6850 (
            .O(N__28219),
            .I(N__28179));
    InMux I__6849 (
            .O(N__28218),
            .I(N__28179));
    LocalMux I__6848 (
            .O(N__28213),
            .I(N__28176));
    Span4Mux_v I__6847 (
            .O(N__28210),
            .I(N__28165));
    Span4Mux_h I__6846 (
            .O(N__28207),
            .I(N__28165));
    Span4Mux_v I__6845 (
            .O(N__28202),
            .I(N__28165));
    Span4Mux_s3_h I__6844 (
            .O(N__28199),
            .I(N__28165));
    Span4Mux_v I__6843 (
            .O(N__28196),
            .I(N__28165));
    LocalMux I__6842 (
            .O(N__28193),
            .I(N__28162));
    Span4Mux_h I__6841 (
            .O(N__28184),
            .I(N__28159));
    LocalMux I__6840 (
            .O(N__28179),
            .I(\tok.A_low_6 ));
    Odrv4 I__6839 (
            .O(N__28176),
            .I(\tok.A_low_6 ));
    Odrv4 I__6838 (
            .O(N__28165),
            .I(\tok.A_low_6 ));
    Odrv4 I__6837 (
            .O(N__28162),
            .I(\tok.A_low_6 ));
    Odrv4 I__6836 (
            .O(N__28159),
            .I(\tok.A_low_6 ));
    CascadeMux I__6835 (
            .O(N__28148),
            .I(N__28145));
    InMux I__6834 (
            .O(N__28145),
            .I(N__28142));
    LocalMux I__6833 (
            .O(N__28142),
            .I(N__28139));
    Span4Mux_v I__6832 (
            .O(N__28139),
            .I(N__28136));
    Span4Mux_h I__6831 (
            .O(N__28136),
            .I(N__28133));
    Odrv4 I__6830 (
            .O(N__28133),
            .I(\tok.n179 ));
    InMux I__6829 (
            .O(N__28130),
            .I(N__28127));
    LocalMux I__6828 (
            .O(N__28127),
            .I(N__28124));
    Span4Mux_h I__6827 (
            .O(N__28124),
            .I(N__28121));
    Odrv4 I__6826 (
            .O(N__28121),
            .I(\tok.n10_adj_675 ));
    InMux I__6825 (
            .O(N__28118),
            .I(N__28111));
    InMux I__6824 (
            .O(N__28117),
            .I(N__28111));
    InMux I__6823 (
            .O(N__28116),
            .I(N__28108));
    LocalMux I__6822 (
            .O(N__28111),
            .I(N__28105));
    LocalMux I__6821 (
            .O(N__28108),
            .I(N__28099));
    Span4Mux_h I__6820 (
            .O(N__28105),
            .I(N__28096));
    InMux I__6819 (
            .O(N__28104),
            .I(N__28093));
    InMux I__6818 (
            .O(N__28103),
            .I(N__28088));
    InMux I__6817 (
            .O(N__28102),
            .I(N__28088));
    Odrv4 I__6816 (
            .O(N__28099),
            .I(\tok.n9 ));
    Odrv4 I__6815 (
            .O(N__28096),
            .I(\tok.n9 ));
    LocalMux I__6814 (
            .O(N__28093),
            .I(\tok.n9 ));
    LocalMux I__6813 (
            .O(N__28088),
            .I(\tok.n9 ));
    CascadeMux I__6812 (
            .O(N__28079),
            .I(\tok.n10_adj_675_cascade_ ));
    InMux I__6811 (
            .O(N__28076),
            .I(N__28068));
    InMux I__6810 (
            .O(N__28075),
            .I(N__28068));
    InMux I__6809 (
            .O(N__28074),
            .I(N__28065));
    InMux I__6808 (
            .O(N__28073),
            .I(N__28062));
    LocalMux I__6807 (
            .O(N__28068),
            .I(N__28059));
    LocalMux I__6806 (
            .O(N__28065),
            .I(N__28051));
    LocalMux I__6805 (
            .O(N__28062),
            .I(N__28048));
    Span4Mux_h I__6804 (
            .O(N__28059),
            .I(N__28045));
    InMux I__6803 (
            .O(N__28058),
            .I(N__28040));
    InMux I__6802 (
            .O(N__28057),
            .I(N__28040));
    InMux I__6801 (
            .O(N__28056),
            .I(N__28037));
    InMux I__6800 (
            .O(N__28055),
            .I(N__28032));
    InMux I__6799 (
            .O(N__28054),
            .I(N__28032));
    Odrv12 I__6798 (
            .O(N__28051),
            .I(\tok.n2586 ));
    Odrv4 I__6797 (
            .O(N__28048),
            .I(\tok.n2586 ));
    Odrv4 I__6796 (
            .O(N__28045),
            .I(\tok.n2586 ));
    LocalMux I__6795 (
            .O(N__28040),
            .I(\tok.n2586 ));
    LocalMux I__6794 (
            .O(N__28037),
            .I(\tok.n2586 ));
    LocalMux I__6793 (
            .O(N__28032),
            .I(\tok.n2586 ));
    InMux I__6792 (
            .O(N__28019),
            .I(N__28008));
    InMux I__6791 (
            .O(N__28018),
            .I(N__28005));
    InMux I__6790 (
            .O(N__28017),
            .I(N__28002));
    InMux I__6789 (
            .O(N__28016),
            .I(N__27994));
    InMux I__6788 (
            .O(N__28015),
            .I(N__27994));
    InMux I__6787 (
            .O(N__28014),
            .I(N__27989));
    CascadeMux I__6786 (
            .O(N__28013),
            .I(N__27983));
    CascadeMux I__6785 (
            .O(N__28012),
            .I(N__27980));
    CascadeMux I__6784 (
            .O(N__28011),
            .I(N__27976));
    LocalMux I__6783 (
            .O(N__28008),
            .I(N__27969));
    LocalMux I__6782 (
            .O(N__28005),
            .I(N__27969));
    LocalMux I__6781 (
            .O(N__28002),
            .I(N__27969));
    InMux I__6780 (
            .O(N__28001),
            .I(N__27966));
    InMux I__6779 (
            .O(N__28000),
            .I(N__27963));
    InMux I__6778 (
            .O(N__27999),
            .I(N__27960));
    LocalMux I__6777 (
            .O(N__27994),
            .I(N__27957));
    InMux I__6776 (
            .O(N__27993),
            .I(N__27952));
    InMux I__6775 (
            .O(N__27992),
            .I(N__27952));
    LocalMux I__6774 (
            .O(N__27989),
            .I(N__27949));
    InMux I__6773 (
            .O(N__27988),
            .I(N__27946));
    InMux I__6772 (
            .O(N__27987),
            .I(N__27939));
    InMux I__6771 (
            .O(N__27986),
            .I(N__27939));
    InMux I__6770 (
            .O(N__27983),
            .I(N__27939));
    InMux I__6769 (
            .O(N__27980),
            .I(N__27936));
    InMux I__6768 (
            .O(N__27979),
            .I(N__27931));
    InMux I__6767 (
            .O(N__27976),
            .I(N__27931));
    Span4Mux_s3_v I__6766 (
            .O(N__27969),
            .I(N__27920));
    LocalMux I__6765 (
            .O(N__27966),
            .I(N__27915));
    LocalMux I__6764 (
            .O(N__27963),
            .I(N__27915));
    LocalMux I__6763 (
            .O(N__27960),
            .I(N__27908));
    Span4Mux_v I__6762 (
            .O(N__27957),
            .I(N__27908));
    LocalMux I__6761 (
            .O(N__27952),
            .I(N__27908));
    Span4Mux_v I__6760 (
            .O(N__27949),
            .I(N__27905));
    LocalMux I__6759 (
            .O(N__27946),
            .I(N__27900));
    LocalMux I__6758 (
            .O(N__27939),
            .I(N__27900));
    LocalMux I__6757 (
            .O(N__27936),
            .I(N__27897));
    LocalMux I__6756 (
            .O(N__27931),
            .I(N__27894));
    CascadeMux I__6755 (
            .O(N__27930),
            .I(N__27891));
    CascadeMux I__6754 (
            .O(N__27929),
            .I(N__27888));
    CascadeMux I__6753 (
            .O(N__27928),
            .I(N__27885));
    CascadeMux I__6752 (
            .O(N__27927),
            .I(N__27881));
    CascadeMux I__6751 (
            .O(N__27926),
            .I(N__27876));
    CascadeMux I__6750 (
            .O(N__27925),
            .I(N__27873));
    CascadeMux I__6749 (
            .O(N__27924),
            .I(N__27870));
    CascadeMux I__6748 (
            .O(N__27923),
            .I(N__27865));
    Span4Mux_v I__6747 (
            .O(N__27920),
            .I(N__27860));
    Span4Mux_v I__6746 (
            .O(N__27915),
            .I(N__27860));
    Span4Mux_h I__6745 (
            .O(N__27908),
            .I(N__27857));
    Span4Mux_h I__6744 (
            .O(N__27905),
            .I(N__27848));
    Span4Mux_v I__6743 (
            .O(N__27900),
            .I(N__27848));
    Span4Mux_v I__6742 (
            .O(N__27897),
            .I(N__27848));
    Span4Mux_v I__6741 (
            .O(N__27894),
            .I(N__27848));
    InMux I__6740 (
            .O(N__27891),
            .I(N__27841));
    InMux I__6739 (
            .O(N__27888),
            .I(N__27841));
    InMux I__6738 (
            .O(N__27885),
            .I(N__27841));
    InMux I__6737 (
            .O(N__27884),
            .I(N__27834));
    InMux I__6736 (
            .O(N__27881),
            .I(N__27834));
    InMux I__6735 (
            .O(N__27880),
            .I(N__27834));
    InMux I__6734 (
            .O(N__27879),
            .I(N__27819));
    InMux I__6733 (
            .O(N__27876),
            .I(N__27819));
    InMux I__6732 (
            .O(N__27873),
            .I(N__27819));
    InMux I__6731 (
            .O(N__27870),
            .I(N__27819));
    InMux I__6730 (
            .O(N__27869),
            .I(N__27819));
    InMux I__6729 (
            .O(N__27868),
            .I(N__27819));
    InMux I__6728 (
            .O(N__27865),
            .I(N__27819));
    Odrv4 I__6727 (
            .O(N__27860),
            .I(\tok.T_3 ));
    Odrv4 I__6726 (
            .O(N__27857),
            .I(\tok.T_3 ));
    Odrv4 I__6725 (
            .O(N__27848),
            .I(\tok.T_3 ));
    LocalMux I__6724 (
            .O(N__27841),
            .I(\tok.T_3 ));
    LocalMux I__6723 (
            .O(N__27834),
            .I(\tok.T_3 ));
    LocalMux I__6722 (
            .O(N__27819),
            .I(\tok.T_3 ));
    InMux I__6721 (
            .O(N__27806),
            .I(N__27801));
    InMux I__6720 (
            .O(N__27805),
            .I(N__27796));
    InMux I__6719 (
            .O(N__27804),
            .I(N__27796));
    LocalMux I__6718 (
            .O(N__27801),
            .I(N__27791));
    LocalMux I__6717 (
            .O(N__27796),
            .I(N__27788));
    InMux I__6716 (
            .O(N__27795),
            .I(N__27785));
    InMux I__6715 (
            .O(N__27794),
            .I(N__27782));
    Span4Mux_h I__6714 (
            .O(N__27791),
            .I(N__27777));
    Span4Mux_h I__6713 (
            .O(N__27788),
            .I(N__27774));
    LocalMux I__6712 (
            .O(N__27785),
            .I(N__27771));
    LocalMux I__6711 (
            .O(N__27782),
            .I(N__27768));
    InMux I__6710 (
            .O(N__27781),
            .I(N__27763));
    InMux I__6709 (
            .O(N__27780),
            .I(N__27763));
    Span4Mux_h I__6708 (
            .O(N__27777),
            .I(N__27759));
    Span4Mux_h I__6707 (
            .O(N__27774),
            .I(N__27756));
    Span4Mux_v I__6706 (
            .O(N__27771),
            .I(N__27749));
    Span4Mux_v I__6705 (
            .O(N__27768),
            .I(N__27749));
    LocalMux I__6704 (
            .O(N__27763),
            .I(N__27749));
    InMux I__6703 (
            .O(N__27762),
            .I(N__27746));
    Odrv4 I__6702 (
            .O(N__27759),
            .I(\tok.n2178 ));
    Odrv4 I__6701 (
            .O(N__27756),
            .I(\tok.n2178 ));
    Odrv4 I__6700 (
            .O(N__27749),
            .I(\tok.n2178 ));
    LocalMux I__6699 (
            .O(N__27746),
            .I(\tok.n2178 ));
    InMux I__6698 (
            .O(N__27737),
            .I(N__27734));
    LocalMux I__6697 (
            .O(N__27734),
            .I(N__27731));
    Odrv12 I__6696 (
            .O(N__27731),
            .I(\tok.n41 ));
    InMux I__6695 (
            .O(N__27728),
            .I(N__27725));
    LocalMux I__6694 (
            .O(N__27725),
            .I(\tok.n4484 ));
    CascadeMux I__6693 (
            .O(N__27722),
            .I(N__27719));
    InMux I__6692 (
            .O(N__27719),
            .I(N__27716));
    LocalMux I__6691 (
            .O(N__27716),
            .I(\tok.n40_adj_661 ));
    InMux I__6690 (
            .O(N__27713),
            .I(N__27710));
    LocalMux I__6689 (
            .O(N__27710),
            .I(N__27707));
    Odrv12 I__6688 (
            .O(N__27707),
            .I(\tok.n42 ));
    InMux I__6687 (
            .O(N__27704),
            .I(N__27701));
    LocalMux I__6686 (
            .O(N__27701),
            .I(\tok.n4688 ));
    InMux I__6685 (
            .O(N__27698),
            .I(N__27695));
    LocalMux I__6684 (
            .O(N__27695),
            .I(N__27692));
    Span4Mux_s3_h I__6683 (
            .O(N__27692),
            .I(N__27687));
    InMux I__6682 (
            .O(N__27691),
            .I(N__27684));
    InMux I__6681 (
            .O(N__27690),
            .I(N__27681));
    Span4Mux_v I__6680 (
            .O(N__27687),
            .I(N__27676));
    LocalMux I__6679 (
            .O(N__27684),
            .I(N__27676));
    LocalMux I__6678 (
            .O(N__27681),
            .I(\tok.n10 ));
    Odrv4 I__6677 (
            .O(N__27676),
            .I(\tok.n10 ));
    CascadeMux I__6676 (
            .O(N__27671),
            .I(\tok.n14_adj_658_cascade_ ));
    InMux I__6675 (
            .O(N__27668),
            .I(N__27646));
    InMux I__6674 (
            .O(N__27667),
            .I(N__27646));
    InMux I__6673 (
            .O(N__27666),
            .I(N__27646));
    InMux I__6672 (
            .O(N__27665),
            .I(N__27637));
    InMux I__6671 (
            .O(N__27664),
            .I(N__27637));
    InMux I__6670 (
            .O(N__27663),
            .I(N__27637));
    InMux I__6669 (
            .O(N__27662),
            .I(N__27637));
    InMux I__6668 (
            .O(N__27661),
            .I(N__27626));
    InMux I__6667 (
            .O(N__27660),
            .I(N__27626));
    InMux I__6666 (
            .O(N__27659),
            .I(N__27626));
    InMux I__6665 (
            .O(N__27658),
            .I(N__27626));
    InMux I__6664 (
            .O(N__27657),
            .I(N__27626));
    InMux I__6663 (
            .O(N__27656),
            .I(N__27617));
    InMux I__6662 (
            .O(N__27655),
            .I(N__27617));
    InMux I__6661 (
            .O(N__27654),
            .I(N__27617));
    InMux I__6660 (
            .O(N__27653),
            .I(N__27617));
    LocalMux I__6659 (
            .O(N__27646),
            .I(N__27614));
    LocalMux I__6658 (
            .O(N__27637),
            .I(N__27607));
    LocalMux I__6657 (
            .O(N__27626),
            .I(N__27607));
    LocalMux I__6656 (
            .O(N__27617),
            .I(N__27607));
    Span4Mux_v I__6655 (
            .O(N__27614),
            .I(N__27602));
    Span4Mux_v I__6654 (
            .O(N__27607),
            .I(N__27602));
    Span4Mux_h I__6653 (
            .O(N__27602),
            .I(N__27599));
    Odrv4 I__6652 (
            .O(N__27599),
            .I(\tok.n399 ));
    CascadeMux I__6651 (
            .O(N__27596),
            .I(N__27593));
    InMux I__6650 (
            .O(N__27593),
            .I(N__27590));
    LocalMux I__6649 (
            .O(N__27590),
            .I(N__27586));
    InMux I__6648 (
            .O(N__27589),
            .I(N__27583));
    Odrv12 I__6647 (
            .O(N__27586),
            .I(\tok.n14 ));
    LocalMux I__6646 (
            .O(N__27583),
            .I(\tok.n14 ));
    CascadeMux I__6645 (
            .O(N__27578),
            .I(\tok.n4422_cascade_ ));
    InMux I__6644 (
            .O(N__27575),
            .I(N__27572));
    LocalMux I__6643 (
            .O(N__27572),
            .I(N__27567));
    InMux I__6642 (
            .O(N__27571),
            .I(N__27562));
    InMux I__6641 (
            .O(N__27570),
            .I(N__27562));
    Span4Mux_s3_v I__6640 (
            .O(N__27567),
            .I(N__27557));
    LocalMux I__6639 (
            .O(N__27562),
            .I(N__27557));
    Span4Mux_v I__6638 (
            .O(N__27557),
            .I(N__27552));
    InMux I__6637 (
            .O(N__27556),
            .I(N__27549));
    InMux I__6636 (
            .O(N__27555),
            .I(N__27546));
    Odrv4 I__6635 (
            .O(N__27552),
            .I(\tok.n11_adj_648 ));
    LocalMux I__6634 (
            .O(N__27549),
            .I(\tok.n11_adj_648 ));
    LocalMux I__6633 (
            .O(N__27546),
            .I(\tok.n11_adj_648 ));
    InMux I__6632 (
            .O(N__27539),
            .I(N__27533));
    InMux I__6631 (
            .O(N__27538),
            .I(N__27533));
    LocalMux I__6630 (
            .O(N__27533),
            .I(\tok.n4558 ));
    InMux I__6629 (
            .O(N__27530),
            .I(N__27525));
    InMux I__6628 (
            .O(N__27529),
            .I(N__27520));
    InMux I__6627 (
            .O(N__27528),
            .I(N__27520));
    LocalMux I__6626 (
            .O(N__27525),
            .I(N__27517));
    LocalMux I__6625 (
            .O(N__27520),
            .I(N__27514));
    Odrv12 I__6624 (
            .O(N__27517),
            .I(\tok.n14_adj_650 ));
    Odrv4 I__6623 (
            .O(N__27514),
            .I(\tok.n14_adj_650 ));
    CascadeMux I__6622 (
            .O(N__27509),
            .I(\tok.n51_cascade_ ));
    InMux I__6621 (
            .O(N__27506),
            .I(N__27503));
    LocalMux I__6620 (
            .O(N__27503),
            .I(\tok.n4424 ));
    InMux I__6619 (
            .O(N__27500),
            .I(N__27497));
    LocalMux I__6618 (
            .O(N__27497),
            .I(\tok.n48 ));
    InMux I__6617 (
            .O(N__27494),
            .I(N__27491));
    LocalMux I__6616 (
            .O(N__27491),
            .I(N__27488));
    Span4Mux_s3_h I__6615 (
            .O(N__27488),
            .I(N__27485));
    Sp12to4 I__6614 (
            .O(N__27485),
            .I(N__27482));
    Odrv12 I__6613 (
            .O(N__27482),
            .I(\tok.table_rd_12 ));
    InMux I__6612 (
            .O(N__27479),
            .I(N__27476));
    LocalMux I__6611 (
            .O(N__27476),
            .I(N__27473));
    Odrv12 I__6610 (
            .O(N__27473),
            .I(\tok.n5_adj_694 ));
    InMux I__6609 (
            .O(N__27470),
            .I(N__27467));
    LocalMux I__6608 (
            .O(N__27467),
            .I(N__27464));
    Span4Mux_s2_h I__6607 (
            .O(N__27464),
            .I(N__27461));
    Span4Mux_h I__6606 (
            .O(N__27461),
            .I(N__27458));
    Odrv4 I__6605 (
            .O(N__27458),
            .I(\tok.n10_adj_697 ));
    CascadeMux I__6604 (
            .O(N__27455),
            .I(\tok.n14_adj_695_cascade_ ));
    InMux I__6603 (
            .O(N__27452),
            .I(N__27449));
    LocalMux I__6602 (
            .O(N__27449),
            .I(N__27442));
    InMux I__6601 (
            .O(N__27448),
            .I(N__27439));
    InMux I__6600 (
            .O(N__27447),
            .I(N__27436));
    CascadeMux I__6599 (
            .O(N__27446),
            .I(N__27430));
    InMux I__6598 (
            .O(N__27445),
            .I(N__27424));
    Span4Mux_h I__6597 (
            .O(N__27442),
            .I(N__27418));
    LocalMux I__6596 (
            .O(N__27439),
            .I(N__27418));
    LocalMux I__6595 (
            .O(N__27436),
            .I(N__27415));
    InMux I__6594 (
            .O(N__27435),
            .I(N__27412));
    InMux I__6593 (
            .O(N__27434),
            .I(N__27408));
    InMux I__6592 (
            .O(N__27433),
            .I(N__27403));
    InMux I__6591 (
            .O(N__27430),
            .I(N__27403));
    InMux I__6590 (
            .O(N__27429),
            .I(N__27400));
    InMux I__6589 (
            .O(N__27428),
            .I(N__27396));
    InMux I__6588 (
            .O(N__27427),
            .I(N__27393));
    LocalMux I__6587 (
            .O(N__27424),
            .I(N__27389));
    InMux I__6586 (
            .O(N__27423),
            .I(N__27386));
    Span4Mux_v I__6585 (
            .O(N__27418),
            .I(N__27383));
    Span4Mux_v I__6584 (
            .O(N__27415),
            .I(N__27378));
    LocalMux I__6583 (
            .O(N__27412),
            .I(N__27378));
    InMux I__6582 (
            .O(N__27411),
            .I(N__27375));
    LocalMux I__6581 (
            .O(N__27408),
            .I(N__27370));
    LocalMux I__6580 (
            .O(N__27403),
            .I(N__27370));
    LocalMux I__6579 (
            .O(N__27400),
            .I(N__27367));
    InMux I__6578 (
            .O(N__27399),
            .I(N__27364));
    LocalMux I__6577 (
            .O(N__27396),
            .I(N__27359));
    LocalMux I__6576 (
            .O(N__27393),
            .I(N__27359));
    InMux I__6575 (
            .O(N__27392),
            .I(N__27356));
    Span12Mux_s4_v I__6574 (
            .O(N__27389),
            .I(N__27353));
    LocalMux I__6573 (
            .O(N__27386),
            .I(N__27346));
    Span4Mux_h I__6572 (
            .O(N__27383),
            .I(N__27346));
    Span4Mux_h I__6571 (
            .O(N__27378),
            .I(N__27346));
    LocalMux I__6570 (
            .O(N__27375),
            .I(N__27341));
    Span4Mux_h I__6569 (
            .O(N__27370),
            .I(N__27341));
    Sp12to4 I__6568 (
            .O(N__27367),
            .I(N__27334));
    LocalMux I__6567 (
            .O(N__27364),
            .I(N__27334));
    Span12Mux_s8_h I__6566 (
            .O(N__27359),
            .I(N__27334));
    LocalMux I__6565 (
            .O(N__27356),
            .I(\tok.A_low_4 ));
    Odrv12 I__6564 (
            .O(N__27353),
            .I(\tok.A_low_4 ));
    Odrv4 I__6563 (
            .O(N__27346),
            .I(\tok.A_low_4 ));
    Odrv4 I__6562 (
            .O(N__27341),
            .I(\tok.A_low_4 ));
    Odrv12 I__6561 (
            .O(N__27334),
            .I(\tok.A_low_4 ));
    InMux I__6560 (
            .O(N__27323),
            .I(N__27320));
    LocalMux I__6559 (
            .O(N__27320),
            .I(N__27317));
    Span4Mux_h I__6558 (
            .O(N__27317),
            .I(N__27314));
    Odrv4 I__6557 (
            .O(N__27314),
            .I(\tok.n18_adj_698 ));
    InMux I__6556 (
            .O(N__27311),
            .I(N__27307));
    InMux I__6555 (
            .O(N__27310),
            .I(N__27304));
    LocalMux I__6554 (
            .O(N__27307),
            .I(N__27299));
    LocalMux I__6553 (
            .O(N__27304),
            .I(N__27299));
    Span4Mux_v I__6552 (
            .O(N__27299),
            .I(N__27296));
    Span4Mux_h I__6551 (
            .O(N__27296),
            .I(N__27293));
    Odrv4 I__6550 (
            .O(N__27293),
            .I(\tok.n2177 ));
    InMux I__6549 (
            .O(N__27290),
            .I(N__27286));
    InMux I__6548 (
            .O(N__27289),
            .I(N__27283));
    LocalMux I__6547 (
            .O(N__27286),
            .I(\tok.n14_adj_825 ));
    LocalMux I__6546 (
            .O(N__27283),
            .I(\tok.n14_adj_825 ));
    CascadeMux I__6545 (
            .O(N__27278),
            .I(\tok.n2177_cascade_ ));
    InMux I__6544 (
            .O(N__27275),
            .I(N__27272));
    LocalMux I__6543 (
            .O(N__27272),
            .I(N__27269));
    Span4Mux_h I__6542 (
            .O(N__27269),
            .I(N__27263));
    InMux I__6541 (
            .O(N__27268),
            .I(N__27260));
    InMux I__6540 (
            .O(N__27267),
            .I(N__27257));
    InMux I__6539 (
            .O(N__27266),
            .I(N__27254));
    Odrv4 I__6538 (
            .O(N__27263),
            .I(\tok.n10_adj_646 ));
    LocalMux I__6537 (
            .O(N__27260),
            .I(\tok.n10_adj_646 ));
    LocalMux I__6536 (
            .O(N__27257),
            .I(\tok.n10_adj_646 ));
    LocalMux I__6535 (
            .O(N__27254),
            .I(\tok.n10_adj_646 ));
    InMux I__6534 (
            .O(N__27245),
            .I(N__27239));
    InMux I__6533 (
            .O(N__27244),
            .I(N__27236));
    InMux I__6532 (
            .O(N__27243),
            .I(N__27233));
    InMux I__6531 (
            .O(N__27242),
            .I(N__27229));
    LocalMux I__6530 (
            .O(N__27239),
            .I(N__27225));
    LocalMux I__6529 (
            .O(N__27236),
            .I(N__27222));
    LocalMux I__6528 (
            .O(N__27233),
            .I(N__27219));
    InMux I__6527 (
            .O(N__27232),
            .I(N__27212));
    LocalMux I__6526 (
            .O(N__27229),
            .I(N__27205));
    InMux I__6525 (
            .O(N__27228),
            .I(N__27202));
    Span4Mux_h I__6524 (
            .O(N__27225),
            .I(N__27199));
    Span4Mux_h I__6523 (
            .O(N__27222),
            .I(N__27196));
    Span4Mux_h I__6522 (
            .O(N__27219),
            .I(N__27193));
    CascadeMux I__6521 (
            .O(N__27218),
            .I(N__27189));
    InMux I__6520 (
            .O(N__27217),
            .I(N__27181));
    InMux I__6519 (
            .O(N__27216),
            .I(N__27181));
    InMux I__6518 (
            .O(N__27215),
            .I(N__27181));
    LocalMux I__6517 (
            .O(N__27212),
            .I(N__27178));
    InMux I__6516 (
            .O(N__27211),
            .I(N__27169));
    InMux I__6515 (
            .O(N__27210),
            .I(N__27169));
    InMux I__6514 (
            .O(N__27209),
            .I(N__27169));
    InMux I__6513 (
            .O(N__27208),
            .I(N__27169));
    Span4Mux_h I__6512 (
            .O(N__27205),
            .I(N__27163));
    LocalMux I__6511 (
            .O(N__27202),
            .I(N__27163));
    Span4Mux_h I__6510 (
            .O(N__27199),
            .I(N__27160));
    Span4Mux_h I__6509 (
            .O(N__27196),
            .I(N__27155));
    Span4Mux_h I__6508 (
            .O(N__27193),
            .I(N__27155));
    InMux I__6507 (
            .O(N__27192),
            .I(N__27148));
    InMux I__6506 (
            .O(N__27189),
            .I(N__27148));
    InMux I__6505 (
            .O(N__27188),
            .I(N__27148));
    LocalMux I__6504 (
            .O(N__27181),
            .I(N__27141));
    Span12Mux_s5_v I__6503 (
            .O(N__27178),
            .I(N__27141));
    LocalMux I__6502 (
            .O(N__27169),
            .I(N__27141));
    InMux I__6501 (
            .O(N__27168),
            .I(N__27138));
    Span4Mux_h I__6500 (
            .O(N__27163),
            .I(N__27135));
    Odrv4 I__6499 (
            .O(N__27160),
            .I(\tok.n132 ));
    Odrv4 I__6498 (
            .O(N__27155),
            .I(\tok.n132 ));
    LocalMux I__6497 (
            .O(N__27148),
            .I(\tok.n132 ));
    Odrv12 I__6496 (
            .O(N__27141),
            .I(\tok.n132 ));
    LocalMux I__6495 (
            .O(N__27138),
            .I(\tok.n132 ));
    Odrv4 I__6494 (
            .O(N__27135),
            .I(\tok.n132 ));
    InMux I__6493 (
            .O(N__27122),
            .I(N__27119));
    LocalMux I__6492 (
            .O(N__27119),
            .I(N__27116));
    Span12Mux_s1_h I__6491 (
            .O(N__27116),
            .I(N__27113));
    Odrv12 I__6490 (
            .O(N__27113),
            .I(\tok.table_rd_8 ));
    CascadeMux I__6489 (
            .O(N__27110),
            .I(\tok.n132_cascade_ ));
    InMux I__6488 (
            .O(N__27107),
            .I(N__27104));
    LocalMux I__6487 (
            .O(N__27104),
            .I(N__27101));
    Odrv4 I__6486 (
            .O(N__27101),
            .I(\tok.n5 ));
    InMux I__6485 (
            .O(N__27098),
            .I(N__27095));
    LocalMux I__6484 (
            .O(N__27095),
            .I(N__27092));
    Span4Mux_h I__6483 (
            .O(N__27092),
            .I(N__27089));
    Span4Mux_h I__6482 (
            .O(N__27089),
            .I(N__27086));
    Odrv4 I__6481 (
            .O(N__27086),
            .I(\tok.n10_adj_652 ));
    InMux I__6480 (
            .O(N__27083),
            .I(N__27080));
    LocalMux I__6479 (
            .O(N__27080),
            .I(N__27077));
    Odrv4 I__6478 (
            .O(N__27077),
            .I(\tok.n14_adj_651 ));
    CascadeMux I__6477 (
            .O(N__27074),
            .I(N__27068));
    CascadeMux I__6476 (
            .O(N__27073),
            .I(N__27064));
    CascadeMux I__6475 (
            .O(N__27072),
            .I(N__27058));
    CascadeMux I__6474 (
            .O(N__27071),
            .I(N__27054));
    InMux I__6473 (
            .O(N__27068),
            .I(N__27051));
    InMux I__6472 (
            .O(N__27067),
            .I(N__27047));
    InMux I__6471 (
            .O(N__27064),
            .I(N__27042));
    InMux I__6470 (
            .O(N__27063),
            .I(N__27039));
    InMux I__6469 (
            .O(N__27062),
            .I(N__27036));
    CascadeMux I__6468 (
            .O(N__27061),
            .I(N__27033));
    InMux I__6467 (
            .O(N__27058),
            .I(N__27030));
    InMux I__6466 (
            .O(N__27057),
            .I(N__27027));
    InMux I__6465 (
            .O(N__27054),
            .I(N__27024));
    LocalMux I__6464 (
            .O(N__27051),
            .I(N__27021));
    InMux I__6463 (
            .O(N__27050),
            .I(N__27018));
    LocalMux I__6462 (
            .O(N__27047),
            .I(N__27015));
    InMux I__6461 (
            .O(N__27046),
            .I(N__27012));
    InMux I__6460 (
            .O(N__27045),
            .I(N__27009));
    LocalMux I__6459 (
            .O(N__27042),
            .I(N__27006));
    LocalMux I__6458 (
            .O(N__27039),
            .I(N__27001));
    LocalMux I__6457 (
            .O(N__27036),
            .I(N__27001));
    InMux I__6456 (
            .O(N__27033),
            .I(N__26998));
    LocalMux I__6455 (
            .O(N__27030),
            .I(N__26991));
    LocalMux I__6454 (
            .O(N__27027),
            .I(N__26991));
    LocalMux I__6453 (
            .O(N__27024),
            .I(N__26991));
    Span4Mux_v I__6452 (
            .O(N__27021),
            .I(N__26988));
    LocalMux I__6451 (
            .O(N__27018),
            .I(N__26985));
    Span4Mux_v I__6450 (
            .O(N__27015),
            .I(N__26980));
    LocalMux I__6449 (
            .O(N__27012),
            .I(N__26980));
    LocalMux I__6448 (
            .O(N__27009),
            .I(N__26977));
    Span4Mux_v I__6447 (
            .O(N__27006),
            .I(N__26974));
    Span4Mux_h I__6446 (
            .O(N__27001),
            .I(N__26971));
    LocalMux I__6445 (
            .O(N__26998),
            .I(N__26968));
    Span4Mux_v I__6444 (
            .O(N__26991),
            .I(N__26963));
    Span4Mux_h I__6443 (
            .O(N__26988),
            .I(N__26963));
    Span4Mux_v I__6442 (
            .O(N__26985),
            .I(N__26958));
    Span4Mux_h I__6441 (
            .O(N__26980),
            .I(N__26958));
    Span4Mux_s3_h I__6440 (
            .O(N__26977),
            .I(N__26955));
    Odrv4 I__6439 (
            .O(N__26974),
            .I(\tok.n109 ));
    Odrv4 I__6438 (
            .O(N__26971),
            .I(\tok.n109 ));
    Odrv4 I__6437 (
            .O(N__26968),
            .I(\tok.n109 ));
    Odrv4 I__6436 (
            .O(N__26963),
            .I(\tok.n109 ));
    Odrv4 I__6435 (
            .O(N__26958),
            .I(\tok.n109 ));
    Odrv4 I__6434 (
            .O(N__26955),
            .I(\tok.n109 ));
    InMux I__6433 (
            .O(N__26942),
            .I(N__26938));
    InMux I__6432 (
            .O(N__26941),
            .I(N__26935));
    LocalMux I__6431 (
            .O(N__26938),
            .I(N__26930));
    LocalMux I__6430 (
            .O(N__26935),
            .I(N__26922));
    InMux I__6429 (
            .O(N__26934),
            .I(N__26916));
    InMux I__6428 (
            .O(N__26933),
            .I(N__26913));
    Span4Mux_v I__6427 (
            .O(N__26930),
            .I(N__26910));
    InMux I__6426 (
            .O(N__26929),
            .I(N__26907));
    InMux I__6425 (
            .O(N__26928),
            .I(N__26904));
    InMux I__6424 (
            .O(N__26927),
            .I(N__26901));
    InMux I__6423 (
            .O(N__26926),
            .I(N__26894));
    InMux I__6422 (
            .O(N__26925),
            .I(N__26894));
    Span4Mux_v I__6421 (
            .O(N__26922),
            .I(N__26891));
    InMux I__6420 (
            .O(N__26921),
            .I(N__26886));
    InMux I__6419 (
            .O(N__26920),
            .I(N__26886));
    InMux I__6418 (
            .O(N__26919),
            .I(N__26883));
    LocalMux I__6417 (
            .O(N__26916),
            .I(N__26879));
    LocalMux I__6416 (
            .O(N__26913),
            .I(N__26876));
    Span4Mux_h I__6415 (
            .O(N__26910),
            .I(N__26871));
    LocalMux I__6414 (
            .O(N__26907),
            .I(N__26871));
    LocalMux I__6413 (
            .O(N__26904),
            .I(N__26866));
    LocalMux I__6412 (
            .O(N__26901),
            .I(N__26866));
    InMux I__6411 (
            .O(N__26900),
            .I(N__26863));
    InMux I__6410 (
            .O(N__26899),
            .I(N__26860));
    LocalMux I__6409 (
            .O(N__26894),
            .I(N__26857));
    Span4Mux_h I__6408 (
            .O(N__26891),
            .I(N__26850));
    LocalMux I__6407 (
            .O(N__26886),
            .I(N__26850));
    LocalMux I__6406 (
            .O(N__26883),
            .I(N__26850));
    InMux I__6405 (
            .O(N__26882),
            .I(N__26847));
    Span4Mux_v I__6404 (
            .O(N__26879),
            .I(N__26840));
    Span4Mux_s3_h I__6403 (
            .O(N__26876),
            .I(N__26840));
    Span4Mux_v I__6402 (
            .O(N__26871),
            .I(N__26840));
    Span4Mux_h I__6401 (
            .O(N__26866),
            .I(N__26835));
    LocalMux I__6400 (
            .O(N__26863),
            .I(N__26835));
    LocalMux I__6399 (
            .O(N__26860),
            .I(N__26832));
    Odrv4 I__6398 (
            .O(N__26857),
            .I(\tok.A_low_0 ));
    Odrv4 I__6397 (
            .O(N__26850),
            .I(\tok.A_low_0 ));
    LocalMux I__6396 (
            .O(N__26847),
            .I(\tok.A_low_0 ));
    Odrv4 I__6395 (
            .O(N__26840),
            .I(\tok.A_low_0 ));
    Odrv4 I__6394 (
            .O(N__26835),
            .I(\tok.A_low_0 ));
    Odrv4 I__6393 (
            .O(N__26832),
            .I(\tok.A_low_0 ));
    CascadeMux I__6392 (
            .O(N__26819),
            .I(\tok.ram.n14_adj_631_cascade_ ));
    InMux I__6391 (
            .O(N__26816),
            .I(N__26805));
    InMux I__6390 (
            .O(N__26815),
            .I(N__26805));
    InMux I__6389 (
            .O(N__26814),
            .I(N__26800));
    InMux I__6388 (
            .O(N__26813),
            .I(N__26797));
    InMux I__6387 (
            .O(N__26812),
            .I(N__26792));
    InMux I__6386 (
            .O(N__26811),
            .I(N__26784));
    InMux I__6385 (
            .O(N__26810),
            .I(N__26784));
    LocalMux I__6384 (
            .O(N__26805),
            .I(N__26781));
    InMux I__6383 (
            .O(N__26804),
            .I(N__26776));
    InMux I__6382 (
            .O(N__26803),
            .I(N__26776));
    LocalMux I__6381 (
            .O(N__26800),
            .I(N__26773));
    LocalMux I__6380 (
            .O(N__26797),
            .I(N__26770));
    InMux I__6379 (
            .O(N__26796),
            .I(N__26765));
    InMux I__6378 (
            .O(N__26795),
            .I(N__26765));
    LocalMux I__6377 (
            .O(N__26792),
            .I(N__26762));
    InMux I__6376 (
            .O(N__26791),
            .I(N__26759));
    InMux I__6375 (
            .O(N__26790),
            .I(N__26754));
    InMux I__6374 (
            .O(N__26789),
            .I(N__26754));
    LocalMux I__6373 (
            .O(N__26784),
            .I(N__26749));
    Span4Mux_s3_v I__6372 (
            .O(N__26781),
            .I(N__26749));
    LocalMux I__6371 (
            .O(N__26776),
            .I(N__26742));
    Span4Mux_h I__6370 (
            .O(N__26773),
            .I(N__26742));
    Span4Mux_s3_v I__6369 (
            .O(N__26770),
            .I(N__26742));
    LocalMux I__6368 (
            .O(N__26765),
            .I(N__26739));
    Span4Mux_h I__6367 (
            .O(N__26762),
            .I(N__26734));
    LocalMux I__6366 (
            .O(N__26759),
            .I(N__26734));
    LocalMux I__6365 (
            .O(N__26754),
            .I(N__26731));
    Span4Mux_v I__6364 (
            .O(N__26749),
            .I(N__26727));
    Span4Mux_v I__6363 (
            .O(N__26742),
            .I(N__26724));
    Span4Mux_v I__6362 (
            .O(N__26739),
            .I(N__26717));
    Span4Mux_v I__6361 (
            .O(N__26734),
            .I(N__26717));
    Span4Mux_h I__6360 (
            .O(N__26731),
            .I(N__26717));
    InMux I__6359 (
            .O(N__26730),
            .I(N__26714));
    Sp12to4 I__6358 (
            .O(N__26727),
            .I(N__26709));
    Sp12to4 I__6357 (
            .O(N__26724),
            .I(N__26709));
    Span4Mux_h I__6356 (
            .O(N__26717),
            .I(N__26706));
    LocalMux I__6355 (
            .O(N__26714),
            .I(N__26703));
    Odrv12 I__6354 (
            .O(N__26709),
            .I(\tok.n2635 ));
    Odrv4 I__6353 (
            .O(N__26706),
            .I(\tok.n2635 ));
    Odrv4 I__6352 (
            .O(N__26703),
            .I(\tok.n2635 ));
    InMux I__6351 (
            .O(N__26696),
            .I(N__26691));
    InMux I__6350 (
            .O(N__26695),
            .I(N__26688));
    InMux I__6349 (
            .O(N__26694),
            .I(N__26685));
    LocalMux I__6348 (
            .O(N__26691),
            .I(N__26679));
    LocalMux I__6347 (
            .O(N__26688),
            .I(N__26674));
    LocalMux I__6346 (
            .O(N__26685),
            .I(N__26674));
    InMux I__6345 (
            .O(N__26684),
            .I(N__26670));
    InMux I__6344 (
            .O(N__26683),
            .I(N__26667));
    InMux I__6343 (
            .O(N__26682),
            .I(N__26664));
    Span4Mux_h I__6342 (
            .O(N__26679),
            .I(N__26659));
    Span4Mux_v I__6341 (
            .O(N__26674),
            .I(N__26659));
    InMux I__6340 (
            .O(N__26673),
            .I(N__26656));
    LocalMux I__6339 (
            .O(N__26670),
            .I(N__26651));
    LocalMux I__6338 (
            .O(N__26667),
            .I(N__26651));
    LocalMux I__6337 (
            .O(N__26664),
            .I(N__26647));
    Span4Mux_h I__6336 (
            .O(N__26659),
            .I(N__26644));
    LocalMux I__6335 (
            .O(N__26656),
            .I(N__26639));
    Span4Mux_h I__6334 (
            .O(N__26651),
            .I(N__26639));
    InMux I__6333 (
            .O(N__26650),
            .I(N__26636));
    Odrv4 I__6332 (
            .O(N__26647),
            .I(\tok.n4_adj_795 ));
    Odrv4 I__6331 (
            .O(N__26644),
            .I(\tok.n4_adj_795 ));
    Odrv4 I__6330 (
            .O(N__26639),
            .I(\tok.n4_adj_795 ));
    LocalMux I__6329 (
            .O(N__26636),
            .I(\tok.n4_adj_795 ));
    CascadeMux I__6328 (
            .O(N__26627),
            .I(\tok.n41_cascade_ ));
    CascadeMux I__6327 (
            .O(N__26624),
            .I(N__26619));
    InMux I__6326 (
            .O(N__26623),
            .I(N__26610));
    InMux I__6325 (
            .O(N__26622),
            .I(N__26610));
    InMux I__6324 (
            .O(N__26619),
            .I(N__26605));
    InMux I__6323 (
            .O(N__26618),
            .I(N__26605));
    InMux I__6322 (
            .O(N__26617),
            .I(N__26592));
    InMux I__6321 (
            .O(N__26616),
            .I(N__26592));
    InMux I__6320 (
            .O(N__26615),
            .I(N__26589));
    LocalMux I__6319 (
            .O(N__26610),
            .I(N__26584));
    LocalMux I__6318 (
            .O(N__26605),
            .I(N__26584));
    InMux I__6317 (
            .O(N__26604),
            .I(N__26581));
    InMux I__6316 (
            .O(N__26603),
            .I(N__26578));
    InMux I__6315 (
            .O(N__26602),
            .I(N__26573));
    InMux I__6314 (
            .O(N__26601),
            .I(N__26573));
    InMux I__6313 (
            .O(N__26600),
            .I(N__26570));
    InMux I__6312 (
            .O(N__26599),
            .I(N__26567));
    InMux I__6311 (
            .O(N__26598),
            .I(N__26564));
    CascadeMux I__6310 (
            .O(N__26597),
            .I(N__26559));
    LocalMux I__6309 (
            .O(N__26592),
            .I(N__26554));
    LocalMux I__6308 (
            .O(N__26589),
            .I(N__26554));
    Span4Mux_h I__6307 (
            .O(N__26584),
            .I(N__26549));
    LocalMux I__6306 (
            .O(N__26581),
            .I(N__26549));
    LocalMux I__6305 (
            .O(N__26578),
            .I(N__26544));
    LocalMux I__6304 (
            .O(N__26573),
            .I(N__26544));
    LocalMux I__6303 (
            .O(N__26570),
            .I(N__26539));
    LocalMux I__6302 (
            .O(N__26567),
            .I(N__26539));
    LocalMux I__6301 (
            .O(N__26564),
            .I(N__26536));
    InMux I__6300 (
            .O(N__26563),
            .I(N__26529));
    InMux I__6299 (
            .O(N__26562),
            .I(N__26529));
    InMux I__6298 (
            .O(N__26559),
            .I(N__26529));
    Span4Mux_v I__6297 (
            .O(N__26554),
            .I(N__26526));
    Span4Mux_v I__6296 (
            .O(N__26549),
            .I(N__26521));
    Span4Mux_v I__6295 (
            .O(N__26544),
            .I(N__26521));
    Span4Mux_s3_v I__6294 (
            .O(N__26539),
            .I(N__26514));
    Span4Mux_h I__6293 (
            .O(N__26536),
            .I(N__26514));
    LocalMux I__6292 (
            .O(N__26529),
            .I(N__26514));
    Sp12to4 I__6291 (
            .O(N__26526),
            .I(N__26511));
    Span4Mux_h I__6290 (
            .O(N__26521),
            .I(N__26508));
    Span4Mux_v I__6289 (
            .O(N__26514),
            .I(N__26505));
    Odrv12 I__6288 (
            .O(N__26511),
            .I(\tok.n884 ));
    Odrv4 I__6287 (
            .O(N__26508),
            .I(\tok.n884 ));
    Odrv4 I__6286 (
            .O(N__26505),
            .I(\tok.n884 ));
    InMux I__6285 (
            .O(N__26498),
            .I(N__26494));
    InMux I__6284 (
            .O(N__26497),
            .I(N__26491));
    LocalMux I__6283 (
            .O(N__26494),
            .I(\tok.n14_adj_702 ));
    LocalMux I__6282 (
            .O(N__26491),
            .I(\tok.n14_adj_702 ));
    InMux I__6281 (
            .O(N__26486),
            .I(N__26482));
    InMux I__6280 (
            .O(N__26485),
            .I(N__26479));
    LocalMux I__6279 (
            .O(N__26482),
            .I(N__26476));
    LocalMux I__6278 (
            .O(N__26479),
            .I(N__26473));
    Span4Mux_h I__6277 (
            .O(N__26476),
            .I(N__26470));
    Span4Mux_v I__6276 (
            .O(N__26473),
            .I(N__26467));
    Span4Mux_h I__6275 (
            .O(N__26470),
            .I(N__26464));
    Span4Mux_h I__6274 (
            .O(N__26467),
            .I(N__26461));
    Odrv4 I__6273 (
            .O(N__26464),
            .I(\tok.n15_adj_662 ));
    Odrv4 I__6272 (
            .O(N__26461),
            .I(\tok.n15_adj_662 ));
    CascadeMux I__6271 (
            .O(N__26456),
            .I(N__26452));
    InMux I__6270 (
            .O(N__26455),
            .I(N__26449));
    InMux I__6269 (
            .O(N__26452),
            .I(N__26446));
    LocalMux I__6268 (
            .O(N__26449),
            .I(\tok.n4464 ));
    LocalMux I__6267 (
            .O(N__26446),
            .I(\tok.n4464 ));
    InMux I__6266 (
            .O(N__26441),
            .I(N__26438));
    LocalMux I__6265 (
            .O(N__26438),
            .I(\tok.n4573 ));
    InMux I__6264 (
            .O(N__26435),
            .I(N__26431));
    CascadeMux I__6263 (
            .O(N__26434),
            .I(N__26428));
    LocalMux I__6262 (
            .O(N__26431),
            .I(N__26425));
    InMux I__6261 (
            .O(N__26428),
            .I(N__26422));
    Odrv12 I__6260 (
            .O(N__26425),
            .I(\tok.n9_adj_645 ));
    LocalMux I__6259 (
            .O(N__26422),
            .I(\tok.n9_adj_645 ));
    InMux I__6258 (
            .O(N__26417),
            .I(N__26411));
    InMux I__6257 (
            .O(N__26416),
            .I(N__26411));
    LocalMux I__6256 (
            .O(N__26411),
            .I(N__26407));
    InMux I__6255 (
            .O(N__26410),
            .I(N__26404));
    Span4Mux_h I__6254 (
            .O(N__26407),
            .I(N__26401));
    LocalMux I__6253 (
            .O(N__26404),
            .I(N__26398));
    Span4Mux_h I__6252 (
            .O(N__26401),
            .I(N__26394));
    Span4Mux_v I__6251 (
            .O(N__26398),
            .I(N__26391));
    InMux I__6250 (
            .O(N__26397),
            .I(N__26388));
    Odrv4 I__6249 (
            .O(N__26394),
            .I(\tok.n11 ));
    Odrv4 I__6248 (
            .O(N__26391),
            .I(\tok.n11 ));
    LocalMux I__6247 (
            .O(N__26388),
            .I(\tok.n11 ));
    CascadeMux I__6246 (
            .O(N__26381),
            .I(\tok.n6_cascade_ ));
    InMux I__6245 (
            .O(N__26378),
            .I(N__26375));
    LocalMux I__6244 (
            .O(N__26375),
            .I(N__26371));
    InMux I__6243 (
            .O(N__26374),
            .I(N__26368));
    Odrv12 I__6242 (
            .O(N__26371),
            .I(\tok.C_stk.tail_2 ));
    LocalMux I__6241 (
            .O(N__26368),
            .I(\tok.C_stk.tail_2 ));
    CascadeMux I__6240 (
            .O(N__26363),
            .I(\tok.C_stk.n4876_cascade_ ));
    InMux I__6239 (
            .O(N__26360),
            .I(N__26353));
    InMux I__6238 (
            .O(N__26359),
            .I(N__26353));
    CascadeMux I__6237 (
            .O(N__26358),
            .I(N__26349));
    LocalMux I__6236 (
            .O(N__26353),
            .I(N__26342));
    InMux I__6235 (
            .O(N__26352),
            .I(N__26337));
    InMux I__6234 (
            .O(N__26349),
            .I(N__26337));
    InMux I__6233 (
            .O(N__26348),
            .I(N__26332));
    InMux I__6232 (
            .O(N__26347),
            .I(N__26332));
    InMux I__6231 (
            .O(N__26346),
            .I(N__26325));
    InMux I__6230 (
            .O(N__26345),
            .I(N__26325));
    Span4Mux_s3_v I__6229 (
            .O(N__26342),
            .I(N__26317));
    LocalMux I__6228 (
            .O(N__26337),
            .I(N__26317));
    LocalMux I__6227 (
            .O(N__26332),
            .I(N__26314));
    InMux I__6226 (
            .O(N__26331),
            .I(N__26309));
    InMux I__6225 (
            .O(N__26330),
            .I(N__26309));
    LocalMux I__6224 (
            .O(N__26325),
            .I(N__26306));
    InMux I__6223 (
            .O(N__26324),
            .I(N__26296));
    InMux I__6222 (
            .O(N__26323),
            .I(N__26296));
    InMux I__6221 (
            .O(N__26322),
            .I(N__26296));
    Span4Mux_v I__6220 (
            .O(N__26317),
            .I(N__26291));
    Span4Mux_s3_v I__6219 (
            .O(N__26314),
            .I(N__26291));
    LocalMux I__6218 (
            .O(N__26309),
            .I(N__26286));
    Span4Mux_h I__6217 (
            .O(N__26306),
            .I(N__26286));
    InMux I__6216 (
            .O(N__26305),
            .I(N__26279));
    InMux I__6215 (
            .O(N__26304),
            .I(N__26279));
    InMux I__6214 (
            .O(N__26303),
            .I(N__26279));
    LocalMux I__6213 (
            .O(N__26296),
            .I(\tok.C_stk.n600 ));
    Odrv4 I__6212 (
            .O(N__26291),
            .I(\tok.C_stk.n600 ));
    Odrv4 I__6211 (
            .O(N__26286),
            .I(\tok.C_stk.n600 ));
    LocalMux I__6210 (
            .O(N__26279),
            .I(\tok.C_stk.n600 ));
    ClkMux I__6209 (
            .O(N__26270),
            .I(N__26042));
    ClkMux I__6208 (
            .O(N__26269),
            .I(N__26042));
    ClkMux I__6207 (
            .O(N__26268),
            .I(N__26042));
    ClkMux I__6206 (
            .O(N__26267),
            .I(N__26042));
    ClkMux I__6205 (
            .O(N__26266),
            .I(N__26042));
    ClkMux I__6204 (
            .O(N__26265),
            .I(N__26042));
    ClkMux I__6203 (
            .O(N__26264),
            .I(N__26042));
    ClkMux I__6202 (
            .O(N__26263),
            .I(N__26042));
    ClkMux I__6201 (
            .O(N__26262),
            .I(N__26042));
    ClkMux I__6200 (
            .O(N__26261),
            .I(N__26042));
    ClkMux I__6199 (
            .O(N__26260),
            .I(N__26042));
    ClkMux I__6198 (
            .O(N__26259),
            .I(N__26042));
    ClkMux I__6197 (
            .O(N__26258),
            .I(N__26042));
    ClkMux I__6196 (
            .O(N__26257),
            .I(N__26042));
    ClkMux I__6195 (
            .O(N__26256),
            .I(N__26042));
    ClkMux I__6194 (
            .O(N__26255),
            .I(N__26042));
    ClkMux I__6193 (
            .O(N__26254),
            .I(N__26042));
    ClkMux I__6192 (
            .O(N__26253),
            .I(N__26042));
    ClkMux I__6191 (
            .O(N__26252),
            .I(N__26042));
    ClkMux I__6190 (
            .O(N__26251),
            .I(N__26042));
    ClkMux I__6189 (
            .O(N__26250),
            .I(N__26042));
    ClkMux I__6188 (
            .O(N__26249),
            .I(N__26042));
    ClkMux I__6187 (
            .O(N__26248),
            .I(N__26042));
    ClkMux I__6186 (
            .O(N__26247),
            .I(N__26042));
    ClkMux I__6185 (
            .O(N__26246),
            .I(N__26042));
    ClkMux I__6184 (
            .O(N__26245),
            .I(N__26042));
    ClkMux I__6183 (
            .O(N__26244),
            .I(N__26042));
    ClkMux I__6182 (
            .O(N__26243),
            .I(N__26042));
    ClkMux I__6181 (
            .O(N__26242),
            .I(N__26042));
    ClkMux I__6180 (
            .O(N__26241),
            .I(N__26042));
    ClkMux I__6179 (
            .O(N__26240),
            .I(N__26042));
    ClkMux I__6178 (
            .O(N__26239),
            .I(N__26042));
    ClkMux I__6177 (
            .O(N__26238),
            .I(N__26042));
    ClkMux I__6176 (
            .O(N__26237),
            .I(N__26042));
    ClkMux I__6175 (
            .O(N__26236),
            .I(N__26042));
    ClkMux I__6174 (
            .O(N__26235),
            .I(N__26042));
    ClkMux I__6173 (
            .O(N__26234),
            .I(N__26042));
    ClkMux I__6172 (
            .O(N__26233),
            .I(N__26042));
    ClkMux I__6171 (
            .O(N__26232),
            .I(N__26042));
    ClkMux I__6170 (
            .O(N__26231),
            .I(N__26042));
    ClkMux I__6169 (
            .O(N__26230),
            .I(N__26042));
    ClkMux I__6168 (
            .O(N__26229),
            .I(N__26042));
    ClkMux I__6167 (
            .O(N__26228),
            .I(N__26042));
    ClkMux I__6166 (
            .O(N__26227),
            .I(N__26042));
    ClkMux I__6165 (
            .O(N__26226),
            .I(N__26042));
    ClkMux I__6164 (
            .O(N__26225),
            .I(N__26042));
    ClkMux I__6163 (
            .O(N__26224),
            .I(N__26042));
    ClkMux I__6162 (
            .O(N__26223),
            .I(N__26042));
    ClkMux I__6161 (
            .O(N__26222),
            .I(N__26042));
    ClkMux I__6160 (
            .O(N__26221),
            .I(N__26042));
    ClkMux I__6159 (
            .O(N__26220),
            .I(N__26042));
    ClkMux I__6158 (
            .O(N__26219),
            .I(N__26042));
    ClkMux I__6157 (
            .O(N__26218),
            .I(N__26042));
    ClkMux I__6156 (
            .O(N__26217),
            .I(N__26042));
    ClkMux I__6155 (
            .O(N__26216),
            .I(N__26042));
    ClkMux I__6154 (
            .O(N__26215),
            .I(N__26042));
    ClkMux I__6153 (
            .O(N__26214),
            .I(N__26042));
    ClkMux I__6152 (
            .O(N__26213),
            .I(N__26042));
    ClkMux I__6151 (
            .O(N__26212),
            .I(N__26042));
    ClkMux I__6150 (
            .O(N__26211),
            .I(N__26042));
    ClkMux I__6149 (
            .O(N__26210),
            .I(N__26042));
    ClkMux I__6148 (
            .O(N__26209),
            .I(N__26042));
    ClkMux I__6147 (
            .O(N__26208),
            .I(N__26042));
    ClkMux I__6146 (
            .O(N__26207),
            .I(N__26042));
    ClkMux I__6145 (
            .O(N__26206),
            .I(N__26042));
    ClkMux I__6144 (
            .O(N__26205),
            .I(N__26042));
    ClkMux I__6143 (
            .O(N__26204),
            .I(N__26042));
    ClkMux I__6142 (
            .O(N__26203),
            .I(N__26042));
    ClkMux I__6141 (
            .O(N__26202),
            .I(N__26042));
    ClkMux I__6140 (
            .O(N__26201),
            .I(N__26042));
    ClkMux I__6139 (
            .O(N__26200),
            .I(N__26042));
    ClkMux I__6138 (
            .O(N__26199),
            .I(N__26042));
    ClkMux I__6137 (
            .O(N__26198),
            .I(N__26042));
    ClkMux I__6136 (
            .O(N__26197),
            .I(N__26042));
    ClkMux I__6135 (
            .O(N__26196),
            .I(N__26042));
    ClkMux I__6134 (
            .O(N__26195),
            .I(N__26042));
    GlobalMux I__6133 (
            .O(N__26042),
            .I(N__26039));
    DummyBuf I__6132 (
            .O(N__26039),
            .I(clk));
    CascadeMux I__6131 (
            .O(N__26036),
            .I(N__26033));
    InMux I__6130 (
            .O(N__26033),
            .I(N__26027));
    InMux I__6129 (
            .O(N__26032),
            .I(N__26024));
    InMux I__6128 (
            .O(N__26031),
            .I(N__26019));
    InMux I__6127 (
            .O(N__26030),
            .I(N__26019));
    LocalMux I__6126 (
            .O(N__26027),
            .I(N__26016));
    LocalMux I__6125 (
            .O(N__26024),
            .I(N__26011));
    LocalMux I__6124 (
            .O(N__26019),
            .I(N__26011));
    Span4Mux_v I__6123 (
            .O(N__26016),
            .I(N__26008));
    Span4Mux_s3_h I__6122 (
            .O(N__26011),
            .I(N__26005));
    Odrv4 I__6121 (
            .O(N__26008),
            .I(\tok.tc_plus_1_2 ));
    Odrv4 I__6120 (
            .O(N__26005),
            .I(\tok.tc_plus_1_2 ));
    InMux I__6119 (
            .O(N__26000),
            .I(N__25997));
    LocalMux I__6118 (
            .O(N__25997),
            .I(N__25991));
    InMux I__6117 (
            .O(N__25996),
            .I(N__25987));
    InMux I__6116 (
            .O(N__25995),
            .I(N__25984));
    InMux I__6115 (
            .O(N__25994),
            .I(N__25980));
    Span4Mux_v I__6114 (
            .O(N__25991),
            .I(N__25975));
    InMux I__6113 (
            .O(N__25990),
            .I(N__25972));
    LocalMux I__6112 (
            .O(N__25987),
            .I(N__25969));
    LocalMux I__6111 (
            .O(N__25984),
            .I(N__25966));
    InMux I__6110 (
            .O(N__25983),
            .I(N__25963));
    LocalMux I__6109 (
            .O(N__25980),
            .I(N__25960));
    InMux I__6108 (
            .O(N__25979),
            .I(N__25957));
    InMux I__6107 (
            .O(N__25978),
            .I(N__25954));
    Span4Mux_h I__6106 (
            .O(N__25975),
            .I(N__25949));
    LocalMux I__6105 (
            .O(N__25972),
            .I(N__25949));
    Span4Mux_h I__6104 (
            .O(N__25969),
            .I(N__25946));
    Span4Mux_h I__6103 (
            .O(N__25966),
            .I(N__25943));
    LocalMux I__6102 (
            .O(N__25963),
            .I(N__25938));
    Span4Mux_v I__6101 (
            .O(N__25960),
            .I(N__25938));
    LocalMux I__6100 (
            .O(N__25957),
            .I(N__25933));
    LocalMux I__6099 (
            .O(N__25954),
            .I(N__25933));
    Odrv4 I__6098 (
            .O(N__25949),
            .I(\tok.tc__7__N_134 ));
    Odrv4 I__6097 (
            .O(N__25946),
            .I(\tok.tc__7__N_134 ));
    Odrv4 I__6096 (
            .O(N__25943),
            .I(\tok.tc__7__N_134 ));
    Odrv4 I__6095 (
            .O(N__25938),
            .I(\tok.tc__7__N_134 ));
    Odrv12 I__6094 (
            .O(N__25933),
            .I(\tok.tc__7__N_134 ));
    CascadeMux I__6093 (
            .O(N__25922),
            .I(\tok.ram.n4711_cascade_ ));
    CascadeMux I__6092 (
            .O(N__25919),
            .I(\tok.n1_adj_724_cascade_ ));
    InMux I__6091 (
            .O(N__25916),
            .I(N__25913));
    LocalMux I__6090 (
            .O(N__25913),
            .I(\tok.n13_adj_725 ));
    InMux I__6089 (
            .O(N__25910),
            .I(N__25905));
    InMux I__6088 (
            .O(N__25909),
            .I(N__25900));
    InMux I__6087 (
            .O(N__25908),
            .I(N__25900));
    LocalMux I__6086 (
            .O(N__25905),
            .I(N__25894));
    LocalMux I__6085 (
            .O(N__25900),
            .I(N__25891));
    InMux I__6084 (
            .O(N__25899),
            .I(N__25888));
    InMux I__6083 (
            .O(N__25898),
            .I(N__25885));
    InMux I__6082 (
            .O(N__25897),
            .I(N__25881));
    Span4Mux_s1_h I__6081 (
            .O(N__25894),
            .I(N__25874));
    Span4Mux_v I__6080 (
            .O(N__25891),
            .I(N__25874));
    LocalMux I__6079 (
            .O(N__25888),
            .I(N__25874));
    LocalMux I__6078 (
            .O(N__25885),
            .I(N__25869));
    InMux I__6077 (
            .O(N__25884),
            .I(N__25866));
    LocalMux I__6076 (
            .O(N__25881),
            .I(N__25861));
    Span4Mux_h I__6075 (
            .O(N__25874),
            .I(N__25861));
    InMux I__6074 (
            .O(N__25873),
            .I(N__25858));
    InMux I__6073 (
            .O(N__25872),
            .I(N__25855));
    Odrv4 I__6072 (
            .O(N__25869),
            .I(\tok.n101_adj_776 ));
    LocalMux I__6071 (
            .O(N__25866),
            .I(\tok.n101_adj_776 ));
    Odrv4 I__6070 (
            .O(N__25861),
            .I(\tok.n101_adj_776 ));
    LocalMux I__6069 (
            .O(N__25858),
            .I(\tok.n101_adj_776 ));
    LocalMux I__6068 (
            .O(N__25855),
            .I(\tok.n101_adj_776 ));
    InMux I__6067 (
            .O(N__25844),
            .I(N__25841));
    LocalMux I__6066 (
            .O(N__25841),
            .I(\tok.ram.n4708 ));
    InMux I__6065 (
            .O(N__25838),
            .I(N__25835));
    LocalMux I__6064 (
            .O(N__25835),
            .I(\tok.n1_adj_736 ));
    InMux I__6063 (
            .O(N__25832),
            .I(N__25829));
    LocalMux I__6062 (
            .O(N__25829),
            .I(\tok.n5_adj_737 ));
    InMux I__6061 (
            .O(N__25826),
            .I(N__25822));
    CascadeMux I__6060 (
            .O(N__25825),
            .I(N__25817));
    LocalMux I__6059 (
            .O(N__25822),
            .I(N__25813));
    InMux I__6058 (
            .O(N__25821),
            .I(N__25806));
    InMux I__6057 (
            .O(N__25820),
            .I(N__25806));
    InMux I__6056 (
            .O(N__25817),
            .I(N__25806));
    InMux I__6055 (
            .O(N__25816),
            .I(N__25803));
    Odrv4 I__6054 (
            .O(N__25813),
            .I(\tok.c_stk_r_2 ));
    LocalMux I__6053 (
            .O(N__25806),
            .I(\tok.c_stk_r_2 ));
    LocalMux I__6052 (
            .O(N__25803),
            .I(\tok.c_stk_r_2 ));
    CascadeMux I__6051 (
            .O(N__25796),
            .I(N__25793));
    InMux I__6050 (
            .O(N__25793),
            .I(N__25789));
    InMux I__6049 (
            .O(N__25792),
            .I(N__25786));
    LocalMux I__6048 (
            .O(N__25789),
            .I(N__25783));
    LocalMux I__6047 (
            .O(N__25786),
            .I(N__25780));
    Span4Mux_v I__6046 (
            .O(N__25783),
            .I(N__25777));
    Span4Mux_v I__6045 (
            .O(N__25780),
            .I(N__25774));
    Span4Mux_h I__6044 (
            .O(N__25777),
            .I(N__25771));
    Span4Mux_h I__6043 (
            .O(N__25774),
            .I(N__25768));
    Span4Mux_h I__6042 (
            .O(N__25771),
            .I(N__25765));
    Odrv4 I__6041 (
            .O(N__25768),
            .I(\tok.table_rd_2 ));
    Odrv4 I__6040 (
            .O(N__25765),
            .I(\tok.table_rd_2 ));
    CascadeMux I__6039 (
            .O(N__25760),
            .I(\tok.n83_adj_721_cascade_ ));
    InMux I__6038 (
            .O(N__25757),
            .I(N__25754));
    LocalMux I__6037 (
            .O(N__25754),
            .I(\tok.n4692 ));
    InMux I__6036 (
            .O(N__25751),
            .I(N__25748));
    LocalMux I__6035 (
            .O(N__25748),
            .I(N__25744));
    InMux I__6034 (
            .O(N__25747),
            .I(N__25741));
    Span4Mux_s2_v I__6033 (
            .O(N__25744),
            .I(N__25738));
    LocalMux I__6032 (
            .O(N__25741),
            .I(\tok.tail_10 ));
    Odrv4 I__6031 (
            .O(N__25738),
            .I(\tok.tail_10 ));
    CascadeMux I__6030 (
            .O(N__25733),
            .I(N__25701));
    CascadeMux I__6029 (
            .O(N__25732),
            .I(N__25698));
    InMux I__6028 (
            .O(N__25731),
            .I(N__25678));
    InMux I__6027 (
            .O(N__25730),
            .I(N__25678));
    InMux I__6026 (
            .O(N__25729),
            .I(N__25678));
    InMux I__6025 (
            .O(N__25728),
            .I(N__25678));
    InMux I__6024 (
            .O(N__25727),
            .I(N__25678));
    InMux I__6023 (
            .O(N__25726),
            .I(N__25678));
    InMux I__6022 (
            .O(N__25725),
            .I(N__25678));
    InMux I__6021 (
            .O(N__25724),
            .I(N__25678));
    InMux I__6020 (
            .O(N__25723),
            .I(N__25661));
    InMux I__6019 (
            .O(N__25722),
            .I(N__25661));
    InMux I__6018 (
            .O(N__25721),
            .I(N__25661));
    InMux I__6017 (
            .O(N__25720),
            .I(N__25661));
    InMux I__6016 (
            .O(N__25719),
            .I(N__25661));
    InMux I__6015 (
            .O(N__25718),
            .I(N__25661));
    InMux I__6014 (
            .O(N__25717),
            .I(N__25661));
    InMux I__6013 (
            .O(N__25716),
            .I(N__25661));
    InMux I__6012 (
            .O(N__25715),
            .I(N__25643));
    InMux I__6011 (
            .O(N__25714),
            .I(N__25643));
    InMux I__6010 (
            .O(N__25713),
            .I(N__25643));
    InMux I__6009 (
            .O(N__25712),
            .I(N__25643));
    InMux I__6008 (
            .O(N__25711),
            .I(N__25643));
    InMux I__6007 (
            .O(N__25710),
            .I(N__25643));
    InMux I__6006 (
            .O(N__25709),
            .I(N__25643));
    InMux I__6005 (
            .O(N__25708),
            .I(N__25643));
    CascadeMux I__6004 (
            .O(N__25707),
            .I(N__25632));
    CascadeMux I__6003 (
            .O(N__25706),
            .I(N__25629));
    CascadeMux I__6002 (
            .O(N__25705),
            .I(N__25626));
    CascadeMux I__6001 (
            .O(N__25704),
            .I(N__25623));
    InMux I__6000 (
            .O(N__25701),
            .I(N__25608));
    InMux I__5999 (
            .O(N__25698),
            .I(N__25608));
    InMux I__5998 (
            .O(N__25697),
            .I(N__25608));
    InMux I__5997 (
            .O(N__25696),
            .I(N__25608));
    InMux I__5996 (
            .O(N__25695),
            .I(N__25608));
    LocalMux I__5995 (
            .O(N__25678),
            .I(N__25605));
    LocalMux I__5994 (
            .O(N__25661),
            .I(N__25602));
    CascadeMux I__5993 (
            .O(N__25660),
            .I(N__25599));
    LocalMux I__5992 (
            .O(N__25643),
            .I(N__25578));
    InMux I__5991 (
            .O(N__25642),
            .I(N__25561));
    InMux I__5990 (
            .O(N__25641),
            .I(N__25561));
    InMux I__5989 (
            .O(N__25640),
            .I(N__25561));
    InMux I__5988 (
            .O(N__25639),
            .I(N__25561));
    InMux I__5987 (
            .O(N__25638),
            .I(N__25561));
    InMux I__5986 (
            .O(N__25637),
            .I(N__25561));
    InMux I__5985 (
            .O(N__25636),
            .I(N__25561));
    InMux I__5984 (
            .O(N__25635),
            .I(N__25561));
    InMux I__5983 (
            .O(N__25632),
            .I(N__25544));
    InMux I__5982 (
            .O(N__25629),
            .I(N__25544));
    InMux I__5981 (
            .O(N__25626),
            .I(N__25544));
    InMux I__5980 (
            .O(N__25623),
            .I(N__25544));
    InMux I__5979 (
            .O(N__25622),
            .I(N__25544));
    InMux I__5978 (
            .O(N__25621),
            .I(N__25544));
    InMux I__5977 (
            .O(N__25620),
            .I(N__25544));
    InMux I__5976 (
            .O(N__25619),
            .I(N__25544));
    LocalMux I__5975 (
            .O(N__25608),
            .I(N__25537));
    Span4Mux_s3_v I__5974 (
            .O(N__25605),
            .I(N__25537));
    Span4Mux_s1_h I__5973 (
            .O(N__25602),
            .I(N__25537));
    InMux I__5972 (
            .O(N__25599),
            .I(N__25530));
    InMux I__5971 (
            .O(N__25598),
            .I(N__25530));
    InMux I__5970 (
            .O(N__25597),
            .I(N__25530));
    InMux I__5969 (
            .O(N__25596),
            .I(N__25513));
    InMux I__5968 (
            .O(N__25595),
            .I(N__25513));
    InMux I__5967 (
            .O(N__25594),
            .I(N__25513));
    InMux I__5966 (
            .O(N__25593),
            .I(N__25513));
    InMux I__5965 (
            .O(N__25592),
            .I(N__25513));
    InMux I__5964 (
            .O(N__25591),
            .I(N__25513));
    InMux I__5963 (
            .O(N__25590),
            .I(N__25513));
    InMux I__5962 (
            .O(N__25589),
            .I(N__25513));
    InMux I__5961 (
            .O(N__25588),
            .I(N__25496));
    InMux I__5960 (
            .O(N__25587),
            .I(N__25496));
    InMux I__5959 (
            .O(N__25586),
            .I(N__25496));
    InMux I__5958 (
            .O(N__25585),
            .I(N__25496));
    InMux I__5957 (
            .O(N__25584),
            .I(N__25496));
    InMux I__5956 (
            .O(N__25583),
            .I(N__25496));
    InMux I__5955 (
            .O(N__25582),
            .I(N__25496));
    InMux I__5954 (
            .O(N__25581),
            .I(N__25496));
    Span4Mux_s2_v I__5953 (
            .O(N__25578),
            .I(N__25493));
    LocalMux I__5952 (
            .O(N__25561),
            .I(N__25488));
    LocalMux I__5951 (
            .O(N__25544),
            .I(N__25488));
    Span4Mux_h I__5950 (
            .O(N__25537),
            .I(N__25485));
    LocalMux I__5949 (
            .O(N__25530),
            .I(\tok.C_stk_delta_1 ));
    LocalMux I__5948 (
            .O(N__25513),
            .I(\tok.C_stk_delta_1 ));
    LocalMux I__5947 (
            .O(N__25496),
            .I(\tok.C_stk_delta_1 ));
    Odrv4 I__5946 (
            .O(N__25493),
            .I(\tok.C_stk_delta_1 ));
    Odrv12 I__5945 (
            .O(N__25488),
            .I(\tok.C_stk_delta_1 ));
    Odrv4 I__5944 (
            .O(N__25485),
            .I(\tok.C_stk_delta_1 ));
    CEMux I__5943 (
            .O(N__25472),
            .I(N__25468));
    CEMux I__5942 (
            .O(N__25471),
            .I(N__25455));
    LocalMux I__5941 (
            .O(N__25468),
            .I(N__25452));
    CEMux I__5940 (
            .O(N__25467),
            .I(N__25449));
    CEMux I__5939 (
            .O(N__25466),
            .I(N__25446));
    CEMux I__5938 (
            .O(N__25465),
            .I(N__25443));
    InMux I__5937 (
            .O(N__25464),
            .I(N__25428));
    InMux I__5936 (
            .O(N__25463),
            .I(N__25428));
    InMux I__5935 (
            .O(N__25462),
            .I(N__25428));
    InMux I__5934 (
            .O(N__25461),
            .I(N__25428));
    InMux I__5933 (
            .O(N__25460),
            .I(N__25428));
    InMux I__5932 (
            .O(N__25459),
            .I(N__25428));
    InMux I__5931 (
            .O(N__25458),
            .I(N__25428));
    LocalMux I__5930 (
            .O(N__25455),
            .I(N__25423));
    Span4Mux_s2_h I__5929 (
            .O(N__25452),
            .I(N__25417));
    LocalMux I__5928 (
            .O(N__25449),
            .I(N__25414));
    LocalMux I__5927 (
            .O(N__25446),
            .I(N__25411));
    LocalMux I__5926 (
            .O(N__25443),
            .I(N__25408));
    LocalMux I__5925 (
            .O(N__25428),
            .I(N__25405));
    CEMux I__5924 (
            .O(N__25427),
            .I(N__25402));
    CEMux I__5923 (
            .O(N__25426),
            .I(N__25399));
    Span4Mux_h I__5922 (
            .O(N__25423),
            .I(N__25396));
    InMux I__5921 (
            .O(N__25422),
            .I(N__25389));
    InMux I__5920 (
            .O(N__25421),
            .I(N__25389));
    InMux I__5919 (
            .O(N__25420),
            .I(N__25389));
    Span4Mux_h I__5918 (
            .O(N__25417),
            .I(N__25386));
    Span4Mux_s2_h I__5917 (
            .O(N__25414),
            .I(N__25377));
    Span4Mux_s2_h I__5916 (
            .O(N__25411),
            .I(N__25377));
    Span4Mux_s2_v I__5915 (
            .O(N__25408),
            .I(N__25377));
    Span4Mux_v I__5914 (
            .O(N__25405),
            .I(N__25377));
    LocalMux I__5913 (
            .O(N__25402),
            .I(\tok.rd_7__N_374 ));
    LocalMux I__5912 (
            .O(N__25399),
            .I(\tok.rd_7__N_374 ));
    Odrv4 I__5911 (
            .O(N__25396),
            .I(\tok.rd_7__N_374 ));
    LocalMux I__5910 (
            .O(N__25389),
            .I(\tok.rd_7__N_374 ));
    Odrv4 I__5909 (
            .O(N__25386),
            .I(\tok.rd_7__N_374 ));
    Odrv4 I__5908 (
            .O(N__25377),
            .I(\tok.rd_7__N_374 ));
    InMux I__5907 (
            .O(N__25364),
            .I(N__25360));
    InMux I__5906 (
            .O(N__25363),
            .I(N__25356));
    LocalMux I__5905 (
            .O(N__25360),
            .I(N__25353));
    InMux I__5904 (
            .O(N__25359),
            .I(N__25349));
    LocalMux I__5903 (
            .O(N__25356),
            .I(N__25344));
    Span4Mux_v I__5902 (
            .O(N__25353),
            .I(N__25344));
    InMux I__5901 (
            .O(N__25352),
            .I(N__25341));
    LocalMux I__5900 (
            .O(N__25349),
            .I(c_stk_w_7_N_18_4));
    Odrv4 I__5899 (
            .O(N__25344),
            .I(c_stk_w_7_N_18_4));
    LocalMux I__5898 (
            .O(N__25341),
            .I(c_stk_w_7_N_18_4));
    InMux I__5897 (
            .O(N__25334),
            .I(N__25331));
    LocalMux I__5896 (
            .O(N__25331),
            .I(N__25328));
    Span12Mux_v I__5895 (
            .O(N__25328),
            .I(N__25324));
    InMux I__5894 (
            .O(N__25327),
            .I(N__25321));
    Odrv12 I__5893 (
            .O(N__25324),
            .I(\tok.C_stk.tail_4 ));
    LocalMux I__5892 (
            .O(N__25321),
            .I(\tok.C_stk.tail_4 ));
    CascadeMux I__5891 (
            .O(N__25316),
            .I(\tok.C_stk.n4888_cascade_ ));
    CascadeMux I__5890 (
            .O(N__25313),
            .I(\tok.ram.n4705_cascade_ ));
    CascadeMux I__5889 (
            .O(N__25310),
            .I(\tok.n1_adj_745_cascade_ ));
    CascadeMux I__5888 (
            .O(N__25307),
            .I(N__25304));
    InMux I__5887 (
            .O(N__25304),
            .I(N__25301));
    LocalMux I__5886 (
            .O(N__25301),
            .I(N__25298));
    Span4Mux_v I__5885 (
            .O(N__25298),
            .I(N__25292));
    InMux I__5884 (
            .O(N__25297),
            .I(N__25285));
    InMux I__5883 (
            .O(N__25296),
            .I(N__25285));
    InMux I__5882 (
            .O(N__25295),
            .I(N__25285));
    Span4Mux_h I__5881 (
            .O(N__25292),
            .I(N__25280));
    LocalMux I__5880 (
            .O(N__25285),
            .I(N__25280));
    Odrv4 I__5879 (
            .O(N__25280),
            .I(\tok.tc_plus_1_4 ));
    InMux I__5878 (
            .O(N__25277),
            .I(N__25272));
    CascadeMux I__5877 (
            .O(N__25276),
            .I(N__25269));
    CascadeMux I__5876 (
            .O(N__25275),
            .I(N__25266));
    LocalMux I__5875 (
            .O(N__25272),
            .I(N__25262));
    InMux I__5874 (
            .O(N__25269),
            .I(N__25252));
    InMux I__5873 (
            .O(N__25266),
            .I(N__25252));
    InMux I__5872 (
            .O(N__25265),
            .I(N__25252));
    Span4Mux_s2_h I__5871 (
            .O(N__25262),
            .I(N__25248));
    InMux I__5870 (
            .O(N__25261),
            .I(N__25245));
    InMux I__5869 (
            .O(N__25260),
            .I(N__25242));
    CascadeMux I__5868 (
            .O(N__25259),
            .I(N__25239));
    LocalMux I__5867 (
            .O(N__25252),
            .I(N__25236));
    InMux I__5866 (
            .O(N__25251),
            .I(N__25233));
    Span4Mux_h I__5865 (
            .O(N__25248),
            .I(N__25230));
    LocalMux I__5864 (
            .O(N__25245),
            .I(N__25225));
    LocalMux I__5863 (
            .O(N__25242),
            .I(N__25225));
    InMux I__5862 (
            .O(N__25239),
            .I(N__25222));
    Span4Mux_v I__5861 (
            .O(N__25236),
            .I(N__25217));
    LocalMux I__5860 (
            .O(N__25233),
            .I(N__25217));
    Odrv4 I__5859 (
            .O(N__25230),
            .I(\tok.n802 ));
    Odrv4 I__5858 (
            .O(N__25225),
            .I(\tok.n802 ));
    LocalMux I__5857 (
            .O(N__25222),
            .I(\tok.n802 ));
    Odrv4 I__5856 (
            .O(N__25217),
            .I(\tok.n802 ));
    CascadeMux I__5855 (
            .O(N__25208),
            .I(\tok.n13_adj_746_cascade_ ));
    InMux I__5854 (
            .O(N__25205),
            .I(N__25195));
    InMux I__5853 (
            .O(N__25204),
            .I(N__25195));
    InMux I__5852 (
            .O(N__25203),
            .I(N__25195));
    InMux I__5851 (
            .O(N__25202),
            .I(N__25192));
    LocalMux I__5850 (
            .O(N__25195),
            .I(N__25184));
    LocalMux I__5849 (
            .O(N__25192),
            .I(N__25184));
    InMux I__5848 (
            .O(N__25191),
            .I(N__25180));
    InMux I__5847 (
            .O(N__25190),
            .I(N__25177));
    InMux I__5846 (
            .O(N__25189),
            .I(N__25174));
    Span4Mux_v I__5845 (
            .O(N__25184),
            .I(N__25171));
    InMux I__5844 (
            .O(N__25183),
            .I(N__25168));
    LocalMux I__5843 (
            .O(N__25180),
            .I(N__25165));
    LocalMux I__5842 (
            .O(N__25177),
            .I(N__25160));
    LocalMux I__5841 (
            .O(N__25174),
            .I(N__25160));
    Odrv4 I__5840 (
            .O(N__25171),
            .I(\tok.n86 ));
    LocalMux I__5839 (
            .O(N__25168),
            .I(\tok.n86 ));
    Odrv4 I__5838 (
            .O(N__25165),
            .I(\tok.n86 ));
    Odrv12 I__5837 (
            .O(N__25160),
            .I(\tok.n86 ));
    InMux I__5836 (
            .O(N__25151),
            .I(N__25148));
    LocalMux I__5835 (
            .O(N__25148),
            .I(N__25145));
    Span4Mux_v I__5834 (
            .O(N__25145),
            .I(N__25141));
    InMux I__5833 (
            .O(N__25144),
            .I(N__25138));
    Odrv4 I__5832 (
            .O(N__25141),
            .I(n10));
    LocalMux I__5831 (
            .O(N__25138),
            .I(n10));
    InMux I__5830 (
            .O(N__25133),
            .I(N__25129));
    InMux I__5829 (
            .O(N__25132),
            .I(N__25126));
    LocalMux I__5828 (
            .O(N__25129),
            .I(\tok.C_stk.tail_3 ));
    LocalMux I__5827 (
            .O(N__25126),
            .I(\tok.C_stk.tail_3 ));
    CascadeMux I__5826 (
            .O(N__25121),
            .I(N__25118));
    InMux I__5825 (
            .O(N__25118),
            .I(N__25115));
    LocalMux I__5824 (
            .O(N__25115),
            .I(\tok.C_stk.n4882 ));
    CascadeMux I__5823 (
            .O(N__25112),
            .I(N__25108));
    CascadeMux I__5822 (
            .O(N__25111),
            .I(N__25102));
    InMux I__5821 (
            .O(N__25108),
            .I(N__25098));
    InMux I__5820 (
            .O(N__25107),
            .I(N__25095));
    InMux I__5819 (
            .O(N__25106),
            .I(N__25092));
    CascadeMux I__5818 (
            .O(N__25105),
            .I(N__25089));
    InMux I__5817 (
            .O(N__25102),
            .I(N__25086));
    InMux I__5816 (
            .O(N__25101),
            .I(N__25083));
    LocalMux I__5815 (
            .O(N__25098),
            .I(N__25078));
    LocalMux I__5814 (
            .O(N__25095),
            .I(N__25078));
    LocalMux I__5813 (
            .O(N__25092),
            .I(N__25075));
    InMux I__5812 (
            .O(N__25089),
            .I(N__25070));
    LocalMux I__5811 (
            .O(N__25086),
            .I(N__25067));
    LocalMux I__5810 (
            .O(N__25083),
            .I(N__25062));
    Span4Mux_v I__5809 (
            .O(N__25078),
            .I(N__25062));
    Span4Mux_s3_v I__5808 (
            .O(N__25075),
            .I(N__25059));
    InMux I__5807 (
            .O(N__25074),
            .I(N__25054));
    InMux I__5806 (
            .O(N__25073),
            .I(N__25054));
    LocalMux I__5805 (
            .O(N__25070),
            .I(\tok.n602 ));
    Odrv4 I__5804 (
            .O(N__25067),
            .I(\tok.n602 ));
    Odrv4 I__5803 (
            .O(N__25062),
            .I(\tok.n602 ));
    Odrv4 I__5802 (
            .O(N__25059),
            .I(\tok.n602 ));
    LocalMux I__5801 (
            .O(N__25054),
            .I(\tok.n602 ));
    InMux I__5800 (
            .O(N__25043),
            .I(N__25038));
    InMux I__5799 (
            .O(N__25042),
            .I(N__25035));
    InMux I__5798 (
            .O(N__25041),
            .I(N__25031));
    LocalMux I__5797 (
            .O(N__25038),
            .I(N__25026));
    LocalMux I__5796 (
            .O(N__25035),
            .I(N__25026));
    InMux I__5795 (
            .O(N__25034),
            .I(N__25023));
    LocalMux I__5794 (
            .O(N__25031),
            .I(c_stk_w_7_N_18_2));
    Odrv4 I__5793 (
            .O(N__25026),
            .I(c_stk_w_7_N_18_2));
    LocalMux I__5792 (
            .O(N__25023),
            .I(c_stk_w_7_N_18_2));
    InMux I__5791 (
            .O(N__25016),
            .I(N__25012));
    InMux I__5790 (
            .O(N__25015),
            .I(N__25009));
    LocalMux I__5789 (
            .O(N__25012),
            .I(\tok.tail_61 ));
    LocalMux I__5788 (
            .O(N__25009),
            .I(\tok.tail_61 ));
    InMux I__5787 (
            .O(N__25004),
            .I(N__24998));
    InMux I__5786 (
            .O(N__25003),
            .I(N__24998));
    LocalMux I__5785 (
            .O(N__24998),
            .I(\tok.tail_45 ));
    CascadeMux I__5784 (
            .O(N__24995),
            .I(N__24992));
    InMux I__5783 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__5782 (
            .O(N__24989),
            .I(N__24986));
    Span4Mux_h I__5781 (
            .O(N__24986),
            .I(N__24982));
    InMux I__5780 (
            .O(N__24985),
            .I(N__24979));
    Odrv4 I__5779 (
            .O(N__24982),
            .I(\tok.tail_53 ));
    LocalMux I__5778 (
            .O(N__24979),
            .I(\tok.tail_53 ));
    InMux I__5777 (
            .O(N__24974),
            .I(N__24970));
    InMux I__5776 (
            .O(N__24973),
            .I(N__24967));
    LocalMux I__5775 (
            .O(N__24970),
            .I(\tok.C_stk.tail_22 ));
    LocalMux I__5774 (
            .O(N__24967),
            .I(\tok.C_stk.tail_22 ));
    InMux I__5773 (
            .O(N__24962),
            .I(N__24959));
    LocalMux I__5772 (
            .O(N__24959),
            .I(N__24956));
    Span4Mux_h I__5771 (
            .O(N__24956),
            .I(N__24953));
    Span4Mux_s2_h I__5770 (
            .O(N__24953),
            .I(N__24949));
    InMux I__5769 (
            .O(N__24952),
            .I(N__24946));
    Odrv4 I__5768 (
            .O(N__24949),
            .I(\tok.C_stk.tail_6 ));
    LocalMux I__5767 (
            .O(N__24946),
            .I(\tok.C_stk.tail_6 ));
    InMux I__5766 (
            .O(N__24941),
            .I(N__24935));
    InMux I__5765 (
            .O(N__24940),
            .I(N__24935));
    LocalMux I__5764 (
            .O(N__24935),
            .I(\tok.tail_14 ));
    InMux I__5763 (
            .O(N__24932),
            .I(N__24926));
    InMux I__5762 (
            .O(N__24931),
            .I(N__24926));
    LocalMux I__5761 (
            .O(N__24926),
            .I(\tok.tail_11 ));
    InMux I__5760 (
            .O(N__24923),
            .I(N__24917));
    InMux I__5759 (
            .O(N__24922),
            .I(N__24917));
    LocalMux I__5758 (
            .O(N__24917),
            .I(\tok.C_stk.tail_19 ));
    InMux I__5757 (
            .O(N__24914),
            .I(N__24908));
    InMux I__5756 (
            .O(N__24913),
            .I(N__24908));
    LocalMux I__5755 (
            .O(N__24908),
            .I(\tok.tail_27 ));
    InMux I__5754 (
            .O(N__24905),
            .I(N__24899));
    InMux I__5753 (
            .O(N__24904),
            .I(N__24899));
    LocalMux I__5752 (
            .O(N__24899),
            .I(\tok.C_stk.tail_35 ));
    InMux I__5751 (
            .O(N__24896),
            .I(N__24892));
    InMux I__5750 (
            .O(N__24895),
            .I(N__24889));
    LocalMux I__5749 (
            .O(N__24892),
            .I(\tok.tail_59 ));
    LocalMux I__5748 (
            .O(N__24889),
            .I(\tok.tail_59 ));
    InMux I__5747 (
            .O(N__24884),
            .I(N__24878));
    InMux I__5746 (
            .O(N__24883),
            .I(N__24878));
    LocalMux I__5745 (
            .O(N__24878),
            .I(\tok.tail_43 ));
    CascadeMux I__5744 (
            .O(N__24875),
            .I(N__24872));
    InMux I__5743 (
            .O(N__24872),
            .I(N__24869));
    LocalMux I__5742 (
            .O(N__24869),
            .I(N__24865));
    InMux I__5741 (
            .O(N__24868),
            .I(N__24862));
    Odrv4 I__5740 (
            .O(N__24865),
            .I(\tok.tail_51 ));
    LocalMux I__5739 (
            .O(N__24862),
            .I(\tok.tail_51 ));
    InMux I__5738 (
            .O(N__24857),
            .I(N__24851));
    CascadeMux I__5737 (
            .O(N__24856),
            .I(N__24848));
    InMux I__5736 (
            .O(N__24855),
            .I(N__24840));
    InMux I__5735 (
            .O(N__24854),
            .I(N__24836));
    LocalMux I__5734 (
            .O(N__24851),
            .I(N__24832));
    InMux I__5733 (
            .O(N__24848),
            .I(N__24829));
    CascadeMux I__5732 (
            .O(N__24847),
            .I(N__24826));
    InMux I__5731 (
            .O(N__24846),
            .I(N__24823));
    InMux I__5730 (
            .O(N__24845),
            .I(N__24820));
    InMux I__5729 (
            .O(N__24844),
            .I(N__24815));
    InMux I__5728 (
            .O(N__24843),
            .I(N__24815));
    LocalMux I__5727 (
            .O(N__24840),
            .I(N__24812));
    InMux I__5726 (
            .O(N__24839),
            .I(N__24809));
    LocalMux I__5725 (
            .O(N__24836),
            .I(N__24806));
    InMux I__5724 (
            .O(N__24835),
            .I(N__24803));
    Span4Mux_s3_h I__5723 (
            .O(N__24832),
            .I(N__24798));
    LocalMux I__5722 (
            .O(N__24829),
            .I(N__24798));
    InMux I__5721 (
            .O(N__24826),
            .I(N__24795));
    LocalMux I__5720 (
            .O(N__24823),
            .I(N__24791));
    LocalMux I__5719 (
            .O(N__24820),
            .I(N__24786));
    LocalMux I__5718 (
            .O(N__24815),
            .I(N__24786));
    Span4Mux_s3_h I__5717 (
            .O(N__24812),
            .I(N__24782));
    LocalMux I__5716 (
            .O(N__24809),
            .I(N__24775));
    Span4Mux_v I__5715 (
            .O(N__24806),
            .I(N__24775));
    LocalMux I__5714 (
            .O(N__24803),
            .I(N__24775));
    Span4Mux_v I__5713 (
            .O(N__24798),
            .I(N__24770));
    LocalMux I__5712 (
            .O(N__24795),
            .I(N__24770));
    InMux I__5711 (
            .O(N__24794),
            .I(N__24767));
    Span4Mux_h I__5710 (
            .O(N__24791),
            .I(N__24762));
    Span4Mux_h I__5709 (
            .O(N__24786),
            .I(N__24762));
    InMux I__5708 (
            .O(N__24785),
            .I(N__24759));
    Span4Mux_h I__5707 (
            .O(N__24782),
            .I(N__24754));
    Span4Mux_h I__5706 (
            .O(N__24775),
            .I(N__24754));
    Span4Mux_h I__5705 (
            .O(N__24770),
            .I(N__24751));
    LocalMux I__5704 (
            .O(N__24767),
            .I(N__24748));
    Odrv4 I__5703 (
            .O(N__24762),
            .I(\tok.n60 ));
    LocalMux I__5702 (
            .O(N__24759),
            .I(\tok.n60 ));
    Odrv4 I__5701 (
            .O(N__24754),
            .I(\tok.n60 ));
    Odrv4 I__5700 (
            .O(N__24751),
            .I(\tok.n60 ));
    Odrv12 I__5699 (
            .O(N__24748),
            .I(\tok.n60 ));
    InMux I__5698 (
            .O(N__24737),
            .I(N__24730));
    InMux I__5697 (
            .O(N__24736),
            .I(N__24730));
    InMux I__5696 (
            .O(N__24735),
            .I(N__24721));
    LocalMux I__5695 (
            .O(N__24730),
            .I(N__24718));
    InMux I__5694 (
            .O(N__24729),
            .I(N__24713));
    InMux I__5693 (
            .O(N__24728),
            .I(N__24713));
    InMux I__5692 (
            .O(N__24727),
            .I(N__24709));
    InMux I__5691 (
            .O(N__24726),
            .I(N__24706));
    InMux I__5690 (
            .O(N__24725),
            .I(N__24698));
    InMux I__5689 (
            .O(N__24724),
            .I(N__24698));
    LocalMux I__5688 (
            .O(N__24721),
            .I(N__24695));
    Span4Mux_v I__5687 (
            .O(N__24718),
            .I(N__24692));
    LocalMux I__5686 (
            .O(N__24713),
            .I(N__24689));
    InMux I__5685 (
            .O(N__24712),
            .I(N__24686));
    LocalMux I__5684 (
            .O(N__24709),
            .I(N__24683));
    LocalMux I__5683 (
            .O(N__24706),
            .I(N__24680));
    InMux I__5682 (
            .O(N__24705),
            .I(N__24677));
    InMux I__5681 (
            .O(N__24704),
            .I(N__24672));
    InMux I__5680 (
            .O(N__24703),
            .I(N__24672));
    LocalMux I__5679 (
            .O(N__24698),
            .I(N__24667));
    Span4Mux_s2_v I__5678 (
            .O(N__24695),
            .I(N__24667));
    Span4Mux_h I__5677 (
            .O(N__24692),
            .I(N__24660));
    Span4Mux_v I__5676 (
            .O(N__24689),
            .I(N__24660));
    LocalMux I__5675 (
            .O(N__24686),
            .I(N__24660));
    Span12Mux_s5_v I__5674 (
            .O(N__24683),
            .I(N__24652));
    Span12Mux_s5_h I__5673 (
            .O(N__24680),
            .I(N__24652));
    LocalMux I__5672 (
            .O(N__24677),
            .I(N__24652));
    LocalMux I__5671 (
            .O(N__24672),
            .I(N__24645));
    Span4Mux_h I__5670 (
            .O(N__24667),
            .I(N__24645));
    Span4Mux_h I__5669 (
            .O(N__24660),
            .I(N__24645));
    InMux I__5668 (
            .O(N__24659),
            .I(N__24642));
    Odrv12 I__5667 (
            .O(N__24652),
            .I(\tok.n83 ));
    Odrv4 I__5666 (
            .O(N__24645),
            .I(\tok.n83 ));
    LocalMux I__5665 (
            .O(N__24642),
            .I(\tok.n83 ));
    InMux I__5664 (
            .O(N__24635),
            .I(N__24632));
    LocalMux I__5663 (
            .O(N__24632),
            .I(N__24629));
    Span4Mux_s3_v I__5662 (
            .O(N__24629),
            .I(N__24626));
    Odrv4 I__5661 (
            .O(N__24626),
            .I(\tok.n3 ));
    InMux I__5660 (
            .O(N__24623),
            .I(N__24618));
    InMux I__5659 (
            .O(N__24622),
            .I(N__24615));
    CascadeMux I__5658 (
            .O(N__24621),
            .I(N__24612));
    LocalMux I__5657 (
            .O(N__24618),
            .I(N__24609));
    LocalMux I__5656 (
            .O(N__24615),
            .I(N__24606));
    InMux I__5655 (
            .O(N__24612),
            .I(N__24603));
    Span12Mux_s5_v I__5654 (
            .O(N__24609),
            .I(N__24600));
    Span4Mux_v I__5653 (
            .O(N__24606),
            .I(N__24595));
    LocalMux I__5652 (
            .O(N__24603),
            .I(N__24595));
    Odrv12 I__5651 (
            .O(N__24600),
            .I(\tok.n4478 ));
    Odrv4 I__5650 (
            .O(N__24595),
            .I(\tok.n4478 ));
    InMux I__5649 (
            .O(N__24590),
            .I(N__24586));
    CascadeMux I__5648 (
            .O(N__24589),
            .I(N__24580));
    LocalMux I__5647 (
            .O(N__24586),
            .I(N__24577));
    InMux I__5646 (
            .O(N__24585),
            .I(N__24574));
    InMux I__5645 (
            .O(N__24584),
            .I(N__24567));
    InMux I__5644 (
            .O(N__24583),
            .I(N__24567));
    InMux I__5643 (
            .O(N__24580),
            .I(N__24567));
    Odrv4 I__5642 (
            .O(N__24577),
            .I(\tok.c_stk_r_5 ));
    LocalMux I__5641 (
            .O(N__24574),
            .I(\tok.c_stk_r_5 ));
    LocalMux I__5640 (
            .O(N__24567),
            .I(\tok.c_stk_r_5 ));
    InMux I__5639 (
            .O(N__24560),
            .I(N__24557));
    LocalMux I__5638 (
            .O(N__24557),
            .I(N__24554));
    Span4Mux_h I__5637 (
            .O(N__24554),
            .I(N__24550));
    InMux I__5636 (
            .O(N__24553),
            .I(N__24547));
    Odrv4 I__5635 (
            .O(N__24550),
            .I(\tok.C_stk.tail_5 ));
    LocalMux I__5634 (
            .O(N__24547),
            .I(\tok.C_stk.tail_5 ));
    InMux I__5633 (
            .O(N__24542),
            .I(N__24536));
    InMux I__5632 (
            .O(N__24541),
            .I(N__24536));
    LocalMux I__5631 (
            .O(N__24536),
            .I(\tok.tail_13 ));
    InMux I__5630 (
            .O(N__24533),
            .I(N__24527));
    InMux I__5629 (
            .O(N__24532),
            .I(N__24527));
    LocalMux I__5628 (
            .O(N__24527),
            .I(\tok.C_stk.tail_21 ));
    CascadeMux I__5627 (
            .O(N__24524),
            .I(N__24521));
    InMux I__5626 (
            .O(N__24521),
            .I(N__24515));
    InMux I__5625 (
            .O(N__24520),
            .I(N__24515));
    LocalMux I__5624 (
            .O(N__24515),
            .I(N__24512));
    Odrv4 I__5623 (
            .O(N__24512),
            .I(\tok.tail_29 ));
    InMux I__5622 (
            .O(N__24509),
            .I(N__24503));
    InMux I__5621 (
            .O(N__24508),
            .I(N__24503));
    LocalMux I__5620 (
            .O(N__24503),
            .I(\tok.C_stk.tail_37 ));
    CascadeMux I__5619 (
            .O(N__24500),
            .I(\tok.n4460_cascade_ ));
    InMux I__5618 (
            .O(N__24497),
            .I(N__24486));
    InMux I__5617 (
            .O(N__24496),
            .I(N__24486));
    InMux I__5616 (
            .O(N__24495),
            .I(N__24482));
    InMux I__5615 (
            .O(N__24494),
            .I(N__24479));
    InMux I__5614 (
            .O(N__24493),
            .I(N__24474));
    InMux I__5613 (
            .O(N__24492),
            .I(N__24474));
    InMux I__5612 (
            .O(N__24491),
            .I(N__24466));
    LocalMux I__5611 (
            .O(N__24486),
            .I(N__24463));
    InMux I__5610 (
            .O(N__24485),
            .I(N__24460));
    LocalMux I__5609 (
            .O(N__24482),
            .I(N__24457));
    LocalMux I__5608 (
            .O(N__24479),
            .I(N__24451));
    LocalMux I__5607 (
            .O(N__24474),
            .I(N__24451));
    InMux I__5606 (
            .O(N__24473),
            .I(N__24448));
    InMux I__5605 (
            .O(N__24472),
            .I(N__24443));
    InMux I__5604 (
            .O(N__24471),
            .I(N__24443));
    InMux I__5603 (
            .O(N__24470),
            .I(N__24438));
    InMux I__5602 (
            .O(N__24469),
            .I(N__24438));
    LocalMux I__5601 (
            .O(N__24466),
            .I(N__24435));
    Span4Mux_s3_v I__5600 (
            .O(N__24463),
            .I(N__24428));
    LocalMux I__5599 (
            .O(N__24460),
            .I(N__24428));
    Span4Mux_v I__5598 (
            .O(N__24457),
            .I(N__24428));
    InMux I__5597 (
            .O(N__24456),
            .I(N__24425));
    Span4Mux_v I__5596 (
            .O(N__24451),
            .I(N__24420));
    LocalMux I__5595 (
            .O(N__24448),
            .I(N__24420));
    LocalMux I__5594 (
            .O(N__24443),
            .I(N__24415));
    LocalMux I__5593 (
            .O(N__24438),
            .I(N__24415));
    Span4Mux_s3_v I__5592 (
            .O(N__24435),
            .I(N__24408));
    Span4Mux_h I__5591 (
            .O(N__24428),
            .I(N__24408));
    LocalMux I__5590 (
            .O(N__24425),
            .I(N__24408));
    Span4Mux_h I__5589 (
            .O(N__24420),
            .I(N__24403));
    Span4Mux_v I__5588 (
            .O(N__24415),
            .I(N__24403));
    Span4Mux_h I__5587 (
            .O(N__24408),
            .I(N__24400));
    Odrv4 I__5586 (
            .O(N__24403),
            .I(\tok.n2726 ));
    Odrv4 I__5585 (
            .O(N__24400),
            .I(\tok.n2726 ));
    CascadeMux I__5584 (
            .O(N__24395),
            .I(N__24390));
    InMux I__5583 (
            .O(N__24394),
            .I(N__24386));
    CascadeMux I__5582 (
            .O(N__24393),
            .I(N__24383));
    InMux I__5581 (
            .O(N__24390),
            .I(N__24380));
    CascadeMux I__5580 (
            .O(N__24389),
            .I(N__24377));
    LocalMux I__5579 (
            .O(N__24386),
            .I(N__24372));
    InMux I__5578 (
            .O(N__24383),
            .I(N__24369));
    LocalMux I__5577 (
            .O(N__24380),
            .I(N__24363));
    InMux I__5576 (
            .O(N__24377),
            .I(N__24360));
    CascadeMux I__5575 (
            .O(N__24376),
            .I(N__24357));
    InMux I__5574 (
            .O(N__24375),
            .I(N__24354));
    Span4Mux_h I__5573 (
            .O(N__24372),
            .I(N__24349));
    LocalMux I__5572 (
            .O(N__24369),
            .I(N__24349));
    CascadeMux I__5571 (
            .O(N__24368),
            .I(N__24346));
    InMux I__5570 (
            .O(N__24367),
            .I(N__24343));
    InMux I__5569 (
            .O(N__24366),
            .I(N__24340));
    Span4Mux_s3_h I__5568 (
            .O(N__24363),
            .I(N__24335));
    LocalMux I__5567 (
            .O(N__24360),
            .I(N__24335));
    InMux I__5566 (
            .O(N__24357),
            .I(N__24332));
    LocalMux I__5565 (
            .O(N__24354),
            .I(N__24329));
    Span4Mux_v I__5564 (
            .O(N__24349),
            .I(N__24326));
    InMux I__5563 (
            .O(N__24346),
            .I(N__24323));
    LocalMux I__5562 (
            .O(N__24343),
            .I(N__24320));
    LocalMux I__5561 (
            .O(N__24340),
            .I(N__24315));
    Span4Mux_h I__5560 (
            .O(N__24335),
            .I(N__24315));
    LocalMux I__5559 (
            .O(N__24332),
            .I(N__24306));
    Span4Mux_v I__5558 (
            .O(N__24329),
            .I(N__24306));
    Span4Mux_h I__5557 (
            .O(N__24326),
            .I(N__24306));
    LocalMux I__5556 (
            .O(N__24323),
            .I(N__24306));
    Span4Mux_v I__5555 (
            .O(N__24320),
            .I(N__24303));
    Span4Mux_h I__5554 (
            .O(N__24315),
            .I(N__24300));
    Odrv4 I__5553 (
            .O(N__24306),
            .I(\tok.S_4 ));
    Odrv4 I__5552 (
            .O(N__24303),
            .I(\tok.S_4 ));
    Odrv4 I__5551 (
            .O(N__24300),
            .I(\tok.S_4 ));
    InMux I__5550 (
            .O(N__24293),
            .I(N__24290));
    LocalMux I__5549 (
            .O(N__24290),
            .I(N__24287));
    Span4Mux_s3_h I__5548 (
            .O(N__24287),
            .I(N__24284));
    Odrv4 I__5547 (
            .O(N__24284),
            .I(\tok.n13_adj_787 ));
    CascadeMux I__5546 (
            .O(N__24281),
            .I(\tok.n10_adj_829_cascade_ ));
    InMux I__5545 (
            .O(N__24278),
            .I(N__24275));
    LocalMux I__5544 (
            .O(N__24275),
            .I(N__24272));
    Odrv12 I__5543 (
            .O(N__24272),
            .I(\tok.n13_adj_833 ));
    InMux I__5542 (
            .O(N__24269),
            .I(N__24265));
    InMux I__5541 (
            .O(N__24268),
            .I(N__24262));
    LocalMux I__5540 (
            .O(N__24265),
            .I(N__24258));
    LocalMux I__5539 (
            .O(N__24262),
            .I(N__24255));
    InMux I__5538 (
            .O(N__24261),
            .I(N__24252));
    Span4Mux_v I__5537 (
            .O(N__24258),
            .I(N__24247));
    Span4Mux_v I__5536 (
            .O(N__24255),
            .I(N__24247));
    LocalMux I__5535 (
            .O(N__24252),
            .I(\tok.n2746 ));
    Odrv4 I__5534 (
            .O(N__24247),
            .I(\tok.n2746 ));
    InMux I__5533 (
            .O(N__24242),
            .I(N__24239));
    LocalMux I__5532 (
            .O(N__24239),
            .I(N__24236));
    Odrv12 I__5531 (
            .O(N__24236),
            .I(\tok.n8_adj_839 ));
    CascadeMux I__5530 (
            .O(N__24233),
            .I(N__24230));
    InMux I__5529 (
            .O(N__24230),
            .I(N__24227));
    LocalMux I__5528 (
            .O(N__24227),
            .I(N__24223));
    CascadeMux I__5527 (
            .O(N__24226),
            .I(N__24220));
    Span4Mux_s3_v I__5526 (
            .O(N__24223),
            .I(N__24217));
    InMux I__5525 (
            .O(N__24220),
            .I(N__24214));
    Span4Mux_h I__5524 (
            .O(N__24217),
            .I(N__24211));
    LocalMux I__5523 (
            .O(N__24214),
            .I(N__24208));
    Span4Mux_v I__5522 (
            .O(N__24211),
            .I(N__24205));
    Odrv12 I__5521 (
            .O(N__24208),
            .I(\tok.table_rd_0 ));
    Odrv4 I__5520 (
            .O(N__24205),
            .I(\tok.table_rd_0 ));
    InMux I__5519 (
            .O(N__24200),
            .I(N__24197));
    LocalMux I__5518 (
            .O(N__24197),
            .I(N__24194));
    Span4Mux_v I__5517 (
            .O(N__24194),
            .I(N__24191));
    Odrv4 I__5516 (
            .O(N__24191),
            .I(\tok.n18_adj_681 ));
    InMux I__5515 (
            .O(N__24188),
            .I(N__24182));
    InMux I__5514 (
            .O(N__24187),
            .I(N__24177));
    InMux I__5513 (
            .O(N__24186),
            .I(N__24174));
    InMux I__5512 (
            .O(N__24185),
            .I(N__24170));
    LocalMux I__5511 (
            .O(N__24182),
            .I(N__24165));
    InMux I__5510 (
            .O(N__24181),
            .I(N__24162));
    InMux I__5509 (
            .O(N__24180),
            .I(N__24159));
    LocalMux I__5508 (
            .O(N__24177),
            .I(N__24156));
    LocalMux I__5507 (
            .O(N__24174),
            .I(N__24153));
    InMux I__5506 (
            .O(N__24173),
            .I(N__24150));
    LocalMux I__5505 (
            .O(N__24170),
            .I(N__24146));
    InMux I__5504 (
            .O(N__24169),
            .I(N__24141));
    InMux I__5503 (
            .O(N__24168),
            .I(N__24141));
    Span4Mux_s2_v I__5502 (
            .O(N__24165),
            .I(N__24137));
    LocalMux I__5501 (
            .O(N__24162),
            .I(N__24132));
    LocalMux I__5500 (
            .O(N__24159),
            .I(N__24132));
    Span4Mux_h I__5499 (
            .O(N__24156),
            .I(N__24122));
    Span4Mux_v I__5498 (
            .O(N__24153),
            .I(N__24122));
    LocalMux I__5497 (
            .O(N__24150),
            .I(N__24122));
    CascadeMux I__5496 (
            .O(N__24149),
            .I(N__24119));
    Span4Mux_v I__5495 (
            .O(N__24146),
            .I(N__24113));
    LocalMux I__5494 (
            .O(N__24141),
            .I(N__24113));
    InMux I__5493 (
            .O(N__24140),
            .I(N__24110));
    Span4Mux_v I__5492 (
            .O(N__24137),
            .I(N__24105));
    Span4Mux_v I__5491 (
            .O(N__24132),
            .I(N__24105));
    InMux I__5490 (
            .O(N__24131),
            .I(N__24102));
    InMux I__5489 (
            .O(N__24130),
            .I(N__24097));
    InMux I__5488 (
            .O(N__24129),
            .I(N__24097));
    Span4Mux_h I__5487 (
            .O(N__24122),
            .I(N__24094));
    InMux I__5486 (
            .O(N__24119),
            .I(N__24089));
    InMux I__5485 (
            .O(N__24118),
            .I(N__24089));
    Odrv4 I__5484 (
            .O(N__24113),
            .I(\tok.A_low_1 ));
    LocalMux I__5483 (
            .O(N__24110),
            .I(\tok.A_low_1 ));
    Odrv4 I__5482 (
            .O(N__24105),
            .I(\tok.A_low_1 ));
    LocalMux I__5481 (
            .O(N__24102),
            .I(\tok.A_low_1 ));
    LocalMux I__5480 (
            .O(N__24097),
            .I(\tok.A_low_1 ));
    Odrv4 I__5479 (
            .O(N__24094),
            .I(\tok.A_low_1 ));
    LocalMux I__5478 (
            .O(N__24089),
            .I(\tok.A_low_1 ));
    InMux I__5477 (
            .O(N__24074),
            .I(N__24070));
    InMux I__5476 (
            .O(N__24073),
            .I(N__24063));
    LocalMux I__5475 (
            .O(N__24070),
            .I(N__24060));
    InMux I__5474 (
            .O(N__24069),
            .I(N__24057));
    InMux I__5473 (
            .O(N__24068),
            .I(N__24054));
    InMux I__5472 (
            .O(N__24067),
            .I(N__24051));
    InMux I__5471 (
            .O(N__24066),
            .I(N__24048));
    LocalMux I__5470 (
            .O(N__24063),
            .I(N__24045));
    Span4Mux_v I__5469 (
            .O(N__24060),
            .I(N__24042));
    LocalMux I__5468 (
            .O(N__24057),
            .I(N__24039));
    LocalMux I__5467 (
            .O(N__24054),
            .I(N__24036));
    LocalMux I__5466 (
            .O(N__24051),
            .I(N__24031));
    LocalMux I__5465 (
            .O(N__24048),
            .I(N__24031));
    Span4Mux_v I__5464 (
            .O(N__24045),
            .I(N__24022));
    Span4Mux_h I__5463 (
            .O(N__24042),
            .I(N__24022));
    Span4Mux_v I__5462 (
            .O(N__24039),
            .I(N__24022));
    Span4Mux_s2_h I__5461 (
            .O(N__24036),
            .I(N__24022));
    Span4Mux_v I__5460 (
            .O(N__24031),
            .I(N__24019));
    Odrv4 I__5459 (
            .O(N__24022),
            .I(\tok.n101 ));
    Odrv4 I__5458 (
            .O(N__24019),
            .I(\tok.n101 ));
    CascadeMux I__5457 (
            .O(N__24014),
            .I(N__24010));
    InMux I__5456 (
            .O(N__24013),
            .I(N__24005));
    InMux I__5455 (
            .O(N__24010),
            .I(N__24000));
    CascadeMux I__5454 (
            .O(N__24009),
            .I(N__23997));
    InMux I__5453 (
            .O(N__24008),
            .I(N__23994));
    LocalMux I__5452 (
            .O(N__24005),
            .I(N__23991));
    InMux I__5451 (
            .O(N__24004),
            .I(N__23988));
    InMux I__5450 (
            .O(N__24003),
            .I(N__23985));
    LocalMux I__5449 (
            .O(N__24000),
            .I(N__23979));
    InMux I__5448 (
            .O(N__23997),
            .I(N__23976));
    LocalMux I__5447 (
            .O(N__23994),
            .I(N__23971));
    Span4Mux_v I__5446 (
            .O(N__23991),
            .I(N__23971));
    LocalMux I__5445 (
            .O(N__23988),
            .I(N__23968));
    LocalMux I__5444 (
            .O(N__23985),
            .I(N__23965));
    InMux I__5443 (
            .O(N__23984),
            .I(N__23962));
    InMux I__5442 (
            .O(N__23983),
            .I(N__23959));
    CascadeMux I__5441 (
            .O(N__23982),
            .I(N__23956));
    Span4Mux_h I__5440 (
            .O(N__23979),
            .I(N__23953));
    LocalMux I__5439 (
            .O(N__23976),
            .I(N__23947));
    Span4Mux_h I__5438 (
            .O(N__23971),
            .I(N__23947));
    Span4Mux_h I__5437 (
            .O(N__23968),
            .I(N__23942));
    Span4Mux_v I__5436 (
            .O(N__23965),
            .I(N__23942));
    LocalMux I__5435 (
            .O(N__23962),
            .I(N__23937));
    LocalMux I__5434 (
            .O(N__23959),
            .I(N__23937));
    InMux I__5433 (
            .O(N__23956),
            .I(N__23934));
    Span4Mux_h I__5432 (
            .O(N__23953),
            .I(N__23931));
    InMux I__5431 (
            .O(N__23952),
            .I(N__23928));
    Span4Mux_v I__5430 (
            .O(N__23947),
            .I(N__23925));
    Odrv4 I__5429 (
            .O(N__23942),
            .I(\tok.n54 ));
    Odrv12 I__5428 (
            .O(N__23937),
            .I(\tok.n54 ));
    LocalMux I__5427 (
            .O(N__23934),
            .I(\tok.n54 ));
    Odrv4 I__5426 (
            .O(N__23931),
            .I(\tok.n54 ));
    LocalMux I__5425 (
            .O(N__23928),
            .I(\tok.n54 ));
    Odrv4 I__5424 (
            .O(N__23925),
            .I(\tok.n54 ));
    CascadeMux I__5423 (
            .O(N__23912),
            .I(\tok.n244_cascade_ ));
    InMux I__5422 (
            .O(N__23909),
            .I(N__23906));
    LocalMux I__5421 (
            .O(N__23906),
            .I(N__23903));
    Odrv12 I__5420 (
            .O(N__23903),
            .I(\tok.n17_adj_785 ));
    InMux I__5419 (
            .O(N__23900),
            .I(N__23890));
    InMux I__5418 (
            .O(N__23899),
            .I(N__23879));
    InMux I__5417 (
            .O(N__23898),
            .I(N__23879));
    InMux I__5416 (
            .O(N__23897),
            .I(N__23879));
    InMux I__5415 (
            .O(N__23896),
            .I(N__23879));
    InMux I__5414 (
            .O(N__23895),
            .I(N__23879));
    CascadeMux I__5413 (
            .O(N__23894),
            .I(N__23872));
    InMux I__5412 (
            .O(N__23893),
            .I(N__23862));
    LocalMux I__5411 (
            .O(N__23890),
            .I(N__23859));
    LocalMux I__5410 (
            .O(N__23879),
            .I(N__23856));
    InMux I__5409 (
            .O(N__23878),
            .I(N__23847));
    InMux I__5408 (
            .O(N__23877),
            .I(N__23847));
    InMux I__5407 (
            .O(N__23876),
            .I(N__23847));
    InMux I__5406 (
            .O(N__23875),
            .I(N__23847));
    InMux I__5405 (
            .O(N__23872),
            .I(N__23838));
    InMux I__5404 (
            .O(N__23871),
            .I(N__23838));
    InMux I__5403 (
            .O(N__23870),
            .I(N__23838));
    InMux I__5402 (
            .O(N__23869),
            .I(N__23838));
    InMux I__5401 (
            .O(N__23868),
            .I(N__23833));
    InMux I__5400 (
            .O(N__23867),
            .I(N__23833));
    InMux I__5399 (
            .O(N__23866),
            .I(N__23828));
    InMux I__5398 (
            .O(N__23865),
            .I(N__23828));
    LocalMux I__5397 (
            .O(N__23862),
            .I(N__23825));
    Span4Mux_v I__5396 (
            .O(N__23859),
            .I(N__23818));
    Span4Mux_v I__5395 (
            .O(N__23856),
            .I(N__23818));
    LocalMux I__5394 (
            .O(N__23847),
            .I(N__23818));
    LocalMux I__5393 (
            .O(N__23838),
            .I(N__23815));
    LocalMux I__5392 (
            .O(N__23833),
            .I(N__23812));
    LocalMux I__5391 (
            .O(N__23828),
            .I(N__23809));
    Span4Mux_v I__5390 (
            .O(N__23825),
            .I(N__23802));
    Span4Mux_h I__5389 (
            .O(N__23818),
            .I(N__23802));
    Span4Mux_v I__5388 (
            .O(N__23815),
            .I(N__23802));
    Span4Mux_v I__5387 (
            .O(N__23812),
            .I(N__23798));
    Span4Mux_h I__5386 (
            .O(N__23809),
            .I(N__23795));
    Span4Mux_h I__5385 (
            .O(N__23802),
            .I(N__23792));
    InMux I__5384 (
            .O(N__23801),
            .I(N__23789));
    Odrv4 I__5383 (
            .O(N__23798),
            .I(\tok.n11_adj_647 ));
    Odrv4 I__5382 (
            .O(N__23795),
            .I(\tok.n11_adj_647 ));
    Odrv4 I__5381 (
            .O(N__23792),
            .I(\tok.n11_adj_647 ));
    LocalMux I__5380 (
            .O(N__23789),
            .I(\tok.n11_adj_647 ));
    CascadeMux I__5379 (
            .O(N__23780),
            .I(\tok.n4575_cascade_ ));
    CascadeMux I__5378 (
            .O(N__23777),
            .I(\tok.n83_cascade_ ));
    InMux I__5377 (
            .O(N__23774),
            .I(N__23768));
    InMux I__5376 (
            .O(N__23773),
            .I(N__23768));
    LocalMux I__5375 (
            .O(N__23768),
            .I(N__23765));
    Span4Mux_s3_h I__5374 (
            .O(N__23765),
            .I(N__23762));
    Odrv4 I__5373 (
            .O(N__23762),
            .I(\tok.n40 ));
    CascadeMux I__5372 (
            .O(N__23759),
            .I(\tok.n4571_cascade_ ));
    InMux I__5371 (
            .O(N__23756),
            .I(N__23753));
    LocalMux I__5370 (
            .O(N__23753),
            .I(\tok.n4393 ));
    InMux I__5369 (
            .O(N__23750),
            .I(N__23747));
    LocalMux I__5368 (
            .O(N__23747),
            .I(N__23741));
    InMux I__5367 (
            .O(N__23746),
            .I(N__23736));
    InMux I__5366 (
            .O(N__23745),
            .I(N__23736));
    InMux I__5365 (
            .O(N__23744),
            .I(N__23733));
    Span4Mux_v I__5364 (
            .O(N__23741),
            .I(N__23728));
    LocalMux I__5363 (
            .O(N__23736),
            .I(N__23728));
    LocalMux I__5362 (
            .O(N__23733),
            .I(N__23725));
    Span4Mux_h I__5361 (
            .O(N__23728),
            .I(N__23720));
    Span4Mux_h I__5360 (
            .O(N__23725),
            .I(N__23720));
    Odrv4 I__5359 (
            .O(N__23720),
            .I(\tok.n9_adj_797 ));
    InMux I__5358 (
            .O(N__23717),
            .I(N__23714));
    LocalMux I__5357 (
            .O(N__23714),
            .I(\tok.n13_adj_758 ));
    InMux I__5356 (
            .O(N__23711),
            .I(N__23708));
    LocalMux I__5355 (
            .O(N__23708),
            .I(N__23705));
    Odrv12 I__5354 (
            .O(N__23705),
            .I(n10_adj_873));
    CascadeMux I__5353 (
            .O(N__23702),
            .I(n10_adj_873_cascade_));
    CascadeMux I__5352 (
            .O(N__23699),
            .I(N__23696));
    InMux I__5351 (
            .O(N__23696),
            .I(N__23693));
    LocalMux I__5350 (
            .O(N__23693),
            .I(N__23688));
    InMux I__5349 (
            .O(N__23692),
            .I(N__23685));
    InMux I__5348 (
            .O(N__23691),
            .I(N__23681));
    Span4Mux_s3_h I__5347 (
            .O(N__23688),
            .I(N__23678));
    LocalMux I__5346 (
            .O(N__23685),
            .I(N__23675));
    InMux I__5345 (
            .O(N__23684),
            .I(N__23672));
    LocalMux I__5344 (
            .O(N__23681),
            .I(c_stk_w_7_N_18_5));
    Odrv4 I__5343 (
            .O(N__23678),
            .I(c_stk_w_7_N_18_5));
    Odrv12 I__5342 (
            .O(N__23675),
            .I(c_stk_w_7_N_18_5));
    LocalMux I__5341 (
            .O(N__23672),
            .I(c_stk_w_7_N_18_5));
    CascadeMux I__5340 (
            .O(N__23663),
            .I(N__23660));
    InMux I__5339 (
            .O(N__23660),
            .I(N__23657));
    LocalMux I__5338 (
            .O(N__23657),
            .I(\tok.tc_5 ));
    InMux I__5337 (
            .O(N__23654),
            .I(N__23651));
    LocalMux I__5336 (
            .O(N__23651),
            .I(N__23648));
    Span4Mux_h I__5335 (
            .O(N__23648),
            .I(N__23645));
    Odrv4 I__5334 (
            .O(N__23645),
            .I(n10_adj_874));
    CascadeMux I__5333 (
            .O(N__23642),
            .I(n10_adj_874_cascade_));
    CascadeMux I__5332 (
            .O(N__23639),
            .I(N__23636));
    InMux I__5331 (
            .O(N__23636),
            .I(N__23633));
    LocalMux I__5330 (
            .O(N__23633),
            .I(N__23630));
    Odrv4 I__5329 (
            .O(N__23630),
            .I(\tok.tc_2 ));
    CascadeMux I__5328 (
            .O(N__23627),
            .I(N__23624));
    InMux I__5327 (
            .O(N__23624),
            .I(N__23621));
    LocalMux I__5326 (
            .O(N__23621),
            .I(N__23616));
    InMux I__5325 (
            .O(N__23620),
            .I(N__23610));
    InMux I__5324 (
            .O(N__23619),
            .I(N__23610));
    Span4Mux_v I__5323 (
            .O(N__23616),
            .I(N__23607));
    InMux I__5322 (
            .O(N__23615),
            .I(N__23604));
    LocalMux I__5321 (
            .O(N__23610),
            .I(N__23601));
    Span4Mux_v I__5320 (
            .O(N__23607),
            .I(N__23598));
    LocalMux I__5319 (
            .O(N__23604),
            .I(N__23595));
    Span4Mux_s3_h I__5318 (
            .O(N__23601),
            .I(N__23592));
    Odrv4 I__5317 (
            .O(N__23598),
            .I(\tok.tc_plus_1_3 ));
    Odrv4 I__5316 (
            .O(N__23595),
            .I(\tok.tc_plus_1_3 ));
    Odrv4 I__5315 (
            .O(N__23592),
            .I(\tok.tc_plus_1_3 ));
    CascadeMux I__5314 (
            .O(N__23585),
            .I(N__23582));
    InMux I__5313 (
            .O(N__23582),
            .I(N__23579));
    LocalMux I__5312 (
            .O(N__23579),
            .I(N__23576));
    Odrv4 I__5311 (
            .O(N__23576),
            .I(n92_adj_870));
    CascadeMux I__5310 (
            .O(N__23573),
            .I(n92_adj_870_cascade_));
    CascadeMux I__5309 (
            .O(N__23570),
            .I(N__23567));
    InMux I__5308 (
            .O(N__23567),
            .I(N__23564));
    LocalMux I__5307 (
            .O(N__23564),
            .I(N__23559));
    InMux I__5306 (
            .O(N__23563),
            .I(N__23556));
    InMux I__5305 (
            .O(N__23562),
            .I(N__23552));
    Span4Mux_v I__5304 (
            .O(N__23559),
            .I(N__23549));
    LocalMux I__5303 (
            .O(N__23556),
            .I(N__23546));
    InMux I__5302 (
            .O(N__23555),
            .I(N__23543));
    LocalMux I__5301 (
            .O(N__23552),
            .I(c_stk_w_7_N_18_3));
    Odrv4 I__5300 (
            .O(N__23549),
            .I(c_stk_w_7_N_18_3));
    Odrv12 I__5299 (
            .O(N__23546),
            .I(c_stk_w_7_N_18_3));
    LocalMux I__5298 (
            .O(N__23543),
            .I(c_stk_w_7_N_18_3));
    CascadeMux I__5297 (
            .O(N__23534),
            .I(N__23531));
    InMux I__5296 (
            .O(N__23531),
            .I(N__23528));
    LocalMux I__5295 (
            .O(N__23528),
            .I(N__23525));
    Odrv4 I__5294 (
            .O(N__23525),
            .I(\tok.tc_3 ));
    InMux I__5293 (
            .O(N__23522),
            .I(N__23507));
    InMux I__5292 (
            .O(N__23521),
            .I(N__23507));
    InMux I__5291 (
            .O(N__23520),
            .I(N__23507));
    InMux I__5290 (
            .O(N__23519),
            .I(N__23507));
    InMux I__5289 (
            .O(N__23518),
            .I(N__23493));
    InMux I__5288 (
            .O(N__23517),
            .I(N__23493));
    InMux I__5287 (
            .O(N__23516),
            .I(N__23490));
    LocalMux I__5286 (
            .O(N__23507),
            .I(N__23487));
    InMux I__5285 (
            .O(N__23506),
            .I(N__23470));
    InMux I__5284 (
            .O(N__23505),
            .I(N__23470));
    InMux I__5283 (
            .O(N__23504),
            .I(N__23470));
    InMux I__5282 (
            .O(N__23503),
            .I(N__23470));
    InMux I__5281 (
            .O(N__23502),
            .I(N__23470));
    InMux I__5280 (
            .O(N__23501),
            .I(N__23470));
    InMux I__5279 (
            .O(N__23500),
            .I(N__23470));
    InMux I__5278 (
            .O(N__23499),
            .I(N__23470));
    InMux I__5277 (
            .O(N__23498),
            .I(N__23467));
    LocalMux I__5276 (
            .O(N__23493),
            .I(N__23464));
    LocalMux I__5275 (
            .O(N__23490),
            .I(N__23461));
    Span4Mux_v I__5274 (
            .O(N__23487),
            .I(N__23458));
    LocalMux I__5273 (
            .O(N__23470),
            .I(stall_));
    LocalMux I__5272 (
            .O(N__23467),
            .I(stall_));
    Odrv4 I__5271 (
            .O(N__23464),
            .I(stall_));
    Odrv4 I__5270 (
            .O(N__23461),
            .I(stall_));
    Odrv4 I__5269 (
            .O(N__23458),
            .I(stall_));
    CascadeMux I__5268 (
            .O(N__23447),
            .I(N__23444));
    InMux I__5267 (
            .O(N__23444),
            .I(N__23441));
    LocalMux I__5266 (
            .O(N__23441),
            .I(\tok.tc_4 ));
    CascadeMux I__5265 (
            .O(N__23438),
            .I(\tok.C_stk.n4900_cascade_ ));
    CascadeMux I__5264 (
            .O(N__23435),
            .I(N__23432));
    InMux I__5263 (
            .O(N__23432),
            .I(N__23429));
    LocalMux I__5262 (
            .O(N__23429),
            .I(N__23425));
    InMux I__5261 (
            .O(N__23428),
            .I(N__23422));
    Span4Mux_v I__5260 (
            .O(N__23425),
            .I(N__23419));
    LocalMux I__5259 (
            .O(N__23422),
            .I(N__23416));
    Span4Mux_h I__5258 (
            .O(N__23419),
            .I(N__23413));
    Span4Mux_v I__5257 (
            .O(N__23416),
            .I(N__23410));
    Span4Mux_h I__5256 (
            .O(N__23413),
            .I(N__23407));
    Odrv4 I__5255 (
            .O(N__23410),
            .I(\tok.table_rd_5 ));
    Odrv4 I__5254 (
            .O(N__23407),
            .I(\tok.table_rd_5 ));
    CascadeMux I__5253 (
            .O(N__23402),
            .I(\tok.n83_adj_742_cascade_ ));
    CascadeMux I__5252 (
            .O(N__23399),
            .I(\tok.n4651_cascade_ ));
    CascadeMux I__5251 (
            .O(N__23396),
            .I(\tok.ram.n4702_cascade_ ));
    InMux I__5250 (
            .O(N__23393),
            .I(N__23390));
    LocalMux I__5249 (
            .O(N__23390),
            .I(\tok.n1_adj_757 ));
    CascadeMux I__5248 (
            .O(N__23387),
            .I(N__23384));
    InMux I__5247 (
            .O(N__23384),
            .I(N__23380));
    InMux I__5246 (
            .O(N__23383),
            .I(N__23377));
    LocalMux I__5245 (
            .O(N__23380),
            .I(N__23374));
    LocalMux I__5244 (
            .O(N__23377),
            .I(N__23369));
    Span4Mux_v I__5243 (
            .O(N__23374),
            .I(N__23366));
    InMux I__5242 (
            .O(N__23373),
            .I(N__23361));
    InMux I__5241 (
            .O(N__23372),
            .I(N__23361));
    Span4Mux_v I__5240 (
            .O(N__23369),
            .I(N__23356));
    Span4Mux_s2_h I__5239 (
            .O(N__23366),
            .I(N__23356));
    LocalMux I__5238 (
            .O(N__23361),
            .I(N__23353));
    Odrv4 I__5237 (
            .O(N__23356),
            .I(\tok.tc_plus_1_5 ));
    Odrv4 I__5236 (
            .O(N__23353),
            .I(\tok.tc_plus_1_5 ));
    InMux I__5235 (
            .O(N__23348),
            .I(N__23345));
    LocalMux I__5234 (
            .O(N__23345),
            .I(N__23341));
    InMux I__5233 (
            .O(N__23344),
            .I(N__23338));
    Span4Mux_v I__5232 (
            .O(N__23341),
            .I(N__23335));
    LocalMux I__5231 (
            .O(N__23338),
            .I(\tok.tail_44 ));
    Odrv4 I__5230 (
            .O(N__23335),
            .I(\tok.tail_44 ));
    InMux I__5229 (
            .O(N__23330),
            .I(N__23327));
    LocalMux I__5228 (
            .O(N__23327),
            .I(N__23324));
    Span4Mux_s3_h I__5227 (
            .O(N__23324),
            .I(N__23320));
    InMux I__5226 (
            .O(N__23323),
            .I(N__23317));
    Odrv4 I__5225 (
            .O(N__23320),
            .I(\tok.C_stk.tail_18 ));
    LocalMux I__5224 (
            .O(N__23317),
            .I(\tok.C_stk.tail_18 ));
    CascadeMux I__5223 (
            .O(N__23312),
            .I(N__23308));
    InMux I__5222 (
            .O(N__23311),
            .I(N__23303));
    InMux I__5221 (
            .O(N__23308),
            .I(N__23303));
    LocalMux I__5220 (
            .O(N__23303),
            .I(N__23300));
    Span4Mux_s2_h I__5219 (
            .O(N__23300),
            .I(N__23297));
    Span4Mux_h I__5218 (
            .O(N__23297),
            .I(N__23294));
    Odrv4 I__5217 (
            .O(N__23294),
            .I(\tok.n240 ));
    CascadeMux I__5216 (
            .O(N__23291),
            .I(N__23287));
    InMux I__5215 (
            .O(N__23290),
            .I(N__23284));
    InMux I__5214 (
            .O(N__23287),
            .I(N__23281));
    LocalMux I__5213 (
            .O(N__23284),
            .I(N__23278));
    LocalMux I__5212 (
            .O(N__23281),
            .I(N__23275));
    Odrv4 I__5211 (
            .O(N__23278),
            .I(\tok.tail_55 ));
    Odrv12 I__5210 (
            .O(N__23275),
            .I(\tok.tail_55 ));
    InMux I__5209 (
            .O(N__23270),
            .I(N__23267));
    LocalMux I__5208 (
            .O(N__23267),
            .I(N__23263));
    InMux I__5207 (
            .O(N__23266),
            .I(N__23260));
    Odrv4 I__5206 (
            .O(N__23263),
            .I(\tok.tail_63 ));
    LocalMux I__5205 (
            .O(N__23260),
            .I(\tok.tail_63 ));
    InMux I__5204 (
            .O(N__23255),
            .I(N__23251));
    InMux I__5203 (
            .O(N__23254),
            .I(N__23248));
    LocalMux I__5202 (
            .O(N__23251),
            .I(\tok.tail_54 ));
    LocalMux I__5201 (
            .O(N__23248),
            .I(\tok.tail_54 ));
    InMux I__5200 (
            .O(N__23243),
            .I(N__23239));
    InMux I__5199 (
            .O(N__23242),
            .I(N__23236));
    LocalMux I__5198 (
            .O(N__23239),
            .I(\tok.tail_62 ));
    LocalMux I__5197 (
            .O(N__23236),
            .I(\tok.tail_62 ));
    InMux I__5196 (
            .O(N__23231),
            .I(N__23227));
    InMux I__5195 (
            .O(N__23230),
            .I(N__23224));
    LocalMux I__5194 (
            .O(N__23227),
            .I(N__23221));
    LocalMux I__5193 (
            .O(N__23224),
            .I(N__23218));
    Span4Mux_h I__5192 (
            .O(N__23221),
            .I(N__23215));
    Odrv4 I__5191 (
            .O(N__23218),
            .I(\tok.tail_52 ));
    Odrv4 I__5190 (
            .O(N__23215),
            .I(\tok.tail_52 ));
    InMux I__5189 (
            .O(N__23210),
            .I(N__23206));
    InMux I__5188 (
            .O(N__23209),
            .I(N__23203));
    LocalMux I__5187 (
            .O(N__23206),
            .I(\tok.tail_60 ));
    LocalMux I__5186 (
            .O(N__23203),
            .I(\tok.tail_60 ));
    InMux I__5185 (
            .O(N__23198),
            .I(N__23192));
    InMux I__5184 (
            .O(N__23197),
            .I(N__23192));
    LocalMux I__5183 (
            .O(N__23192),
            .I(\tok.C_stk.tail_39 ));
    InMux I__5182 (
            .O(N__23189),
            .I(N__23183));
    InMux I__5181 (
            .O(N__23188),
            .I(N__23183));
    LocalMux I__5180 (
            .O(N__23183),
            .I(\tok.tail_47 ));
    InMux I__5179 (
            .O(N__23180),
            .I(N__23174));
    InMux I__5178 (
            .O(N__23179),
            .I(N__23174));
    LocalMux I__5177 (
            .O(N__23174),
            .I(\tok.C_stk.tail_16 ));
    InMux I__5176 (
            .O(N__23171),
            .I(N__23168));
    LocalMux I__5175 (
            .O(N__23168),
            .I(N__23164));
    InMux I__5174 (
            .O(N__23167),
            .I(N__23161));
    Odrv4 I__5173 (
            .O(N__23164),
            .I(\tok.C_stk.tail_32 ));
    LocalMux I__5172 (
            .O(N__23161),
            .I(\tok.C_stk.tail_32 ));
    InMux I__5171 (
            .O(N__23156),
            .I(N__23152));
    InMux I__5170 (
            .O(N__23155),
            .I(N__23149));
    LocalMux I__5169 (
            .O(N__23152),
            .I(N__23146));
    LocalMux I__5168 (
            .O(N__23149),
            .I(\tok.tail_24 ));
    Odrv4 I__5167 (
            .O(N__23146),
            .I(\tok.tail_24 ));
    CascadeMux I__5166 (
            .O(N__23141),
            .I(N__23138));
    InMux I__5165 (
            .O(N__23138),
            .I(N__23132));
    InMux I__5164 (
            .O(N__23137),
            .I(N__23132));
    LocalMux I__5163 (
            .O(N__23132),
            .I(\tok.tail_30 ));
    InMux I__5162 (
            .O(N__23129),
            .I(N__23123));
    InMux I__5161 (
            .O(N__23128),
            .I(N__23123));
    LocalMux I__5160 (
            .O(N__23123),
            .I(\tok.C_stk.tail_38 ));
    InMux I__5159 (
            .O(N__23120),
            .I(N__23114));
    InMux I__5158 (
            .O(N__23119),
            .I(N__23114));
    LocalMux I__5157 (
            .O(N__23114),
            .I(\tok.tail_46 ));
    InMux I__5156 (
            .O(N__23111),
            .I(N__23107));
    InMux I__5155 (
            .O(N__23110),
            .I(N__23103));
    LocalMux I__5154 (
            .O(N__23107),
            .I(N__23100));
    CascadeMux I__5153 (
            .O(N__23106),
            .I(N__23095));
    LocalMux I__5152 (
            .O(N__23103),
            .I(N__23092));
    Span4Mux_h I__5151 (
            .O(N__23100),
            .I(N__23089));
    InMux I__5150 (
            .O(N__23099),
            .I(N__23086));
    InMux I__5149 (
            .O(N__23098),
            .I(N__23081));
    InMux I__5148 (
            .O(N__23095),
            .I(N__23081));
    Span4Mux_v I__5147 (
            .O(N__23092),
            .I(N__23078));
    Odrv4 I__5146 (
            .O(N__23089),
            .I(\tok.c_stk_r_6 ));
    LocalMux I__5145 (
            .O(N__23086),
            .I(\tok.c_stk_r_6 ));
    LocalMux I__5144 (
            .O(N__23081),
            .I(\tok.c_stk_r_6 ));
    Odrv4 I__5143 (
            .O(N__23078),
            .I(\tok.c_stk_r_6 ));
    InMux I__5142 (
            .O(N__23069),
            .I(N__23066));
    LocalMux I__5141 (
            .O(N__23066),
            .I(N__23063));
    Span12Mux_s6_v I__5140 (
            .O(N__23063),
            .I(N__23060));
    Odrv12 I__5139 (
            .O(N__23060),
            .I(\tok.n9_adj_807 ));
    InMux I__5138 (
            .O(N__23057),
            .I(N__23051));
    InMux I__5137 (
            .O(N__23056),
            .I(N__23051));
    LocalMux I__5136 (
            .O(N__23051),
            .I(uart_rx_data_4));
    InMux I__5135 (
            .O(N__23048),
            .I(N__23045));
    LocalMux I__5134 (
            .O(N__23045),
            .I(N__23042));
    Span4Mux_h I__5133 (
            .O(N__23042),
            .I(N__23039));
    Span4Mux_h I__5132 (
            .O(N__23039),
            .I(N__23036));
    Odrv4 I__5131 (
            .O(N__23036),
            .I(\tok.n3_adj_826 ));
    CascadeMux I__5130 (
            .O(N__23033),
            .I(\tok.n6_adj_827_cascade_ ));
    InMux I__5129 (
            .O(N__23030),
            .I(N__23027));
    LocalMux I__5128 (
            .O(N__23027),
            .I(N__23024));
    Odrv4 I__5127 (
            .O(N__23024),
            .I(\tok.n36 ));
    CascadeMux I__5126 (
            .O(N__23021),
            .I(\tok.n33_adj_828_cascade_ ));
    InMux I__5125 (
            .O(N__23018),
            .I(N__23015));
    LocalMux I__5124 (
            .O(N__23015),
            .I(N__23012));
    Span4Mux_h I__5123 (
            .O(N__23012),
            .I(N__23009));
    Odrv4 I__5122 (
            .O(N__23009),
            .I(\tok.n11_adj_831 ));
    InMux I__5121 (
            .O(N__23006),
            .I(N__23000));
    InMux I__5120 (
            .O(N__23005),
            .I(N__22997));
    InMux I__5119 (
            .O(N__23004),
            .I(N__22989));
    InMux I__5118 (
            .O(N__23003),
            .I(N__22989));
    LocalMux I__5117 (
            .O(N__23000),
            .I(N__22986));
    LocalMux I__5116 (
            .O(N__22997),
            .I(N__22983));
    InMux I__5115 (
            .O(N__22996),
            .I(N__22980));
    InMux I__5114 (
            .O(N__22995),
            .I(N__22976));
    InMux I__5113 (
            .O(N__22994),
            .I(N__22973));
    LocalMux I__5112 (
            .O(N__22989),
            .I(N__22970));
    Span4Mux_s1_v I__5111 (
            .O(N__22986),
            .I(N__22966));
    Span4Mux_v I__5110 (
            .O(N__22983),
            .I(N__22961));
    LocalMux I__5109 (
            .O(N__22980),
            .I(N__22961));
    InMux I__5108 (
            .O(N__22979),
            .I(N__22958));
    LocalMux I__5107 (
            .O(N__22976),
            .I(N__22955));
    LocalMux I__5106 (
            .O(N__22973),
            .I(N__22952));
    Span4Mux_v I__5105 (
            .O(N__22970),
            .I(N__22949));
    InMux I__5104 (
            .O(N__22969),
            .I(N__22946));
    Span4Mux_v I__5103 (
            .O(N__22966),
            .I(N__22939));
    Span4Mux_h I__5102 (
            .O(N__22961),
            .I(N__22939));
    LocalMux I__5101 (
            .O(N__22958),
            .I(N__22939));
    Span4Mux_h I__5100 (
            .O(N__22955),
            .I(N__22936));
    Span4Mux_s3_v I__5099 (
            .O(N__22952),
            .I(N__22933));
    Span4Mux_h I__5098 (
            .O(N__22949),
            .I(N__22925));
    LocalMux I__5097 (
            .O(N__22946),
            .I(N__22925));
    Span4Mux_v I__5096 (
            .O(N__22939),
            .I(N__22925));
    Span4Mux_v I__5095 (
            .O(N__22936),
            .I(N__22920));
    Span4Mux_h I__5094 (
            .O(N__22933),
            .I(N__22920));
    InMux I__5093 (
            .O(N__22932),
            .I(N__22917));
    Span4Mux_h I__5092 (
            .O(N__22925),
            .I(N__22914));
    Odrv4 I__5091 (
            .O(N__22920),
            .I(\tok.n56 ));
    LocalMux I__5090 (
            .O(N__22917),
            .I(\tok.n56 ));
    Odrv4 I__5089 (
            .O(N__22914),
            .I(\tok.n56 ));
    InMux I__5088 (
            .O(N__22907),
            .I(N__22904));
    LocalMux I__5087 (
            .O(N__22904),
            .I(N__22901));
    Span4Mux_h I__5086 (
            .O(N__22901),
            .I(N__22898));
    Span4Mux_h I__5085 (
            .O(N__22898),
            .I(N__22895));
    Odrv4 I__5084 (
            .O(N__22895),
            .I(\tok.n2514 ));
    InMux I__5083 (
            .O(N__22892),
            .I(N__22889));
    LocalMux I__5082 (
            .O(N__22889),
            .I(N__22885));
    InMux I__5081 (
            .O(N__22888),
            .I(N__22882));
    Span4Mux_s3_h I__5080 (
            .O(N__22885),
            .I(N__22879));
    LocalMux I__5079 (
            .O(N__22882),
            .I(\tok.C_stk.tail_0 ));
    Odrv4 I__5078 (
            .O(N__22879),
            .I(\tok.C_stk.tail_0 ));
    InMux I__5077 (
            .O(N__22874),
            .I(N__22871));
    LocalMux I__5076 (
            .O(N__22871),
            .I(N__22868));
    Span4Mux_s1_v I__5075 (
            .O(N__22868),
            .I(N__22864));
    InMux I__5074 (
            .O(N__22867),
            .I(N__22861));
    Odrv4 I__5073 (
            .O(N__22864),
            .I(\tok.tail_8 ));
    LocalMux I__5072 (
            .O(N__22861),
            .I(\tok.tail_8 ));
    InMux I__5071 (
            .O(N__22856),
            .I(N__22852));
    CascadeMux I__5070 (
            .O(N__22855),
            .I(N__22849));
    LocalMux I__5069 (
            .O(N__22852),
            .I(N__22846));
    InMux I__5068 (
            .O(N__22849),
            .I(N__22843));
    Odrv4 I__5067 (
            .O(N__22846),
            .I(\tok.tail_15 ));
    LocalMux I__5066 (
            .O(N__22843),
            .I(\tok.tail_15 ));
    InMux I__5065 (
            .O(N__22838),
            .I(N__22835));
    LocalMux I__5064 (
            .O(N__22835),
            .I(N__22832));
    Span4Mux_s1_v I__5063 (
            .O(N__22832),
            .I(N__22828));
    InMux I__5062 (
            .O(N__22831),
            .I(N__22825));
    Odrv4 I__5061 (
            .O(N__22828),
            .I(\tok.C_stk.tail_23 ));
    LocalMux I__5060 (
            .O(N__22825),
            .I(\tok.C_stk.tail_23 ));
    InMux I__5059 (
            .O(N__22820),
            .I(N__22814));
    InMux I__5058 (
            .O(N__22819),
            .I(N__22814));
    LocalMux I__5057 (
            .O(N__22814),
            .I(\tok.tail_31 ));
    InMux I__5056 (
            .O(N__22811),
            .I(N__22808));
    LocalMux I__5055 (
            .O(N__22808),
            .I(\tok.n211 ));
    InMux I__5054 (
            .O(N__22805),
            .I(N__22802));
    LocalMux I__5053 (
            .O(N__22802),
            .I(N__22799));
    Odrv4 I__5052 (
            .O(N__22799),
            .I(\tok.n2_adj_810 ));
    InMux I__5051 (
            .O(N__22796),
            .I(N__22793));
    LocalMux I__5050 (
            .O(N__22793),
            .I(N__22790));
    Odrv4 I__5049 (
            .O(N__22790),
            .I(\tok.n5_adj_710 ));
    InMux I__5048 (
            .O(N__22787),
            .I(N__22784));
    LocalMux I__5047 (
            .O(N__22784),
            .I(N__22781));
    Span4Mux_h I__5046 (
            .O(N__22781),
            .I(N__22778));
    Odrv4 I__5045 (
            .O(N__22778),
            .I(\tok.n6_adj_711 ));
    InMux I__5044 (
            .O(N__22775),
            .I(N__22772));
    LocalMux I__5043 (
            .O(N__22772),
            .I(N__22769));
    Span12Mux_s7_h I__5042 (
            .O(N__22769),
            .I(N__22766));
    Odrv12 I__5041 (
            .O(N__22766),
            .I(\tok.n4664 ));
    InMux I__5040 (
            .O(N__22763),
            .I(N__22760));
    LocalMux I__5039 (
            .O(N__22760),
            .I(N__22757));
    Odrv4 I__5038 (
            .O(N__22757),
            .I(\tok.n4663 ));
    InMux I__5037 (
            .O(N__22754),
            .I(N__22751));
    LocalMux I__5036 (
            .O(N__22751),
            .I(\tok.n33 ));
    InMux I__5035 (
            .O(N__22748),
            .I(N__22745));
    LocalMux I__5034 (
            .O(N__22745),
            .I(N__22742));
    Odrv12 I__5033 (
            .O(N__22742),
            .I(\tok.n27 ));
    CascadeMux I__5032 (
            .O(N__22739),
            .I(N__22736));
    InMux I__5031 (
            .O(N__22736),
            .I(N__22733));
    LocalMux I__5030 (
            .O(N__22733),
            .I(N__22730));
    Span4Mux_h I__5029 (
            .O(N__22730),
            .I(N__22727));
    Span4Mux_h I__5028 (
            .O(N__22727),
            .I(N__22724));
    Odrv4 I__5027 (
            .O(N__22724),
            .I(\tok.n296 ));
    InMux I__5026 (
            .O(N__22721),
            .I(N__22713));
    InMux I__5025 (
            .O(N__22720),
            .I(N__22710));
    InMux I__5024 (
            .O(N__22719),
            .I(N__22705));
    InMux I__5023 (
            .O(N__22718),
            .I(N__22705));
    InMux I__5022 (
            .O(N__22717),
            .I(N__22702));
    CascadeMux I__5021 (
            .O(N__22716),
            .I(N__22698));
    LocalMux I__5020 (
            .O(N__22713),
            .I(N__22694));
    LocalMux I__5019 (
            .O(N__22710),
            .I(N__22691));
    LocalMux I__5018 (
            .O(N__22705),
            .I(N__22688));
    LocalMux I__5017 (
            .O(N__22702),
            .I(N__22685));
    InMux I__5016 (
            .O(N__22701),
            .I(N__22680));
    InMux I__5015 (
            .O(N__22698),
            .I(N__22680));
    InMux I__5014 (
            .O(N__22697),
            .I(N__22677));
    Span4Mux_h I__5013 (
            .O(N__22694),
            .I(N__22672));
    Span4Mux_v I__5012 (
            .O(N__22691),
            .I(N__22672));
    Span12Mux_s5_h I__5011 (
            .O(N__22688),
            .I(N__22665));
    Span12Mux_s11_v I__5010 (
            .O(N__22685),
            .I(N__22665));
    LocalMux I__5009 (
            .O(N__22680),
            .I(N__22665));
    LocalMux I__5008 (
            .O(N__22677),
            .I(\tok.n191 ));
    Odrv4 I__5007 (
            .O(N__22672),
            .I(\tok.n191 ));
    Odrv12 I__5006 (
            .O(N__22665),
            .I(\tok.n191 ));
    CascadeMux I__5005 (
            .O(N__22658),
            .I(N__22652));
    InMux I__5004 (
            .O(N__22657),
            .I(N__22647));
    InMux I__5003 (
            .O(N__22656),
            .I(N__22644));
    InMux I__5002 (
            .O(N__22655),
            .I(N__22641));
    InMux I__5001 (
            .O(N__22652),
            .I(N__22637));
    InMux I__5000 (
            .O(N__22651),
            .I(N__22633));
    InMux I__4999 (
            .O(N__22650),
            .I(N__22628));
    LocalMux I__4998 (
            .O(N__22647),
            .I(N__22625));
    LocalMux I__4997 (
            .O(N__22644),
            .I(N__22622));
    LocalMux I__4996 (
            .O(N__22641),
            .I(N__22619));
    InMux I__4995 (
            .O(N__22640),
            .I(N__22616));
    LocalMux I__4994 (
            .O(N__22637),
            .I(N__22613));
    InMux I__4993 (
            .O(N__22636),
            .I(N__22610));
    LocalMux I__4992 (
            .O(N__22633),
            .I(N__22607));
    InMux I__4991 (
            .O(N__22632),
            .I(N__22604));
    InMux I__4990 (
            .O(N__22631),
            .I(N__22601));
    LocalMux I__4989 (
            .O(N__22628),
            .I(N__22598));
    Span4Mux_v I__4988 (
            .O(N__22625),
            .I(N__22593));
    Span4Mux_v I__4987 (
            .O(N__22622),
            .I(N__22593));
    Span4Mux_h I__4986 (
            .O(N__22619),
            .I(N__22590));
    LocalMux I__4985 (
            .O(N__22616),
            .I(N__22583));
    Span4Mux_h I__4984 (
            .O(N__22613),
            .I(N__22583));
    LocalMux I__4983 (
            .O(N__22610),
            .I(N__22580));
    Span4Mux_s2_h I__4982 (
            .O(N__22607),
            .I(N__22577));
    LocalMux I__4981 (
            .O(N__22604),
            .I(N__22566));
    LocalMux I__4980 (
            .O(N__22601),
            .I(N__22566));
    Span4Mux_v I__4979 (
            .O(N__22598),
            .I(N__22566));
    Span4Mux_h I__4978 (
            .O(N__22593),
            .I(N__22566));
    Span4Mux_v I__4977 (
            .O(N__22590),
            .I(N__22566));
    InMux I__4976 (
            .O(N__22589),
            .I(N__22561));
    InMux I__4975 (
            .O(N__22588),
            .I(N__22561));
    Span4Mux_h I__4974 (
            .O(N__22583),
            .I(N__22558));
    Span4Mux_h I__4973 (
            .O(N__22580),
            .I(N__22555));
    Span4Mux_v I__4972 (
            .O(N__22577),
            .I(N__22550));
    Span4Mux_h I__4971 (
            .O(N__22566),
            .I(N__22550));
    LocalMux I__4970 (
            .O(N__22561),
            .I(\tok.n59 ));
    Odrv4 I__4969 (
            .O(N__22558),
            .I(\tok.n59 ));
    Odrv4 I__4968 (
            .O(N__22555),
            .I(\tok.n59 ));
    Odrv4 I__4967 (
            .O(N__22550),
            .I(\tok.n59 ));
    CascadeMux I__4966 (
            .O(N__22541),
            .I(N__22538));
    InMux I__4965 (
            .O(N__22538),
            .I(N__22535));
    LocalMux I__4964 (
            .O(N__22535),
            .I(N__22532));
    Odrv4 I__4963 (
            .O(N__22532),
            .I(\tok.n2_adj_703 ));
    CascadeMux I__4962 (
            .O(N__22529),
            .I(N__22523));
    InMux I__4961 (
            .O(N__22528),
            .I(N__22516));
    InMux I__4960 (
            .O(N__22527),
            .I(N__22513));
    InMux I__4959 (
            .O(N__22526),
            .I(N__22508));
    InMux I__4958 (
            .O(N__22523),
            .I(N__22508));
    CascadeMux I__4957 (
            .O(N__22522),
            .I(N__22504));
    InMux I__4956 (
            .O(N__22521),
            .I(N__22500));
    InMux I__4955 (
            .O(N__22520),
            .I(N__22497));
    InMux I__4954 (
            .O(N__22519),
            .I(N__22494));
    LocalMux I__4953 (
            .O(N__22516),
            .I(N__22486));
    LocalMux I__4952 (
            .O(N__22513),
            .I(N__22481));
    LocalMux I__4951 (
            .O(N__22508),
            .I(N__22481));
    InMux I__4950 (
            .O(N__22507),
            .I(N__22474));
    InMux I__4949 (
            .O(N__22504),
            .I(N__22474));
    InMux I__4948 (
            .O(N__22503),
            .I(N__22474));
    LocalMux I__4947 (
            .O(N__22500),
            .I(N__22469));
    LocalMux I__4946 (
            .O(N__22497),
            .I(N__22469));
    LocalMux I__4945 (
            .O(N__22494),
            .I(N__22466));
    InMux I__4944 (
            .O(N__22493),
            .I(N__22461));
    InMux I__4943 (
            .O(N__22492),
            .I(N__22461));
    InMux I__4942 (
            .O(N__22491),
            .I(N__22458));
    InMux I__4941 (
            .O(N__22490),
            .I(N__22455));
    CascadeMux I__4940 (
            .O(N__22489),
            .I(N__22452));
    Span4Mux_s3_v I__4939 (
            .O(N__22486),
            .I(N__22443));
    Span4Mux_s3_v I__4938 (
            .O(N__22481),
            .I(N__22443));
    LocalMux I__4937 (
            .O(N__22474),
            .I(N__22443));
    Span4Mux_s2_v I__4936 (
            .O(N__22469),
            .I(N__22440));
    Span4Mux_v I__4935 (
            .O(N__22466),
            .I(N__22435));
    LocalMux I__4934 (
            .O(N__22461),
            .I(N__22435));
    LocalMux I__4933 (
            .O(N__22458),
            .I(N__22430));
    LocalMux I__4932 (
            .O(N__22455),
            .I(N__22430));
    InMux I__4931 (
            .O(N__22452),
            .I(N__22427));
    InMux I__4930 (
            .O(N__22451),
            .I(N__22422));
    InMux I__4929 (
            .O(N__22450),
            .I(N__22422));
    Span4Mux_v I__4928 (
            .O(N__22443),
            .I(N__22417));
    Span4Mux_v I__4927 (
            .O(N__22440),
            .I(N__22417));
    Span4Mux_h I__4926 (
            .O(N__22435),
            .I(N__22414));
    Odrv12 I__4925 (
            .O(N__22430),
            .I(\tok.stall ));
    LocalMux I__4924 (
            .O(N__22427),
            .I(\tok.stall ));
    LocalMux I__4923 (
            .O(N__22422),
            .I(\tok.stall ));
    Odrv4 I__4922 (
            .O(N__22417),
            .I(\tok.stall ));
    Odrv4 I__4921 (
            .O(N__22414),
            .I(\tok.stall ));
    CascadeMux I__4920 (
            .O(N__22403),
            .I(N__22397));
    InMux I__4919 (
            .O(N__22402),
            .I(N__22394));
    InMux I__4918 (
            .O(N__22401),
            .I(N__22390));
    InMux I__4917 (
            .O(N__22400),
            .I(N__22386));
    InMux I__4916 (
            .O(N__22397),
            .I(N__22383));
    LocalMux I__4915 (
            .O(N__22394),
            .I(N__22380));
    InMux I__4914 (
            .O(N__22393),
            .I(N__22377));
    LocalMux I__4913 (
            .O(N__22390),
            .I(N__22370));
    InMux I__4912 (
            .O(N__22389),
            .I(N__22367));
    LocalMux I__4911 (
            .O(N__22386),
            .I(N__22361));
    LocalMux I__4910 (
            .O(N__22383),
            .I(N__22361));
    Span4Mux_v I__4909 (
            .O(N__22380),
            .I(N__22358));
    LocalMux I__4908 (
            .O(N__22377),
            .I(N__22355));
    InMux I__4907 (
            .O(N__22376),
            .I(N__22350));
    InMux I__4906 (
            .O(N__22375),
            .I(N__22350));
    CascadeMux I__4905 (
            .O(N__22374),
            .I(N__22346));
    InMux I__4904 (
            .O(N__22373),
            .I(N__22343));
    Span4Mux_v I__4903 (
            .O(N__22370),
            .I(N__22338));
    LocalMux I__4902 (
            .O(N__22367),
            .I(N__22338));
    InMux I__4901 (
            .O(N__22366),
            .I(N__22335));
    Span4Mux_v I__4900 (
            .O(N__22361),
            .I(N__22329));
    Span4Mux_v I__4899 (
            .O(N__22358),
            .I(N__22322));
    Span4Mux_s2_v I__4898 (
            .O(N__22355),
            .I(N__22322));
    LocalMux I__4897 (
            .O(N__22350),
            .I(N__22322));
    InMux I__4896 (
            .O(N__22349),
            .I(N__22317));
    InMux I__4895 (
            .O(N__22346),
            .I(N__22317));
    LocalMux I__4894 (
            .O(N__22343),
            .I(N__22312));
    Span4Mux_h I__4893 (
            .O(N__22338),
            .I(N__22312));
    LocalMux I__4892 (
            .O(N__22335),
            .I(N__22309));
    InMux I__4891 (
            .O(N__22334),
            .I(N__22304));
    InMux I__4890 (
            .O(N__22333),
            .I(N__22304));
    InMux I__4889 (
            .O(N__22332),
            .I(N__22301));
    Span4Mux_h I__4888 (
            .O(N__22329),
            .I(N__22298));
    Odrv4 I__4887 (
            .O(N__22322),
            .I(\tok.A_low_5 ));
    LocalMux I__4886 (
            .O(N__22317),
            .I(\tok.A_low_5 ));
    Odrv4 I__4885 (
            .O(N__22312),
            .I(\tok.A_low_5 ));
    Odrv12 I__4884 (
            .O(N__22309),
            .I(\tok.A_low_5 ));
    LocalMux I__4883 (
            .O(N__22304),
            .I(\tok.A_low_5 ));
    LocalMux I__4882 (
            .O(N__22301),
            .I(\tok.A_low_5 ));
    Odrv4 I__4881 (
            .O(N__22298),
            .I(\tok.A_low_5 ));
    CascadeMux I__4880 (
            .O(N__22283),
            .I(N__22278));
    CascadeMux I__4879 (
            .O(N__22282),
            .I(N__22274));
    CascadeMux I__4878 (
            .O(N__22281),
            .I(N__22269));
    InMux I__4877 (
            .O(N__22278),
            .I(N__22266));
    CascadeMux I__4876 (
            .O(N__22277),
            .I(N__22263));
    InMux I__4875 (
            .O(N__22274),
            .I(N__22254));
    InMux I__4874 (
            .O(N__22273),
            .I(N__22254));
    InMux I__4873 (
            .O(N__22272),
            .I(N__22254));
    InMux I__4872 (
            .O(N__22269),
            .I(N__22251));
    LocalMux I__4871 (
            .O(N__22266),
            .I(N__22248));
    InMux I__4870 (
            .O(N__22263),
            .I(N__22245));
    InMux I__4869 (
            .O(N__22262),
            .I(N__22240));
    InMux I__4868 (
            .O(N__22261),
            .I(N__22240));
    LocalMux I__4867 (
            .O(N__22254),
            .I(N__22232));
    LocalMux I__4866 (
            .O(N__22251),
            .I(N__22232));
    Span4Mux_h I__4865 (
            .O(N__22248),
            .I(N__22229));
    LocalMux I__4864 (
            .O(N__22245),
            .I(N__22226));
    LocalMux I__4863 (
            .O(N__22240),
            .I(N__22223));
    InMux I__4862 (
            .O(N__22239),
            .I(N__22216));
    InMux I__4861 (
            .O(N__22238),
            .I(N__22216));
    InMux I__4860 (
            .O(N__22237),
            .I(N__22216));
    Span12Mux_s6_h I__4859 (
            .O(N__22232),
            .I(N__22213));
    Span4Mux_v I__4858 (
            .O(N__22229),
            .I(N__22210));
    Span4Mux_s3_v I__4857 (
            .O(N__22226),
            .I(N__22205));
    Span4Mux_h I__4856 (
            .O(N__22223),
            .I(N__22205));
    LocalMux I__4855 (
            .O(N__22216),
            .I(\tok.search_clk ));
    Odrv12 I__4854 (
            .O(N__22213),
            .I(\tok.search_clk ));
    Odrv4 I__4853 (
            .O(N__22210),
            .I(\tok.search_clk ));
    Odrv4 I__4852 (
            .O(N__22205),
            .I(\tok.search_clk ));
    InMux I__4851 (
            .O(N__22196),
            .I(N__22193));
    LocalMux I__4850 (
            .O(N__22193),
            .I(\tok.n33_adj_817 ));
    InMux I__4849 (
            .O(N__22190),
            .I(N__22187));
    LocalMux I__4848 (
            .O(N__22187),
            .I(N__22184));
    Odrv12 I__4847 (
            .O(N__22184),
            .I(\tok.n27_adj_868 ));
    InMux I__4846 (
            .O(N__22181),
            .I(N__22178));
    LocalMux I__4845 (
            .O(N__22178),
            .I(N__22172));
    InMux I__4844 (
            .O(N__22177),
            .I(N__22169));
    InMux I__4843 (
            .O(N__22176),
            .I(N__22164));
    InMux I__4842 (
            .O(N__22175),
            .I(N__22164));
    Span4Mux_h I__4841 (
            .O(N__22172),
            .I(N__22161));
    LocalMux I__4840 (
            .O(N__22169),
            .I(N__22158));
    LocalMux I__4839 (
            .O(N__22164),
            .I(N__22155));
    Odrv4 I__4838 (
            .O(N__22161),
            .I(\tok.n82 ));
    Odrv4 I__4837 (
            .O(N__22158),
            .I(\tok.n82 ));
    Odrv4 I__4836 (
            .O(N__22155),
            .I(\tok.n82 ));
    InMux I__4835 (
            .O(N__22148),
            .I(N__22145));
    LocalMux I__4834 (
            .O(N__22145),
            .I(N__22142));
    Span4Mux_h I__4833 (
            .O(N__22142),
            .I(N__22139));
    Span4Mux_h I__4832 (
            .O(N__22139),
            .I(N__22134));
    InMux I__4831 (
            .O(N__22138),
            .I(N__22129));
    InMux I__4830 (
            .O(N__22137),
            .I(N__22129));
    Odrv4 I__4829 (
            .O(N__22134),
            .I(capture_5));
    LocalMux I__4828 (
            .O(N__22129),
            .I(capture_5));
    InMux I__4827 (
            .O(N__22124),
            .I(N__22118));
    InMux I__4826 (
            .O(N__22123),
            .I(N__22115));
    InMux I__4825 (
            .O(N__22122),
            .I(N__22109));
    InMux I__4824 (
            .O(N__22121),
            .I(N__22106));
    LocalMux I__4823 (
            .O(N__22118),
            .I(N__22103));
    LocalMux I__4822 (
            .O(N__22115),
            .I(N__22098));
    InMux I__4821 (
            .O(N__22114),
            .I(N__22095));
    InMux I__4820 (
            .O(N__22113),
            .I(N__22092));
    InMux I__4819 (
            .O(N__22112),
            .I(N__22089));
    LocalMux I__4818 (
            .O(N__22109),
            .I(N__22086));
    LocalMux I__4817 (
            .O(N__22106),
            .I(N__22083));
    Span4Mux_h I__4816 (
            .O(N__22103),
            .I(N__22080));
    InMux I__4815 (
            .O(N__22102),
            .I(N__22075));
    InMux I__4814 (
            .O(N__22101),
            .I(N__22075));
    Span4Mux_v I__4813 (
            .O(N__22098),
            .I(N__22072));
    LocalMux I__4812 (
            .O(N__22095),
            .I(N__22069));
    LocalMux I__4811 (
            .O(N__22092),
            .I(N__22064));
    LocalMux I__4810 (
            .O(N__22089),
            .I(N__22064));
    Span4Mux_h I__4809 (
            .O(N__22086),
            .I(N__22061));
    Span4Mux_v I__4808 (
            .O(N__22083),
            .I(N__22058));
    Span4Mux_h I__4807 (
            .O(N__22080),
            .I(N__22053));
    LocalMux I__4806 (
            .O(N__22075),
            .I(N__22053));
    Span4Mux_h I__4805 (
            .O(N__22072),
            .I(N__22046));
    Span4Mux_v I__4804 (
            .O(N__22069),
            .I(N__22046));
    Span4Mux_h I__4803 (
            .O(N__22064),
            .I(N__22046));
    Span4Mux_h I__4802 (
            .O(N__22061),
            .I(N__22043));
    Span4Mux_v I__4801 (
            .O(N__22058),
            .I(N__22038));
    Span4Mux_v I__4800 (
            .O(N__22053),
            .I(N__22038));
    Span4Mux_h I__4799 (
            .O(N__22046),
            .I(N__22035));
    Odrv4 I__4798 (
            .O(N__22043),
            .I(rx_data_7__N_511));
    Odrv4 I__4797 (
            .O(N__22038),
            .I(rx_data_7__N_511));
    Odrv4 I__4796 (
            .O(N__22035),
            .I(rx_data_7__N_511));
    InMux I__4795 (
            .O(N__22028),
            .I(N__22025));
    LocalMux I__4794 (
            .O(N__22025),
            .I(N__22022));
    Odrv4 I__4793 (
            .O(N__22022),
            .I(\tok.n13_adj_816 ));
    InMux I__4792 (
            .O(N__22019),
            .I(\tok.n3902 ));
    InMux I__4791 (
            .O(N__22016),
            .I(N__22013));
    LocalMux I__4790 (
            .O(N__22013),
            .I(N__22010));
    Odrv4 I__4789 (
            .O(N__22010),
            .I(\tok.n2_adj_811 ));
    InMux I__4788 (
            .O(N__22007),
            .I(\tok.n3903 ));
    InMux I__4787 (
            .O(N__22004),
            .I(N__22001));
    LocalMux I__4786 (
            .O(N__22001),
            .I(\tok.n26_adj_808 ));
    InMux I__4785 (
            .O(N__21998),
            .I(\tok.n3904 ));
    InMux I__4784 (
            .O(N__21995),
            .I(\tok.n3905 ));
    InMux I__4783 (
            .O(N__21992),
            .I(\tok.n3906 ));
    InMux I__4782 (
            .O(N__21989),
            .I(N__21982));
    InMux I__4781 (
            .O(N__21988),
            .I(N__21978));
    InMux I__4780 (
            .O(N__21987),
            .I(N__21973));
    InMux I__4779 (
            .O(N__21986),
            .I(N__21968));
    InMux I__4778 (
            .O(N__21985),
            .I(N__21964));
    LocalMux I__4777 (
            .O(N__21982),
            .I(N__21961));
    InMux I__4776 (
            .O(N__21981),
            .I(N__21958));
    LocalMux I__4775 (
            .O(N__21978),
            .I(N__21954));
    InMux I__4774 (
            .O(N__21977),
            .I(N__21949));
    InMux I__4773 (
            .O(N__21976),
            .I(N__21949));
    LocalMux I__4772 (
            .O(N__21973),
            .I(N__21946));
    InMux I__4771 (
            .O(N__21972),
            .I(N__21943));
    CascadeMux I__4770 (
            .O(N__21971),
            .I(N__21939));
    LocalMux I__4769 (
            .O(N__21968),
            .I(N__21934));
    InMux I__4768 (
            .O(N__21967),
            .I(N__21931));
    LocalMux I__4767 (
            .O(N__21964),
            .I(N__21924));
    Span4Mux_v I__4766 (
            .O(N__21961),
            .I(N__21924));
    LocalMux I__4765 (
            .O(N__21958),
            .I(N__21924));
    InMux I__4764 (
            .O(N__21957),
            .I(N__21921));
    Span4Mux_v I__4763 (
            .O(N__21954),
            .I(N__21916));
    LocalMux I__4762 (
            .O(N__21949),
            .I(N__21916));
    Span4Mux_h I__4761 (
            .O(N__21946),
            .I(N__21913));
    LocalMux I__4760 (
            .O(N__21943),
            .I(N__21910));
    InMux I__4759 (
            .O(N__21942),
            .I(N__21907));
    InMux I__4758 (
            .O(N__21939),
            .I(N__21904));
    InMux I__4757 (
            .O(N__21938),
            .I(N__21901));
    InMux I__4756 (
            .O(N__21937),
            .I(N__21898));
    Span4Mux_v I__4755 (
            .O(N__21934),
            .I(N__21893));
    LocalMux I__4754 (
            .O(N__21931),
            .I(N__21893));
    Span4Mux_h I__4753 (
            .O(N__21924),
            .I(N__21890));
    LocalMux I__4752 (
            .O(N__21921),
            .I(N__21885));
    Span4Mux_h I__4751 (
            .O(N__21916),
            .I(N__21885));
    Odrv4 I__4750 (
            .O(N__21913),
            .I(\tok.A_low_2 ));
    Odrv12 I__4749 (
            .O(N__21910),
            .I(\tok.A_low_2 ));
    LocalMux I__4748 (
            .O(N__21907),
            .I(\tok.A_low_2 ));
    LocalMux I__4747 (
            .O(N__21904),
            .I(\tok.A_low_2 ));
    LocalMux I__4746 (
            .O(N__21901),
            .I(\tok.A_low_2 ));
    LocalMux I__4745 (
            .O(N__21898),
            .I(\tok.A_low_2 ));
    Odrv4 I__4744 (
            .O(N__21893),
            .I(\tok.A_low_2 ));
    Odrv4 I__4743 (
            .O(N__21890),
            .I(\tok.A_low_2 ));
    Odrv4 I__4742 (
            .O(N__21885),
            .I(\tok.A_low_2 ));
    InMux I__4741 (
            .O(N__21866),
            .I(N__21863));
    LocalMux I__4740 (
            .O(N__21863),
            .I(N__21860));
    Span4Mux_h I__4739 (
            .O(N__21860),
            .I(N__21857));
    Odrv4 I__4738 (
            .O(N__21857),
            .I(\tok.n210 ));
    InMux I__4737 (
            .O(N__21854),
            .I(\tok.n3907 ));
    InMux I__4736 (
            .O(N__21851),
            .I(N__21847));
    InMux I__4735 (
            .O(N__21850),
            .I(N__21842));
    LocalMux I__4734 (
            .O(N__21847),
            .I(N__21836));
    InMux I__4733 (
            .O(N__21846),
            .I(N__21833));
    InMux I__4732 (
            .O(N__21845),
            .I(N__21828));
    LocalMux I__4731 (
            .O(N__21842),
            .I(N__21825));
    InMux I__4730 (
            .O(N__21841),
            .I(N__21820));
    InMux I__4729 (
            .O(N__21840),
            .I(N__21817));
    InMux I__4728 (
            .O(N__21839),
            .I(N__21814));
    Span4Mux_v I__4727 (
            .O(N__21836),
            .I(N__21808));
    LocalMux I__4726 (
            .O(N__21833),
            .I(N__21808));
    InMux I__4725 (
            .O(N__21832),
            .I(N__21803));
    InMux I__4724 (
            .O(N__21831),
            .I(N__21803));
    LocalMux I__4723 (
            .O(N__21828),
            .I(N__21800));
    Span4Mux_v I__4722 (
            .O(N__21825),
            .I(N__21797));
    InMux I__4721 (
            .O(N__21824),
            .I(N__21791));
    InMux I__4720 (
            .O(N__21823),
            .I(N__21788));
    LocalMux I__4719 (
            .O(N__21820),
            .I(N__21785));
    LocalMux I__4718 (
            .O(N__21817),
            .I(N__21782));
    LocalMux I__4717 (
            .O(N__21814),
            .I(N__21779));
    InMux I__4716 (
            .O(N__21813),
            .I(N__21776));
    Span4Mux_h I__4715 (
            .O(N__21808),
            .I(N__21773));
    LocalMux I__4714 (
            .O(N__21803),
            .I(N__21770));
    Span4Mux_h I__4713 (
            .O(N__21800),
            .I(N__21767));
    Sp12to4 I__4712 (
            .O(N__21797),
            .I(N__21764));
    InMux I__4711 (
            .O(N__21796),
            .I(N__21761));
    InMux I__4710 (
            .O(N__21795),
            .I(N__21758));
    InMux I__4709 (
            .O(N__21794),
            .I(N__21755));
    LocalMux I__4708 (
            .O(N__21791),
            .I(N__21752));
    LocalMux I__4707 (
            .O(N__21788),
            .I(N__21743));
    Span4Mux_h I__4706 (
            .O(N__21785),
            .I(N__21743));
    Span4Mux_h I__4705 (
            .O(N__21782),
            .I(N__21743));
    Span4Mux_v I__4704 (
            .O(N__21779),
            .I(N__21743));
    LocalMux I__4703 (
            .O(N__21776),
            .I(N__21736));
    Span4Mux_v I__4702 (
            .O(N__21773),
            .I(N__21736));
    Span4Mux_h I__4701 (
            .O(N__21770),
            .I(N__21736));
    Odrv4 I__4700 (
            .O(N__21767),
            .I(\tok.A_low_3 ));
    Odrv12 I__4699 (
            .O(N__21764),
            .I(\tok.A_low_3 ));
    LocalMux I__4698 (
            .O(N__21761),
            .I(\tok.A_low_3 ));
    LocalMux I__4697 (
            .O(N__21758),
            .I(\tok.A_low_3 ));
    LocalMux I__4696 (
            .O(N__21755),
            .I(\tok.A_low_3 ));
    Odrv4 I__4695 (
            .O(N__21752),
            .I(\tok.A_low_3 ));
    Odrv4 I__4694 (
            .O(N__21743),
            .I(\tok.A_low_3 ));
    Odrv4 I__4693 (
            .O(N__21736),
            .I(\tok.A_low_3 ));
    InMux I__4692 (
            .O(N__21719),
            .I(N__21716));
    LocalMux I__4691 (
            .O(N__21716),
            .I(N__21713));
    Span4Mux_h I__4690 (
            .O(N__21713),
            .I(N__21710));
    Span4Mux_h I__4689 (
            .O(N__21710),
            .I(N__21707));
    Odrv4 I__4688 (
            .O(N__21707),
            .I(\tok.n209 ));
    InMux I__4687 (
            .O(N__21704),
            .I(\tok.n3908 ));
    DummyBuf I__4686 (
            .O(N__21701),
            .I(N__21695));
    DummyBuf I__4685 (
            .O(N__21700),
            .I(N__21692));
    SRMux I__4684 (
            .O(N__21699),
            .I(N__21686));
    SRMux I__4683 (
            .O(N__21698),
            .I(N__21682));
    InMux I__4682 (
            .O(N__21695),
            .I(N__21678));
    InMux I__4681 (
            .O(N__21692),
            .I(N__21675));
    CascadeMux I__4680 (
            .O(N__21691),
            .I(N__21672));
    CascadeMux I__4679 (
            .O(N__21690),
            .I(N__21669));
    CascadeMux I__4678 (
            .O(N__21689),
            .I(N__21666));
    LocalMux I__4677 (
            .O(N__21686),
            .I(N__21662));
    InMux I__4676 (
            .O(N__21685),
            .I(N__21659));
    LocalMux I__4675 (
            .O(N__21682),
            .I(N__21656));
    SRMux I__4674 (
            .O(N__21681),
            .I(N__21653));
    LocalMux I__4673 (
            .O(N__21678),
            .I(N__21650));
    LocalMux I__4672 (
            .O(N__21675),
            .I(N__21647));
    InMux I__4671 (
            .O(N__21672),
            .I(N__21644));
    InMux I__4670 (
            .O(N__21669),
            .I(N__21639));
    InMux I__4669 (
            .O(N__21666),
            .I(N__21639));
    InMux I__4668 (
            .O(N__21665),
            .I(N__21636));
    Span4Mux_v I__4667 (
            .O(N__21662),
            .I(N__21633));
    LocalMux I__4666 (
            .O(N__21659),
            .I(N__21630));
    Span4Mux_v I__4665 (
            .O(N__21656),
            .I(N__21625));
    LocalMux I__4664 (
            .O(N__21653),
            .I(N__21625));
    Span4Mux_s3_v I__4663 (
            .O(N__21650),
            .I(N__21620));
    Span4Mux_s3_v I__4662 (
            .O(N__21647),
            .I(N__21620));
    LocalMux I__4661 (
            .O(N__21644),
            .I(N__21617));
    LocalMux I__4660 (
            .O(N__21639),
            .I(N__21614));
    LocalMux I__4659 (
            .O(N__21636),
            .I(N__21611));
    Span4Mux_h I__4658 (
            .O(N__21633),
            .I(N__21607));
    Span4Mux_v I__4657 (
            .O(N__21630),
            .I(N__21604));
    Span4Mux_v I__4656 (
            .O(N__21625),
            .I(N__21601));
    Span4Mux_v I__4655 (
            .O(N__21620),
            .I(N__21598));
    Span4Mux_v I__4654 (
            .O(N__21617),
            .I(N__21591));
    Span4Mux_v I__4653 (
            .O(N__21614),
            .I(N__21591));
    Span4Mux_h I__4652 (
            .O(N__21611),
            .I(N__21591));
    InMux I__4651 (
            .O(N__21610),
            .I(N__21588));
    Span4Mux_h I__4650 (
            .O(N__21607),
            .I(N__21585));
    Span4Mux_h I__4649 (
            .O(N__21604),
            .I(N__21582));
    Span4Mux_s2_v I__4648 (
            .O(N__21601),
            .I(N__21579));
    Span4Mux_v I__4647 (
            .O(N__21598),
            .I(N__21572));
    Span4Mux_h I__4646 (
            .O(N__21591),
            .I(N__21572));
    LocalMux I__4645 (
            .O(N__21588),
            .I(N__21572));
    Odrv4 I__4644 (
            .O(N__21585),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4643 (
            .O(N__21582),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4642 (
            .O(N__21579),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4641 (
            .O(N__21572),
            .I(CONSTANT_ONE_NET));
    InMux I__4640 (
            .O(N__21563),
            .I(bfn_9_12_0_));
    InMux I__4639 (
            .O(N__21560),
            .I(N__21557));
    LocalMux I__4638 (
            .O(N__21557),
            .I(\tok.n2598 ));
    CascadeMux I__4637 (
            .O(N__21554),
            .I(\tok.n5_adj_837_cascade_ ));
    CascadeMux I__4636 (
            .O(N__21551),
            .I(N__21547));
    CascadeMux I__4635 (
            .O(N__21550),
            .I(N__21541));
    InMux I__4634 (
            .O(N__21547),
            .I(N__21535));
    InMux I__4633 (
            .O(N__21546),
            .I(N__21532));
    InMux I__4632 (
            .O(N__21545),
            .I(N__21529));
    CascadeMux I__4631 (
            .O(N__21544),
            .I(N__21526));
    InMux I__4630 (
            .O(N__21541),
            .I(N__21523));
    CascadeMux I__4629 (
            .O(N__21540),
            .I(N__21520));
    InMux I__4628 (
            .O(N__21539),
            .I(N__21517));
    InMux I__4627 (
            .O(N__21538),
            .I(N__21514));
    LocalMux I__4626 (
            .O(N__21535),
            .I(N__21511));
    LocalMux I__4625 (
            .O(N__21532),
            .I(N__21506));
    LocalMux I__4624 (
            .O(N__21529),
            .I(N__21506));
    InMux I__4623 (
            .O(N__21526),
            .I(N__21503));
    LocalMux I__4622 (
            .O(N__21523),
            .I(N__21500));
    InMux I__4621 (
            .O(N__21520),
            .I(N__21497));
    LocalMux I__4620 (
            .O(N__21517),
            .I(N__21492));
    LocalMux I__4619 (
            .O(N__21514),
            .I(N__21492));
    Span4Mux_h I__4618 (
            .O(N__21511),
            .I(N__21484));
    Span4Mux_v I__4617 (
            .O(N__21506),
            .I(N__21484));
    LocalMux I__4616 (
            .O(N__21503),
            .I(N__21484));
    Span4Mux_h I__4615 (
            .O(N__21500),
            .I(N__21477));
    LocalMux I__4614 (
            .O(N__21497),
            .I(N__21477));
    Span4Mux_s3_v I__4613 (
            .O(N__21492),
            .I(N__21477));
    InMux I__4612 (
            .O(N__21491),
            .I(N__21474));
    Span4Mux_v I__4611 (
            .O(N__21484),
            .I(N__21471));
    Span4Mux_v I__4610 (
            .O(N__21477),
            .I(N__21468));
    LocalMux I__4609 (
            .O(N__21474),
            .I(\tok.S_3 ));
    Odrv4 I__4608 (
            .O(N__21471),
            .I(\tok.S_3 ));
    Odrv4 I__4607 (
            .O(N__21468),
            .I(\tok.S_3 ));
    InMux I__4606 (
            .O(N__21461),
            .I(N__21458));
    LocalMux I__4605 (
            .O(N__21458),
            .I(N__21455));
    Odrv4 I__4604 (
            .O(N__21455),
            .I(\tok.n23_adj_788 ));
    CascadeMux I__4603 (
            .O(N__21452),
            .I(\tok.n10_adj_838_cascade_ ));
    InMux I__4602 (
            .O(N__21449),
            .I(N__21446));
    LocalMux I__4601 (
            .O(N__21446),
            .I(N__21443));
    Odrv4 I__4600 (
            .O(N__21443),
            .I(\tok.n12_adj_840 ));
    InMux I__4599 (
            .O(N__21440),
            .I(N__21437));
    LocalMux I__4598 (
            .O(N__21437),
            .I(N__21431));
    InMux I__4597 (
            .O(N__21436),
            .I(N__21425));
    InMux I__4596 (
            .O(N__21435),
            .I(N__21422));
    InMux I__4595 (
            .O(N__21434),
            .I(N__21419));
    Span4Mux_v I__4594 (
            .O(N__21431),
            .I(N__21416));
    InMux I__4593 (
            .O(N__21430),
            .I(N__21411));
    InMux I__4592 (
            .O(N__21429),
            .I(N__21411));
    InMux I__4591 (
            .O(N__21428),
            .I(N__21407));
    LocalMux I__4590 (
            .O(N__21425),
            .I(N__21404));
    LocalMux I__4589 (
            .O(N__21422),
            .I(N__21397));
    LocalMux I__4588 (
            .O(N__21419),
            .I(N__21394));
    Span4Mux_h I__4587 (
            .O(N__21416),
            .I(N__21389));
    LocalMux I__4586 (
            .O(N__21411),
            .I(N__21389));
    InMux I__4585 (
            .O(N__21410),
            .I(N__21386));
    LocalMux I__4584 (
            .O(N__21407),
            .I(N__21383));
    Span4Mux_h I__4583 (
            .O(N__21404),
            .I(N__21380));
    InMux I__4582 (
            .O(N__21403),
            .I(N__21375));
    InMux I__4581 (
            .O(N__21402),
            .I(N__21375));
    InMux I__4580 (
            .O(N__21401),
            .I(N__21370));
    InMux I__4579 (
            .O(N__21400),
            .I(N__21370));
    Span4Mux_h I__4578 (
            .O(N__21397),
            .I(N__21363));
    Span4Mux_v I__4577 (
            .O(N__21394),
            .I(N__21363));
    Span4Mux_v I__4576 (
            .O(N__21389),
            .I(N__21363));
    LocalMux I__4575 (
            .O(N__21386),
            .I(N__21358));
    Span4Mux_h I__4574 (
            .O(N__21383),
            .I(N__21358));
    Odrv4 I__4573 (
            .O(N__21380),
            .I(\tok.n57 ));
    LocalMux I__4572 (
            .O(N__21375),
            .I(\tok.n57 ));
    LocalMux I__4571 (
            .O(N__21370),
            .I(\tok.n57 ));
    Odrv4 I__4570 (
            .O(N__21363),
            .I(\tok.n57 ));
    Odrv4 I__4569 (
            .O(N__21358),
            .I(\tok.n57 ));
    InMux I__4568 (
            .O(N__21347),
            .I(N__21344));
    LocalMux I__4567 (
            .O(N__21344),
            .I(\tok.n6_adj_835 ));
    InMux I__4566 (
            .O(N__21341),
            .I(N__21337));
    InMux I__4565 (
            .O(N__21340),
            .I(N__21334));
    LocalMux I__4564 (
            .O(N__21337),
            .I(N__21331));
    LocalMux I__4563 (
            .O(N__21334),
            .I(uart_rx_data_6));
    Odrv12 I__4562 (
            .O(N__21331),
            .I(uart_rx_data_6));
    CascadeMux I__4561 (
            .O(N__21326),
            .I(\tok.n109_cascade_ ));
    InMux I__4560 (
            .O(N__21323),
            .I(N__21316));
    CascadeMux I__4559 (
            .O(N__21322),
            .I(N__21313));
    CascadeMux I__4558 (
            .O(N__21321),
            .I(N__21310));
    InMux I__4557 (
            .O(N__21320),
            .I(N__21307));
    InMux I__4556 (
            .O(N__21319),
            .I(N__21304));
    LocalMux I__4555 (
            .O(N__21316),
            .I(N__21300));
    InMux I__4554 (
            .O(N__21313),
            .I(N__21295));
    InMux I__4553 (
            .O(N__21310),
            .I(N__21292));
    LocalMux I__4552 (
            .O(N__21307),
            .I(N__21287));
    LocalMux I__4551 (
            .O(N__21304),
            .I(N__21287));
    CascadeMux I__4550 (
            .O(N__21303),
            .I(N__21284));
    Span4Mux_v I__4549 (
            .O(N__21300),
            .I(N__21281));
    InMux I__4548 (
            .O(N__21299),
            .I(N__21278));
    InMux I__4547 (
            .O(N__21298),
            .I(N__21275));
    LocalMux I__4546 (
            .O(N__21295),
            .I(N__21270));
    LocalMux I__4545 (
            .O(N__21292),
            .I(N__21270));
    Span4Mux_v I__4544 (
            .O(N__21287),
            .I(N__21266));
    InMux I__4543 (
            .O(N__21284),
            .I(N__21263));
    Span4Mux_h I__4542 (
            .O(N__21281),
            .I(N__21258));
    LocalMux I__4541 (
            .O(N__21278),
            .I(N__21258));
    LocalMux I__4540 (
            .O(N__21275),
            .I(N__21253));
    Span4Mux_h I__4539 (
            .O(N__21270),
            .I(N__21253));
    InMux I__4538 (
            .O(N__21269),
            .I(N__21250));
    Sp12to4 I__4537 (
            .O(N__21266),
            .I(N__21245));
    LocalMux I__4536 (
            .O(N__21263),
            .I(N__21245));
    Span4Mux_v I__4535 (
            .O(N__21258),
            .I(N__21240));
    Span4Mux_h I__4534 (
            .O(N__21253),
            .I(N__21240));
    LocalMux I__4533 (
            .O(N__21250),
            .I(\tok.S_6 ));
    Odrv12 I__4532 (
            .O(N__21245),
            .I(\tok.S_6 ));
    Odrv4 I__4531 (
            .O(N__21240),
            .I(\tok.S_6 ));
    InMux I__4530 (
            .O(N__21233),
            .I(N__21230));
    LocalMux I__4529 (
            .O(N__21230),
            .I(N__21227));
    Span4Mux_v I__4528 (
            .O(N__21227),
            .I(N__21224));
    Odrv4 I__4527 (
            .O(N__21224),
            .I(\tok.n18_adj_782 ));
    InMux I__4526 (
            .O(N__21221),
            .I(N__21218));
    LocalMux I__4525 (
            .O(N__21218),
            .I(N__21215));
    Span4Mux_h I__4524 (
            .O(N__21215),
            .I(N__21211));
    InMux I__4523 (
            .O(N__21214),
            .I(N__21208));
    Span4Mux_h I__4522 (
            .O(N__21211),
            .I(N__21202));
    LocalMux I__4521 (
            .O(N__21208),
            .I(N__21202));
    InMux I__4520 (
            .O(N__21207),
            .I(N__21199));
    Odrv4 I__4519 (
            .O(N__21202),
            .I(capture_4));
    LocalMux I__4518 (
            .O(N__21199),
            .I(capture_4));
    CascadeMux I__4517 (
            .O(N__21194),
            .I(N__21190));
    InMux I__4516 (
            .O(N__21193),
            .I(N__21185));
    InMux I__4515 (
            .O(N__21190),
            .I(N__21185));
    LocalMux I__4514 (
            .O(N__21185),
            .I(uart_rx_data_3));
    CascadeMux I__4513 (
            .O(N__21182),
            .I(N__21177));
    InMux I__4512 (
            .O(N__21181),
            .I(N__21174));
    InMux I__4511 (
            .O(N__21180),
            .I(N__21170));
    InMux I__4510 (
            .O(N__21177),
            .I(N__21165));
    LocalMux I__4509 (
            .O(N__21174),
            .I(N__21162));
    InMux I__4508 (
            .O(N__21173),
            .I(N__21159));
    LocalMux I__4507 (
            .O(N__21170),
            .I(N__21155));
    InMux I__4506 (
            .O(N__21169),
            .I(N__21152));
    InMux I__4505 (
            .O(N__21168),
            .I(N__21149));
    LocalMux I__4504 (
            .O(N__21165),
            .I(N__21146));
    Span4Mux_h I__4503 (
            .O(N__21162),
            .I(N__21142));
    LocalMux I__4502 (
            .O(N__21159),
            .I(N__21139));
    InMux I__4501 (
            .O(N__21158),
            .I(N__21136));
    Span4Mux_v I__4500 (
            .O(N__21155),
            .I(N__21129));
    LocalMux I__4499 (
            .O(N__21152),
            .I(N__21129));
    LocalMux I__4498 (
            .O(N__21149),
            .I(N__21129));
    Span4Mux_v I__4497 (
            .O(N__21146),
            .I(N__21126));
    CascadeMux I__4496 (
            .O(N__21145),
            .I(N__21123));
    Span4Mux_s0_h I__4495 (
            .O(N__21142),
            .I(N__21118));
    Span4Mux_h I__4494 (
            .O(N__21139),
            .I(N__21118));
    LocalMux I__4493 (
            .O(N__21136),
            .I(N__21115));
    Span4Mux_v I__4492 (
            .O(N__21129),
            .I(N__21112));
    Span4Mux_h I__4491 (
            .O(N__21126),
            .I(N__21109));
    InMux I__4490 (
            .O(N__21123),
            .I(N__21106));
    Span4Mux_v I__4489 (
            .O(N__21118),
            .I(N__21103));
    Span4Mux_v I__4488 (
            .O(N__21115),
            .I(N__21096));
    Span4Mux_h I__4487 (
            .O(N__21112),
            .I(N__21096));
    Span4Mux_h I__4486 (
            .O(N__21109),
            .I(N__21096));
    LocalMux I__4485 (
            .O(N__21106),
            .I(\tok.S_9 ));
    Odrv4 I__4484 (
            .O(N__21103),
            .I(\tok.S_9 ));
    Odrv4 I__4483 (
            .O(N__21096),
            .I(\tok.S_9 ));
    CascadeMux I__4482 (
            .O(N__21089),
            .I(N__21086));
    InMux I__4481 (
            .O(N__21086),
            .I(N__21083));
    LocalMux I__4480 (
            .O(N__21083),
            .I(N__21080));
    Span4Mux_v I__4479 (
            .O(N__21080),
            .I(N__21077));
    Span4Mux_h I__4478 (
            .O(N__21077),
            .I(N__21074));
    Odrv4 I__4477 (
            .O(N__21074),
            .I(\tok.n21 ));
    InMux I__4476 (
            .O(N__21071),
            .I(\tok.n3933 ));
    InMux I__4475 (
            .O(N__21068),
            .I(N__21064));
    InMux I__4474 (
            .O(N__21067),
            .I(N__21061));
    LocalMux I__4473 (
            .O(N__21064),
            .I(N__21056));
    LocalMux I__4472 (
            .O(N__21061),
            .I(N__21051));
    InMux I__4471 (
            .O(N__21060),
            .I(N__21048));
    InMux I__4470 (
            .O(N__21059),
            .I(N__21044));
    Span4Mux_v I__4469 (
            .O(N__21056),
            .I(N__21041));
    InMux I__4468 (
            .O(N__21055),
            .I(N__21038));
    InMux I__4467 (
            .O(N__21054),
            .I(N__21035));
    Span4Mux_v I__4466 (
            .O(N__21051),
            .I(N__21026));
    LocalMux I__4465 (
            .O(N__21048),
            .I(N__21023));
    InMux I__4464 (
            .O(N__21047),
            .I(N__21020));
    LocalMux I__4463 (
            .O(N__21044),
            .I(N__21017));
    Span4Mux_h I__4462 (
            .O(N__21041),
            .I(N__21012));
    LocalMux I__4461 (
            .O(N__21038),
            .I(N__21012));
    LocalMux I__4460 (
            .O(N__21035),
            .I(N__21009));
    InMux I__4459 (
            .O(N__21034),
            .I(N__21006));
    InMux I__4458 (
            .O(N__21033),
            .I(N__21001));
    InMux I__4457 (
            .O(N__21032),
            .I(N__21001));
    InMux I__4456 (
            .O(N__21031),
            .I(N__20994));
    InMux I__4455 (
            .O(N__21030),
            .I(N__20994));
    InMux I__4454 (
            .O(N__21029),
            .I(N__20994));
    Span4Mux_h I__4453 (
            .O(N__21026),
            .I(N__20987));
    Span4Mux_v I__4452 (
            .O(N__21023),
            .I(N__20987));
    LocalMux I__4451 (
            .O(N__21020),
            .I(N__20987));
    Span4Mux_h I__4450 (
            .O(N__21017),
            .I(N__20982));
    Span4Mux_h I__4449 (
            .O(N__21012),
            .I(N__20982));
    Span4Mux_h I__4448 (
            .O(N__21009),
            .I(N__20977));
    LocalMux I__4447 (
            .O(N__21006),
            .I(N__20977));
    LocalMux I__4446 (
            .O(N__21001),
            .I(\tok.n58 ));
    LocalMux I__4445 (
            .O(N__20994),
            .I(\tok.n58 ));
    Odrv4 I__4444 (
            .O(N__20987),
            .I(\tok.n58 ));
    Odrv4 I__4443 (
            .O(N__20982),
            .I(\tok.n58 ));
    Odrv4 I__4442 (
            .O(N__20977),
            .I(\tok.n58 ));
    CascadeMux I__4441 (
            .O(N__20966),
            .I(N__20962));
    CascadeMux I__4440 (
            .O(N__20965),
            .I(N__20959));
    InMux I__4439 (
            .O(N__20962),
            .I(N__20955));
    InMux I__4438 (
            .O(N__20959),
            .I(N__20949));
    InMux I__4437 (
            .O(N__20958),
            .I(N__20944));
    LocalMux I__4436 (
            .O(N__20955),
            .I(N__20941));
    InMux I__4435 (
            .O(N__20954),
            .I(N__20938));
    InMux I__4434 (
            .O(N__20953),
            .I(N__20935));
    InMux I__4433 (
            .O(N__20952),
            .I(N__20932));
    LocalMux I__4432 (
            .O(N__20949),
            .I(N__20929));
    CascadeMux I__4431 (
            .O(N__20948),
            .I(N__20926));
    InMux I__4430 (
            .O(N__20947),
            .I(N__20923));
    LocalMux I__4429 (
            .O(N__20944),
            .I(N__20918));
    Span4Mux_h I__4428 (
            .O(N__20941),
            .I(N__20918));
    LocalMux I__4427 (
            .O(N__20938),
            .I(N__20913));
    LocalMux I__4426 (
            .O(N__20935),
            .I(N__20913));
    LocalMux I__4425 (
            .O(N__20932),
            .I(N__20908));
    Span4Mux_h I__4424 (
            .O(N__20929),
            .I(N__20908));
    InMux I__4423 (
            .O(N__20926),
            .I(N__20905));
    LocalMux I__4422 (
            .O(N__20923),
            .I(N__20902));
    Span4Mux_v I__4421 (
            .O(N__20918),
            .I(N__20899));
    Span4Mux_h I__4420 (
            .O(N__20913),
            .I(N__20896));
    Span4Mux_h I__4419 (
            .O(N__20908),
            .I(N__20893));
    LocalMux I__4418 (
            .O(N__20905),
            .I(\tok.S_10 ));
    Odrv12 I__4417 (
            .O(N__20902),
            .I(\tok.S_10 ));
    Odrv4 I__4416 (
            .O(N__20899),
            .I(\tok.S_10 ));
    Odrv4 I__4415 (
            .O(N__20896),
            .I(\tok.S_10 ));
    Odrv4 I__4414 (
            .O(N__20893),
            .I(\tok.S_10 ));
    InMux I__4413 (
            .O(N__20882),
            .I(N__20879));
    LocalMux I__4412 (
            .O(N__20879),
            .I(N__20876));
    Odrv4 I__4411 (
            .O(N__20876),
            .I(\tok.n5_adj_668 ));
    InMux I__4410 (
            .O(N__20873),
            .I(\tok.n3934 ));
    InMux I__4409 (
            .O(N__20870),
            .I(N__20864));
    CascadeMux I__4408 (
            .O(N__20869),
            .I(N__20861));
    CascadeMux I__4407 (
            .O(N__20868),
            .I(N__20858));
    InMux I__4406 (
            .O(N__20867),
            .I(N__20854));
    LocalMux I__4405 (
            .O(N__20864),
            .I(N__20850));
    InMux I__4404 (
            .O(N__20861),
            .I(N__20847));
    InMux I__4403 (
            .O(N__20858),
            .I(N__20844));
    InMux I__4402 (
            .O(N__20857),
            .I(N__20839));
    LocalMux I__4401 (
            .O(N__20854),
            .I(N__20836));
    InMux I__4400 (
            .O(N__20853),
            .I(N__20833));
    Span4Mux_s3_v I__4399 (
            .O(N__20850),
            .I(N__20828));
    LocalMux I__4398 (
            .O(N__20847),
            .I(N__20828));
    LocalMux I__4397 (
            .O(N__20844),
            .I(N__20825));
    CascadeMux I__4396 (
            .O(N__20843),
            .I(N__20822));
    InMux I__4395 (
            .O(N__20842),
            .I(N__20819));
    LocalMux I__4394 (
            .O(N__20839),
            .I(N__20816));
    Span4Mux_s3_v I__4393 (
            .O(N__20836),
            .I(N__20811));
    LocalMux I__4392 (
            .O(N__20833),
            .I(N__20811));
    Span4Mux_v I__4391 (
            .O(N__20828),
            .I(N__20808));
    Span4Mux_v I__4390 (
            .O(N__20825),
            .I(N__20805));
    InMux I__4389 (
            .O(N__20822),
            .I(N__20802));
    LocalMux I__4388 (
            .O(N__20819),
            .I(N__20799));
    Span4Mux_h I__4387 (
            .O(N__20816),
            .I(N__20792));
    Span4Mux_v I__4386 (
            .O(N__20811),
            .I(N__20792));
    Span4Mux_h I__4385 (
            .O(N__20808),
            .I(N__20792));
    Span4Mux_h I__4384 (
            .O(N__20805),
            .I(N__20789));
    LocalMux I__4383 (
            .O(N__20802),
            .I(N__20784));
    Span4Mux_v I__4382 (
            .O(N__20799),
            .I(N__20784));
    Span4Mux_h I__4381 (
            .O(N__20792),
            .I(N__20781));
    Odrv4 I__4380 (
            .O(N__20789),
            .I(\tok.S_11 ));
    Odrv4 I__4379 (
            .O(N__20784),
            .I(\tok.S_11 ));
    Odrv4 I__4378 (
            .O(N__20781),
            .I(\tok.S_11 ));
    InMux I__4377 (
            .O(N__20774),
            .I(N__20771));
    LocalMux I__4376 (
            .O(N__20771),
            .I(N__20768));
    Odrv12 I__4375 (
            .O(N__20768),
            .I(\tok.n5_adj_690 ));
    InMux I__4374 (
            .O(N__20765),
            .I(\tok.n3935 ));
    InMux I__4373 (
            .O(N__20762),
            .I(N__20757));
    CascadeMux I__4372 (
            .O(N__20761),
            .I(N__20754));
    CascadeMux I__4371 (
            .O(N__20760),
            .I(N__20748));
    LocalMux I__4370 (
            .O(N__20757),
            .I(N__20745));
    InMux I__4369 (
            .O(N__20754),
            .I(N__20742));
    InMux I__4368 (
            .O(N__20753),
            .I(N__20739));
    InMux I__4367 (
            .O(N__20752),
            .I(N__20736));
    InMux I__4366 (
            .O(N__20751),
            .I(N__20733));
    InMux I__4365 (
            .O(N__20748),
            .I(N__20729));
    Span4Mux_v I__4364 (
            .O(N__20745),
            .I(N__20724));
    LocalMux I__4363 (
            .O(N__20742),
            .I(N__20724));
    LocalMux I__4362 (
            .O(N__20739),
            .I(N__20716));
    LocalMux I__4361 (
            .O(N__20736),
            .I(N__20716));
    LocalMux I__4360 (
            .O(N__20733),
            .I(N__20716));
    InMux I__4359 (
            .O(N__20732),
            .I(N__20713));
    LocalMux I__4358 (
            .O(N__20729),
            .I(N__20710));
    Span4Mux_v I__4357 (
            .O(N__20724),
            .I(N__20707));
    InMux I__4356 (
            .O(N__20723),
            .I(N__20704));
    Span12Mux_v I__4355 (
            .O(N__20716),
            .I(N__20701));
    LocalMux I__4354 (
            .O(N__20713),
            .I(N__20696));
    Span12Mux_s8_h I__4353 (
            .O(N__20710),
            .I(N__20696));
    Span4Mux_v I__4352 (
            .O(N__20707),
            .I(N__20693));
    LocalMux I__4351 (
            .O(N__20704),
            .I(\tok.S_12 ));
    Odrv12 I__4350 (
            .O(N__20701),
            .I(\tok.S_12 ));
    Odrv12 I__4349 (
            .O(N__20696),
            .I(\tok.S_12 ));
    Odrv4 I__4348 (
            .O(N__20693),
            .I(\tok.S_12 ));
    InMux I__4347 (
            .O(N__20684),
            .I(\tok.n3936 ));
    InMux I__4346 (
            .O(N__20681),
            .I(N__20673));
    InMux I__4345 (
            .O(N__20680),
            .I(N__20670));
    InMux I__4344 (
            .O(N__20679),
            .I(N__20667));
    InMux I__4343 (
            .O(N__20678),
            .I(N__20664));
    InMux I__4342 (
            .O(N__20677),
            .I(N__20661));
    InMux I__4341 (
            .O(N__20676),
            .I(N__20658));
    LocalMux I__4340 (
            .O(N__20673),
            .I(N__20653));
    LocalMux I__4339 (
            .O(N__20670),
            .I(N__20653));
    LocalMux I__4338 (
            .O(N__20667),
            .I(N__20647));
    LocalMux I__4337 (
            .O(N__20664),
            .I(N__20647));
    LocalMux I__4336 (
            .O(N__20661),
            .I(N__20644));
    LocalMux I__4335 (
            .O(N__20658),
            .I(N__20638));
    Span4Mux_v I__4334 (
            .O(N__20653),
            .I(N__20635));
    InMux I__4333 (
            .O(N__20652),
            .I(N__20632));
    Span4Mux_v I__4332 (
            .O(N__20647),
            .I(N__20627));
    Span4Mux_h I__4331 (
            .O(N__20644),
            .I(N__20627));
    InMux I__4330 (
            .O(N__20643),
            .I(N__20622));
    InMux I__4329 (
            .O(N__20642),
            .I(N__20622));
    InMux I__4328 (
            .O(N__20641),
            .I(N__20619));
    Span4Mux_h I__4327 (
            .O(N__20638),
            .I(N__20616));
    Span4Mux_v I__4326 (
            .O(N__20635),
            .I(N__20611));
    LocalMux I__4325 (
            .O(N__20632),
            .I(N__20611));
    Span4Mux_v I__4324 (
            .O(N__20627),
            .I(N__20608));
    LocalMux I__4323 (
            .O(N__20622),
            .I(\tok.n55 ));
    LocalMux I__4322 (
            .O(N__20619),
            .I(\tok.n55 ));
    Odrv4 I__4321 (
            .O(N__20616),
            .I(\tok.n55 ));
    Odrv4 I__4320 (
            .O(N__20611),
            .I(\tok.n55 ));
    Odrv4 I__4319 (
            .O(N__20608),
            .I(\tok.n55 ));
    InMux I__4318 (
            .O(N__20597),
            .I(N__20592));
    InMux I__4317 (
            .O(N__20596),
            .I(N__20589));
    CascadeMux I__4316 (
            .O(N__20595),
            .I(N__20584));
    LocalMux I__4315 (
            .O(N__20592),
            .I(N__20580));
    LocalMux I__4314 (
            .O(N__20589),
            .I(N__20577));
    InMux I__4313 (
            .O(N__20588),
            .I(N__20574));
    InMux I__4312 (
            .O(N__20587),
            .I(N__20571));
    InMux I__4311 (
            .O(N__20584),
            .I(N__20568));
    CascadeMux I__4310 (
            .O(N__20583),
            .I(N__20565));
    Span4Mux_v I__4309 (
            .O(N__20580),
            .I(N__20554));
    Span4Mux_s3_h I__4308 (
            .O(N__20577),
            .I(N__20554));
    LocalMux I__4307 (
            .O(N__20574),
            .I(N__20554));
    LocalMux I__4306 (
            .O(N__20571),
            .I(N__20554));
    LocalMux I__4305 (
            .O(N__20568),
            .I(N__20551));
    InMux I__4304 (
            .O(N__20565),
            .I(N__20548));
    CascadeMux I__4303 (
            .O(N__20564),
            .I(N__20545));
    InMux I__4302 (
            .O(N__20563),
            .I(N__20542));
    Span4Mux_h I__4301 (
            .O(N__20554),
            .I(N__20537));
    Span4Mux_h I__4300 (
            .O(N__20551),
            .I(N__20537));
    LocalMux I__4299 (
            .O(N__20548),
            .I(N__20534));
    InMux I__4298 (
            .O(N__20545),
            .I(N__20531));
    LocalMux I__4297 (
            .O(N__20542),
            .I(N__20528));
    Span4Mux_v I__4296 (
            .O(N__20537),
            .I(N__20525));
    Span4Mux_h I__4295 (
            .O(N__20534),
            .I(N__20522));
    LocalMux I__4294 (
            .O(N__20531),
            .I(\tok.S_13 ));
    Odrv12 I__4293 (
            .O(N__20528),
            .I(\tok.S_13 ));
    Odrv4 I__4292 (
            .O(N__20525),
            .I(\tok.S_13 ));
    Odrv4 I__4291 (
            .O(N__20522),
            .I(\tok.S_13 ));
    InMux I__4290 (
            .O(N__20513),
            .I(\tok.n3937 ));
    InMux I__4289 (
            .O(N__20510),
            .I(N__20502));
    InMux I__4288 (
            .O(N__20509),
            .I(N__20499));
    CascadeMux I__4287 (
            .O(N__20508),
            .I(N__20496));
    InMux I__4286 (
            .O(N__20507),
            .I(N__20492));
    InMux I__4285 (
            .O(N__20506),
            .I(N__20489));
    InMux I__4284 (
            .O(N__20505),
            .I(N__20486));
    LocalMux I__4283 (
            .O(N__20502),
            .I(N__20483));
    LocalMux I__4282 (
            .O(N__20499),
            .I(N__20480));
    InMux I__4281 (
            .O(N__20496),
            .I(N__20477));
    InMux I__4280 (
            .O(N__20495),
            .I(N__20474));
    LocalMux I__4279 (
            .O(N__20492),
            .I(N__20471));
    LocalMux I__4278 (
            .O(N__20489),
            .I(N__20468));
    LocalMux I__4277 (
            .O(N__20486),
            .I(N__20465));
    Span4Mux_h I__4276 (
            .O(N__20483),
            .I(N__20462));
    Span4Mux_v I__4275 (
            .O(N__20480),
            .I(N__20457));
    LocalMux I__4274 (
            .O(N__20477),
            .I(N__20457));
    LocalMux I__4273 (
            .O(N__20474),
            .I(N__20453));
    Span4Mux_v I__4272 (
            .O(N__20471),
            .I(N__20450));
    Span4Mux_v I__4271 (
            .O(N__20468),
            .I(N__20445));
    Span4Mux_v I__4270 (
            .O(N__20465),
            .I(N__20445));
    Span4Mux_v I__4269 (
            .O(N__20462),
            .I(N__20442));
    Span4Mux_h I__4268 (
            .O(N__20457),
            .I(N__20439));
    InMux I__4267 (
            .O(N__20456),
            .I(N__20436));
    Span4Mux_v I__4266 (
            .O(N__20453),
            .I(N__20433));
    Span4Mux_v I__4265 (
            .O(N__20450),
            .I(N__20428));
    Span4Mux_v I__4264 (
            .O(N__20445),
            .I(N__20428));
    Span4Mux_h I__4263 (
            .O(N__20442),
            .I(N__20425));
    Span4Mux_h I__4262 (
            .O(N__20439),
            .I(N__20422));
    LocalMux I__4261 (
            .O(N__20436),
            .I(\tok.S_14 ));
    Odrv4 I__4260 (
            .O(N__20433),
            .I(\tok.S_14 ));
    Odrv4 I__4259 (
            .O(N__20428),
            .I(\tok.S_14 ));
    Odrv4 I__4258 (
            .O(N__20425),
            .I(\tok.S_14 ));
    Odrv4 I__4257 (
            .O(N__20422),
            .I(\tok.S_14 ));
    InMux I__4256 (
            .O(N__20411),
            .I(N__20408));
    LocalMux I__4255 (
            .O(N__20408),
            .I(\tok.n5_adj_729 ));
    InMux I__4254 (
            .O(N__20405),
            .I(\tok.n3938 ));
    InMux I__4253 (
            .O(N__20402),
            .I(N__20396));
    InMux I__4252 (
            .O(N__20401),
            .I(N__20391));
    CascadeMux I__4251 (
            .O(N__20400),
            .I(N__20388));
    InMux I__4250 (
            .O(N__20399),
            .I(N__20385));
    LocalMux I__4249 (
            .O(N__20396),
            .I(N__20382));
    InMux I__4248 (
            .O(N__20395),
            .I(N__20379));
    InMux I__4247 (
            .O(N__20394),
            .I(N__20376));
    LocalMux I__4246 (
            .O(N__20391),
            .I(N__20373));
    InMux I__4245 (
            .O(N__20388),
            .I(N__20370));
    LocalMux I__4244 (
            .O(N__20385),
            .I(N__20365));
    Span4Mux_v I__4243 (
            .O(N__20382),
            .I(N__20362));
    LocalMux I__4242 (
            .O(N__20379),
            .I(N__20353));
    LocalMux I__4241 (
            .O(N__20376),
            .I(N__20353));
    Span4Mux_v I__4240 (
            .O(N__20373),
            .I(N__20353));
    LocalMux I__4239 (
            .O(N__20370),
            .I(N__20353));
    CascadeMux I__4238 (
            .O(N__20369),
            .I(N__20350));
    InMux I__4237 (
            .O(N__20368),
            .I(N__20347));
    Span4Mux_v I__4236 (
            .O(N__20365),
            .I(N__20344));
    Span4Mux_h I__4235 (
            .O(N__20362),
            .I(N__20339));
    Span4Mux_v I__4234 (
            .O(N__20353),
            .I(N__20339));
    InMux I__4233 (
            .O(N__20350),
            .I(N__20336));
    LocalMux I__4232 (
            .O(N__20347),
            .I(N__20333));
    Span4Mux_v I__4231 (
            .O(N__20344),
            .I(N__20328));
    Span4Mux_v I__4230 (
            .O(N__20339),
            .I(N__20328));
    LocalMux I__4229 (
            .O(N__20336),
            .I(\tok.S_15 ));
    Odrv12 I__4228 (
            .O(N__20333),
            .I(\tok.S_15 ));
    Odrv4 I__4227 (
            .O(N__20328),
            .I(\tok.S_15 ));
    CascadeMux I__4226 (
            .O(N__20321),
            .I(N__20318));
    InMux I__4225 (
            .O(N__20318),
            .I(N__20315));
    LocalMux I__4224 (
            .O(N__20315),
            .I(N__20306));
    InMux I__4223 (
            .O(N__20314),
            .I(N__20302));
    InMux I__4222 (
            .O(N__20313),
            .I(N__20297));
    InMux I__4221 (
            .O(N__20312),
            .I(N__20297));
    CascadeMux I__4220 (
            .O(N__20311),
            .I(N__20294));
    InMux I__4219 (
            .O(N__20310),
            .I(N__20291));
    CascadeMux I__4218 (
            .O(N__20309),
            .I(N__20288));
    Span4Mux_v I__4217 (
            .O(N__20306),
            .I(N__20284));
    InMux I__4216 (
            .O(N__20305),
            .I(N__20281));
    LocalMux I__4215 (
            .O(N__20302),
            .I(N__20277));
    LocalMux I__4214 (
            .O(N__20297),
            .I(N__20274));
    InMux I__4213 (
            .O(N__20294),
            .I(N__20271));
    LocalMux I__4212 (
            .O(N__20291),
            .I(N__20268));
    InMux I__4211 (
            .O(N__20288),
            .I(N__20265));
    CascadeMux I__4210 (
            .O(N__20287),
            .I(N__20262));
    Span4Mux_s3_h I__4209 (
            .O(N__20284),
            .I(N__20259));
    LocalMux I__4208 (
            .O(N__20281),
            .I(N__20256));
    InMux I__4207 (
            .O(N__20280),
            .I(N__20253));
    Span4Mux_v I__4206 (
            .O(N__20277),
            .I(N__20246));
    Span4Mux_s3_h I__4205 (
            .O(N__20274),
            .I(N__20246));
    LocalMux I__4204 (
            .O(N__20271),
            .I(N__20246));
    Span4Mux_s3_v I__4203 (
            .O(N__20268),
            .I(N__20241));
    LocalMux I__4202 (
            .O(N__20265),
            .I(N__20241));
    InMux I__4201 (
            .O(N__20262),
            .I(N__20238));
    Span4Mux_h I__4200 (
            .O(N__20259),
            .I(N__20235));
    Span4Mux_v I__4199 (
            .O(N__20256),
            .I(N__20230));
    LocalMux I__4198 (
            .O(N__20253),
            .I(N__20230));
    Span4Mux_h I__4197 (
            .O(N__20246),
            .I(N__20225));
    Span4Mux_v I__4196 (
            .O(N__20241),
            .I(N__20225));
    LocalMux I__4195 (
            .O(N__20238),
            .I(\tok.n53 ));
    Odrv4 I__4194 (
            .O(N__20235),
            .I(\tok.n53 ));
    Odrv4 I__4193 (
            .O(N__20230),
            .I(\tok.n53 ));
    Odrv4 I__4192 (
            .O(N__20225),
            .I(\tok.n53 ));
    InMux I__4191 (
            .O(N__20216),
            .I(\tok.n3939 ));
    InMux I__4190 (
            .O(N__20213),
            .I(N__20210));
    LocalMux I__4189 (
            .O(N__20210),
            .I(N__20207));
    Span4Mux_v I__4188 (
            .O(N__20207),
            .I(N__20204));
    Sp12to4 I__4187 (
            .O(N__20204),
            .I(N__20201));
    Odrv12 I__4186 (
            .O(N__20201),
            .I(\tok.n5_adj_750 ));
    InMux I__4185 (
            .O(N__20198),
            .I(N__20195));
    LocalMux I__4184 (
            .O(N__20195),
            .I(N__20192));
    Span4Mux_v I__4183 (
            .O(N__20192),
            .I(N__20189));
    Span4Mux_h I__4182 (
            .O(N__20189),
            .I(N__20186));
    Odrv4 I__4181 (
            .O(N__20186),
            .I(\tok.n6_adj_812 ));
    InMux I__4180 (
            .O(N__20183),
            .I(N__20180));
    LocalMux I__4179 (
            .O(N__20180),
            .I(N__20177));
    Span12Mux_s10_v I__4178 (
            .O(N__20177),
            .I(N__20174));
    Odrv12 I__4177 (
            .O(N__20174),
            .I(\tok.n9_adj_836 ));
    CascadeMux I__4176 (
            .O(N__20171),
            .I(N__20166));
    CascadeMux I__4175 (
            .O(N__20170),
            .I(N__20163));
    CascadeMux I__4174 (
            .O(N__20169),
            .I(N__20159));
    InMux I__4173 (
            .O(N__20166),
            .I(N__20156));
    InMux I__4172 (
            .O(N__20163),
            .I(N__20151));
    InMux I__4171 (
            .O(N__20162),
            .I(N__20147));
    InMux I__4170 (
            .O(N__20159),
            .I(N__20144));
    LocalMux I__4169 (
            .O(N__20156),
            .I(N__20140));
    InMux I__4168 (
            .O(N__20155),
            .I(N__20137));
    InMux I__4167 (
            .O(N__20154),
            .I(N__20134));
    LocalMux I__4166 (
            .O(N__20151),
            .I(N__20131));
    InMux I__4165 (
            .O(N__20150),
            .I(N__20128));
    LocalMux I__4164 (
            .O(N__20147),
            .I(N__20123));
    LocalMux I__4163 (
            .O(N__20144),
            .I(N__20123));
    InMux I__4162 (
            .O(N__20143),
            .I(N__20120));
    Span4Mux_v I__4161 (
            .O(N__20140),
            .I(N__20117));
    LocalMux I__4160 (
            .O(N__20137),
            .I(N__20114));
    LocalMux I__4159 (
            .O(N__20134),
            .I(N__20106));
    Span4Mux_v I__4158 (
            .O(N__20131),
            .I(N__20106));
    LocalMux I__4157 (
            .O(N__20128),
            .I(N__20106));
    Span4Mux_v I__4156 (
            .O(N__20123),
            .I(N__20101));
    LocalMux I__4155 (
            .O(N__20120),
            .I(N__20101));
    Span4Mux_h I__4154 (
            .O(N__20117),
            .I(N__20098));
    Span4Mux_v I__4153 (
            .O(N__20114),
            .I(N__20095));
    InMux I__4152 (
            .O(N__20113),
            .I(N__20092));
    Span4Mux_v I__4151 (
            .O(N__20106),
            .I(N__20087));
    Span4Mux_h I__4150 (
            .O(N__20101),
            .I(N__20087));
    Odrv4 I__4149 (
            .O(N__20098),
            .I(\tok.S_1 ));
    Odrv4 I__4148 (
            .O(N__20095),
            .I(\tok.S_1 ));
    LocalMux I__4147 (
            .O(N__20092),
            .I(\tok.S_1 ));
    Odrv4 I__4146 (
            .O(N__20087),
            .I(\tok.S_1 ));
    InMux I__4145 (
            .O(N__20078),
            .I(N__20075));
    LocalMux I__4144 (
            .O(N__20075),
            .I(\tok.n4_adj_790 ));
    InMux I__4143 (
            .O(N__20072),
            .I(\tok.n3925 ));
    CascadeMux I__4142 (
            .O(N__20069),
            .I(N__20065));
    CascadeMux I__4141 (
            .O(N__20068),
            .I(N__20061));
    InMux I__4140 (
            .O(N__20065),
            .I(N__20056));
    CascadeMux I__4139 (
            .O(N__20064),
            .I(N__20053));
    InMux I__4138 (
            .O(N__20061),
            .I(N__20050));
    CascadeMux I__4137 (
            .O(N__20060),
            .I(N__20047));
    InMux I__4136 (
            .O(N__20059),
            .I(N__20044));
    LocalMux I__4135 (
            .O(N__20056),
            .I(N__20039));
    InMux I__4134 (
            .O(N__20053),
            .I(N__20036));
    LocalMux I__4133 (
            .O(N__20050),
            .I(N__20032));
    InMux I__4132 (
            .O(N__20047),
            .I(N__20029));
    LocalMux I__4131 (
            .O(N__20044),
            .I(N__20025));
    InMux I__4130 (
            .O(N__20043),
            .I(N__20020));
    InMux I__4129 (
            .O(N__20042),
            .I(N__20020));
    Span4Mux_h I__4128 (
            .O(N__20039),
            .I(N__20017));
    LocalMux I__4127 (
            .O(N__20036),
            .I(N__20014));
    InMux I__4126 (
            .O(N__20035),
            .I(N__20011));
    Span4Mux_h I__4125 (
            .O(N__20032),
            .I(N__20006));
    LocalMux I__4124 (
            .O(N__20029),
            .I(N__20006));
    CascadeMux I__4123 (
            .O(N__20028),
            .I(N__20003));
    Span4Mux_h I__4122 (
            .O(N__20025),
            .I(N__19998));
    LocalMux I__4121 (
            .O(N__20020),
            .I(N__19998));
    Span4Mux_h I__4120 (
            .O(N__20017),
            .I(N__19991));
    Span4Mux_v I__4119 (
            .O(N__20014),
            .I(N__19991));
    LocalMux I__4118 (
            .O(N__20011),
            .I(N__19991));
    Span4Mux_v I__4117 (
            .O(N__20006),
            .I(N__19988));
    InMux I__4116 (
            .O(N__20003),
            .I(N__19985));
    Span4Mux_v I__4115 (
            .O(N__19998),
            .I(N__19982));
    Span4Mux_v I__4114 (
            .O(N__19991),
            .I(N__19977));
    Span4Mux_h I__4113 (
            .O(N__19988),
            .I(N__19977));
    LocalMux I__4112 (
            .O(N__19985),
            .I(\tok.S_2 ));
    Odrv4 I__4111 (
            .O(N__19982),
            .I(\tok.S_2 ));
    Odrv4 I__4110 (
            .O(N__19977),
            .I(\tok.S_2 ));
    CascadeMux I__4109 (
            .O(N__19970),
            .I(N__19967));
    InMux I__4108 (
            .O(N__19967),
            .I(N__19964));
    LocalMux I__4107 (
            .O(N__19964),
            .I(\tok.n5_adj_789 ));
    InMux I__4106 (
            .O(N__19961),
            .I(\tok.n3926 ));
    InMux I__4105 (
            .O(N__19958),
            .I(\tok.n3927 ));
    InMux I__4104 (
            .O(N__19955),
            .I(\tok.n3928 ));
    CascadeMux I__4103 (
            .O(N__19952),
            .I(N__19943));
    CascadeMux I__4102 (
            .O(N__19951),
            .I(N__19940));
    CascadeMux I__4101 (
            .O(N__19950),
            .I(N__19937));
    CascadeMux I__4100 (
            .O(N__19949),
            .I(N__19934));
    InMux I__4099 (
            .O(N__19948),
            .I(N__19929));
    InMux I__4098 (
            .O(N__19947),
            .I(N__19929));
    CascadeMux I__4097 (
            .O(N__19946),
            .I(N__19926));
    InMux I__4096 (
            .O(N__19943),
            .I(N__19923));
    InMux I__4095 (
            .O(N__19940),
            .I(N__19920));
    InMux I__4094 (
            .O(N__19937),
            .I(N__19916));
    InMux I__4093 (
            .O(N__19934),
            .I(N__19913));
    LocalMux I__4092 (
            .O(N__19929),
            .I(N__19910));
    InMux I__4091 (
            .O(N__19926),
            .I(N__19907));
    LocalMux I__4090 (
            .O(N__19923),
            .I(N__19901));
    LocalMux I__4089 (
            .O(N__19920),
            .I(N__19901));
    CascadeMux I__4088 (
            .O(N__19919),
            .I(N__19898));
    LocalMux I__4087 (
            .O(N__19916),
            .I(N__19893));
    LocalMux I__4086 (
            .O(N__19913),
            .I(N__19893));
    Span4Mux_h I__4085 (
            .O(N__19910),
            .I(N__19888));
    LocalMux I__4084 (
            .O(N__19907),
            .I(N__19888));
    InMux I__4083 (
            .O(N__19906),
            .I(N__19885));
    Span4Mux_h I__4082 (
            .O(N__19901),
            .I(N__19882));
    InMux I__4081 (
            .O(N__19898),
            .I(N__19879));
    Span12Mux_s9_v I__4080 (
            .O(N__19893),
            .I(N__19876));
    Span4Mux_v I__4079 (
            .O(N__19888),
            .I(N__19869));
    LocalMux I__4078 (
            .O(N__19885),
            .I(N__19869));
    Span4Mux_h I__4077 (
            .O(N__19882),
            .I(N__19869));
    LocalMux I__4076 (
            .O(N__19879),
            .I(\tok.S_5 ));
    Odrv12 I__4075 (
            .O(N__19876),
            .I(\tok.S_5 ));
    Odrv4 I__4074 (
            .O(N__19869),
            .I(\tok.S_5 ));
    CascadeMux I__4073 (
            .O(N__19862),
            .I(N__19859));
    InMux I__4072 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__4071 (
            .O(N__19856),
            .I(N__19853));
    Sp12to4 I__4070 (
            .O(N__19853),
            .I(N__19850));
    Span12Mux_s6_v I__4069 (
            .O(N__19850),
            .I(N__19847));
    Odrv12 I__4068 (
            .O(N__19847),
            .I(\tok.n5_adj_775 ));
    InMux I__4067 (
            .O(N__19844),
            .I(\tok.n3929 ));
    InMux I__4066 (
            .O(N__19841),
            .I(N__19838));
    LocalMux I__4065 (
            .O(N__19838),
            .I(N__19835));
    Span12Mux_s6_v I__4064 (
            .O(N__19835),
            .I(N__19832));
    Odrv12 I__4063 (
            .O(N__19832),
            .I(\tok.n5_adj_773 ));
    InMux I__4062 (
            .O(N__19829),
            .I(\tok.n3930 ));
    InMux I__4061 (
            .O(N__19826),
            .I(N__19821));
    CascadeMux I__4060 (
            .O(N__19825),
            .I(N__19818));
    InMux I__4059 (
            .O(N__19824),
            .I(N__19814));
    LocalMux I__4058 (
            .O(N__19821),
            .I(N__19808));
    InMux I__4057 (
            .O(N__19818),
            .I(N__19803));
    InMux I__4056 (
            .O(N__19817),
            .I(N__19800));
    LocalMux I__4055 (
            .O(N__19814),
            .I(N__19797));
    InMux I__4054 (
            .O(N__19813),
            .I(N__19794));
    CascadeMux I__4053 (
            .O(N__19812),
            .I(N__19791));
    InMux I__4052 (
            .O(N__19811),
            .I(N__19787));
    Span4Mux_h I__4051 (
            .O(N__19808),
            .I(N__19784));
    InMux I__4050 (
            .O(N__19807),
            .I(N__19779));
    InMux I__4049 (
            .O(N__19806),
            .I(N__19779));
    LocalMux I__4048 (
            .O(N__19803),
            .I(N__19776));
    LocalMux I__4047 (
            .O(N__19800),
            .I(N__19771));
    Span4Mux_s3_h I__4046 (
            .O(N__19797),
            .I(N__19766));
    LocalMux I__4045 (
            .O(N__19794),
            .I(N__19766));
    InMux I__4044 (
            .O(N__19791),
            .I(N__19763));
    CascadeMux I__4043 (
            .O(N__19790),
            .I(N__19758));
    LocalMux I__4042 (
            .O(N__19787),
            .I(N__19754));
    Span4Mux_s2_v I__4041 (
            .O(N__19784),
            .I(N__19749));
    LocalMux I__4040 (
            .O(N__19779),
            .I(N__19749));
    Span4Mux_h I__4039 (
            .O(N__19776),
            .I(N__19746));
    InMux I__4038 (
            .O(N__19775),
            .I(N__19743));
    InMux I__4037 (
            .O(N__19774),
            .I(N__19740));
    Span4Mux_s3_v I__4036 (
            .O(N__19771),
            .I(N__19737));
    Span4Mux_h I__4035 (
            .O(N__19766),
            .I(N__19732));
    LocalMux I__4034 (
            .O(N__19763),
            .I(N__19732));
    InMux I__4033 (
            .O(N__19762),
            .I(N__19729));
    InMux I__4032 (
            .O(N__19761),
            .I(N__19722));
    InMux I__4031 (
            .O(N__19758),
            .I(N__19722));
    InMux I__4030 (
            .O(N__19757),
            .I(N__19722));
    Span4Mux_v I__4029 (
            .O(N__19754),
            .I(N__19717));
    Span4Mux_v I__4028 (
            .O(N__19749),
            .I(N__19717));
    Span4Mux_h I__4027 (
            .O(N__19746),
            .I(N__19714));
    LocalMux I__4026 (
            .O(N__19743),
            .I(N__19709));
    LocalMux I__4025 (
            .O(N__19740),
            .I(N__19709));
    Span4Mux_h I__4024 (
            .O(N__19737),
            .I(N__19704));
    Span4Mux_h I__4023 (
            .O(N__19732),
            .I(N__19704));
    LocalMux I__4022 (
            .O(N__19729),
            .I(\tok.A_low_7 ));
    LocalMux I__4021 (
            .O(N__19722),
            .I(\tok.A_low_7 ));
    Odrv4 I__4020 (
            .O(N__19717),
            .I(\tok.A_low_7 ));
    Odrv4 I__4019 (
            .O(N__19714),
            .I(\tok.A_low_7 ));
    Odrv12 I__4018 (
            .O(N__19709),
            .I(\tok.A_low_7 ));
    Odrv4 I__4017 (
            .O(N__19704),
            .I(\tok.A_low_7 ));
    CascadeMux I__4016 (
            .O(N__19691),
            .I(N__19686));
    CascadeMux I__4015 (
            .O(N__19690),
            .I(N__19683));
    CascadeMux I__4014 (
            .O(N__19689),
            .I(N__19680));
    InMux I__4013 (
            .O(N__19686),
            .I(N__19675));
    InMux I__4012 (
            .O(N__19683),
            .I(N__19670));
    InMux I__4011 (
            .O(N__19680),
            .I(N__19667));
    InMux I__4010 (
            .O(N__19679),
            .I(N__19664));
    CascadeMux I__4009 (
            .O(N__19678),
            .I(N__19661));
    LocalMux I__4008 (
            .O(N__19675),
            .I(N__19657));
    InMux I__4007 (
            .O(N__19674),
            .I(N__19652));
    InMux I__4006 (
            .O(N__19673),
            .I(N__19652));
    LocalMux I__4005 (
            .O(N__19670),
            .I(N__19649));
    LocalMux I__4004 (
            .O(N__19667),
            .I(N__19643));
    LocalMux I__4003 (
            .O(N__19664),
            .I(N__19643));
    InMux I__4002 (
            .O(N__19661),
            .I(N__19640));
    CascadeMux I__4001 (
            .O(N__19660),
            .I(N__19637));
    Span4Mux_v I__4000 (
            .O(N__19657),
            .I(N__19631));
    LocalMux I__3999 (
            .O(N__19652),
            .I(N__19631));
    Span4Mux_v I__3998 (
            .O(N__19649),
            .I(N__19628));
    InMux I__3997 (
            .O(N__19648),
            .I(N__19625));
    Span4Mux_v I__3996 (
            .O(N__19643),
            .I(N__19622));
    LocalMux I__3995 (
            .O(N__19640),
            .I(N__19619));
    InMux I__3994 (
            .O(N__19637),
            .I(N__19616));
    InMux I__3993 (
            .O(N__19636),
            .I(N__19613));
    Span4Mux_h I__3992 (
            .O(N__19631),
            .I(N__19610));
    Sp12to4 I__3991 (
            .O(N__19628),
            .I(N__19599));
    LocalMux I__3990 (
            .O(N__19625),
            .I(N__19599));
    Sp12to4 I__3989 (
            .O(N__19622),
            .I(N__19599));
    Span12Mux_s7_v I__3988 (
            .O(N__19619),
            .I(N__19599));
    LocalMux I__3987 (
            .O(N__19616),
            .I(N__19599));
    LocalMux I__3986 (
            .O(N__19613),
            .I(\tok.S_7 ));
    Odrv4 I__3985 (
            .O(N__19610),
            .I(\tok.S_7 ));
    Odrv12 I__3984 (
            .O(N__19599),
            .I(\tok.S_7 ));
    CascadeMux I__3983 (
            .O(N__19592),
            .I(N__19589));
    InMux I__3982 (
            .O(N__19589),
            .I(N__19586));
    LocalMux I__3981 (
            .O(N__19586),
            .I(N__19583));
    Span4Mux_v I__3980 (
            .O(N__19583),
            .I(N__19580));
    Span4Mux_h I__3979 (
            .O(N__19580),
            .I(N__19577));
    Odrv4 I__3978 (
            .O(N__19577),
            .I(\tok.n5_adj_752 ));
    InMux I__3977 (
            .O(N__19574),
            .I(\tok.n3931 ));
    CascadeMux I__3976 (
            .O(N__19571),
            .I(N__19567));
    InMux I__3975 (
            .O(N__19570),
            .I(N__19564));
    InMux I__3974 (
            .O(N__19567),
            .I(N__19559));
    LocalMux I__3973 (
            .O(N__19564),
            .I(N__19556));
    InMux I__3972 (
            .O(N__19563),
            .I(N__19550));
    InMux I__3971 (
            .O(N__19562),
            .I(N__19546));
    LocalMux I__3970 (
            .O(N__19559),
            .I(N__19541));
    Span4Mux_v I__3969 (
            .O(N__19556),
            .I(N__19541));
    InMux I__3968 (
            .O(N__19555),
            .I(N__19538));
    CascadeMux I__3967 (
            .O(N__19554),
            .I(N__19535));
    InMux I__3966 (
            .O(N__19553),
            .I(N__19532));
    LocalMux I__3965 (
            .O(N__19550),
            .I(N__19529));
    InMux I__3964 (
            .O(N__19549),
            .I(N__19526));
    LocalMux I__3963 (
            .O(N__19546),
            .I(N__19523));
    Span4Mux_v I__3962 (
            .O(N__19541),
            .I(N__19518));
    LocalMux I__3961 (
            .O(N__19538),
            .I(N__19518));
    InMux I__3960 (
            .O(N__19535),
            .I(N__19515));
    LocalMux I__3959 (
            .O(N__19532),
            .I(N__19512));
    Span4Mux_v I__3958 (
            .O(N__19529),
            .I(N__19507));
    LocalMux I__3957 (
            .O(N__19526),
            .I(N__19507));
    Span4Mux_v I__3956 (
            .O(N__19523),
            .I(N__19504));
    Span4Mux_h I__3955 (
            .O(N__19518),
            .I(N__19501));
    LocalMux I__3954 (
            .O(N__19515),
            .I(N__19492));
    Span4Mux_v I__3953 (
            .O(N__19512),
            .I(N__19492));
    Span4Mux_v I__3952 (
            .O(N__19507),
            .I(N__19492));
    Span4Mux_h I__3951 (
            .O(N__19504),
            .I(N__19492));
    Odrv4 I__3950 (
            .O(N__19501),
            .I(\tok.S_8 ));
    Odrv4 I__3949 (
            .O(N__19492),
            .I(\tok.S_8 ));
    InMux I__3948 (
            .O(N__19487),
            .I(bfn_9_9_0_));
    InMux I__3947 (
            .O(N__19484),
            .I(N__19481));
    LocalMux I__3946 (
            .O(N__19481),
            .I(N__19477));
    InMux I__3945 (
            .O(N__19480),
            .I(N__19474));
    Odrv4 I__3944 (
            .O(N__19477),
            .I(n10_adj_875));
    LocalMux I__3943 (
            .O(N__19474),
            .I(n10_adj_875));
    CascadeMux I__3942 (
            .O(N__19469),
            .I(N__19465));
    InMux I__3941 (
            .O(N__19468),
            .I(N__19462));
    InMux I__3940 (
            .O(N__19465),
            .I(N__19458));
    LocalMux I__3939 (
            .O(N__19462),
            .I(N__19455));
    InMux I__3938 (
            .O(N__19461),
            .I(N__19451));
    LocalMux I__3937 (
            .O(N__19458),
            .I(N__19448));
    Span4Mux_v I__3936 (
            .O(N__19455),
            .I(N__19445));
    InMux I__3935 (
            .O(N__19454),
            .I(N__19442));
    LocalMux I__3934 (
            .O(N__19451),
            .I(c_stk_w_7_N_18_0));
    Odrv12 I__3933 (
            .O(N__19448),
            .I(c_stk_w_7_N_18_0));
    Odrv4 I__3932 (
            .O(N__19445),
            .I(c_stk_w_7_N_18_0));
    LocalMux I__3931 (
            .O(N__19442),
            .I(c_stk_w_7_N_18_0));
    CascadeMux I__3930 (
            .O(N__19433),
            .I(N__19427));
    CascadeMux I__3929 (
            .O(N__19432),
            .I(N__19424));
    CascadeMux I__3928 (
            .O(N__19431),
            .I(N__19421));
    CascadeMux I__3927 (
            .O(N__19430),
            .I(N__19418));
    InMux I__3926 (
            .O(N__19427),
            .I(N__19409));
    InMux I__3925 (
            .O(N__19424),
            .I(N__19409));
    InMux I__3924 (
            .O(N__19421),
            .I(N__19409));
    InMux I__3923 (
            .O(N__19418),
            .I(N__19409));
    LocalMux I__3922 (
            .O(N__19409),
            .I(N__19402));
    CascadeMux I__3921 (
            .O(N__19408),
            .I(N__19399));
    CascadeMux I__3920 (
            .O(N__19407),
            .I(N__19396));
    CascadeMux I__3919 (
            .O(N__19406),
            .I(N__19393));
    CascadeMux I__3918 (
            .O(N__19405),
            .I(N__19390));
    Span4Mux_v I__3917 (
            .O(N__19402),
            .I(N__19387));
    InMux I__3916 (
            .O(N__19399),
            .I(N__19378));
    InMux I__3915 (
            .O(N__19396),
            .I(N__19378));
    InMux I__3914 (
            .O(N__19393),
            .I(N__19378));
    InMux I__3913 (
            .O(N__19390),
            .I(N__19378));
    Span4Mux_s0_v I__3912 (
            .O(N__19387),
            .I(N__19372));
    LocalMux I__3911 (
            .O(N__19378),
            .I(N__19372));
    InMux I__3910 (
            .O(N__19377),
            .I(N__19368));
    Span4Mux_v I__3909 (
            .O(N__19372),
            .I(N__19365));
    InMux I__3908 (
            .O(N__19371),
            .I(N__19362));
    LocalMux I__3907 (
            .O(N__19368),
            .I(N__19359));
    Span4Mux_h I__3906 (
            .O(N__19365),
            .I(N__19356));
    LocalMux I__3905 (
            .O(N__19362),
            .I(\tok.found_slot ));
    Odrv12 I__3904 (
            .O(N__19359),
            .I(\tok.found_slot ));
    Odrv4 I__3903 (
            .O(N__19356),
            .I(\tok.found_slot ));
    CascadeMux I__3902 (
            .O(N__19349),
            .I(\tok.n5_adj_655_cascade_ ));
    InMux I__3901 (
            .O(N__19346),
            .I(N__19340));
    InMux I__3900 (
            .O(N__19345),
            .I(N__19333));
    InMux I__3899 (
            .O(N__19344),
            .I(N__19333));
    InMux I__3898 (
            .O(N__19343),
            .I(N__19333));
    LocalMux I__3897 (
            .O(N__19340),
            .I(N__19330));
    LocalMux I__3896 (
            .O(N__19333),
            .I(N__19327));
    Span4Mux_h I__3895 (
            .O(N__19330),
            .I(N__19324));
    Span4Mux_h I__3894 (
            .O(N__19327),
            .I(N__19321));
    Span4Mux_h I__3893 (
            .O(N__19324),
            .I(N__19318));
    Odrv4 I__3892 (
            .O(N__19321),
            .I(\tok.uart_tx_busy ));
    Odrv4 I__3891 (
            .O(N__19318),
            .I(\tok.uart_tx_busy ));
    CascadeMux I__3890 (
            .O(N__19313),
            .I(N__19309));
    CascadeMux I__3889 (
            .O(N__19312),
            .I(N__19306));
    InMux I__3888 (
            .O(N__19309),
            .I(N__19303));
    InMux I__3887 (
            .O(N__19306),
            .I(N__19300));
    LocalMux I__3886 (
            .O(N__19303),
            .I(N__19294));
    LocalMux I__3885 (
            .O(N__19300),
            .I(N__19294));
    InMux I__3884 (
            .O(N__19299),
            .I(N__19291));
    Span4Mux_h I__3883 (
            .O(N__19294),
            .I(N__19288));
    LocalMux I__3882 (
            .O(N__19291),
            .I(\tok.uart_rx_valid ));
    Odrv4 I__3881 (
            .O(N__19288),
            .I(\tok.uart_rx_valid ));
    CascadeMux I__3880 (
            .O(N__19283),
            .I(\tok.uart_stall_cascade_ ));
    InMux I__3879 (
            .O(N__19280),
            .I(N__19270));
    InMux I__3878 (
            .O(N__19279),
            .I(N__19270));
    InMux I__3877 (
            .O(N__19278),
            .I(N__19261));
    InMux I__3876 (
            .O(N__19277),
            .I(N__19261));
    InMux I__3875 (
            .O(N__19276),
            .I(N__19261));
    InMux I__3874 (
            .O(N__19275),
            .I(N__19261));
    LocalMux I__3873 (
            .O(N__19270),
            .I(N__19257));
    LocalMux I__3872 (
            .O(N__19261),
            .I(N__19254));
    InMux I__3871 (
            .O(N__19260),
            .I(N__19251));
    Span4Mux_h I__3870 (
            .O(N__19257),
            .I(N__19248));
    Span4Mux_s3_v I__3869 (
            .O(N__19254),
            .I(N__19243));
    LocalMux I__3868 (
            .O(N__19251),
            .I(N__19243));
    Sp12to4 I__3867 (
            .O(N__19248),
            .I(N__19240));
    Span4Mux_v I__3866 (
            .O(N__19243),
            .I(N__19237));
    Odrv12 I__3865 (
            .O(N__19240),
            .I(\tok.n2732 ));
    Odrv4 I__3864 (
            .O(N__19237),
            .I(\tok.n2732 ));
    CascadeMux I__3863 (
            .O(N__19232),
            .I(\tok.n2732_cascade_ ));
    CascadeMux I__3862 (
            .O(N__19229),
            .I(N__19225));
    CascadeMux I__3861 (
            .O(N__19228),
            .I(N__19222));
    CascadeBuf I__3860 (
            .O(N__19225),
            .I(N__19219));
    CascadeBuf I__3859 (
            .O(N__19222),
            .I(N__19216));
    CascadeMux I__3858 (
            .O(N__19219),
            .I(N__19211));
    CascadeMux I__3857 (
            .O(N__19216),
            .I(N__19208));
    InMux I__3856 (
            .O(N__19215),
            .I(N__19205));
    InMux I__3855 (
            .O(N__19214),
            .I(N__19202));
    InMux I__3854 (
            .O(N__19211),
            .I(N__19199));
    InMux I__3853 (
            .O(N__19208),
            .I(N__19196));
    LocalMux I__3852 (
            .O(N__19205),
            .I(N__19191));
    LocalMux I__3851 (
            .O(N__19202),
            .I(N__19191));
    LocalMux I__3850 (
            .O(N__19199),
            .I(N__19188));
    LocalMux I__3849 (
            .O(N__19196),
            .I(N__19185));
    Span4Mux_h I__3848 (
            .O(N__19191),
            .I(N__19181));
    Span4Mux_h I__3847 (
            .O(N__19188),
            .I(N__19178));
    Span4Mux_h I__3846 (
            .O(N__19185),
            .I(N__19175));
    InMux I__3845 (
            .O(N__19184),
            .I(N__19172));
    Span4Mux_v I__3844 (
            .O(N__19181),
            .I(N__19167));
    Span4Mux_h I__3843 (
            .O(N__19178),
            .I(N__19167));
    Span4Mux_h I__3842 (
            .O(N__19175),
            .I(N__19164));
    LocalMux I__3841 (
            .O(N__19172),
            .I(\tok.n43 ));
    Odrv4 I__3840 (
            .O(N__19167),
            .I(\tok.n43 ));
    Odrv4 I__3839 (
            .O(N__19164),
            .I(\tok.n43 ));
    InMux I__3838 (
            .O(N__19157),
            .I(N__19154));
    LocalMux I__3837 (
            .O(N__19154),
            .I(\tok.n5_adj_655 ));
    SRMux I__3836 (
            .O(N__19151),
            .I(N__19148));
    LocalMux I__3835 (
            .O(N__19148),
            .I(N__19145));
    Span4Mux_h I__3834 (
            .O(N__19145),
            .I(N__19139));
    SRMux I__3833 (
            .O(N__19144),
            .I(N__19136));
    SRMux I__3832 (
            .O(N__19143),
            .I(N__19132));
    SRMux I__3831 (
            .O(N__19142),
            .I(N__19127));
    Span4Mux_h I__3830 (
            .O(N__19139),
            .I(N__19122));
    LocalMux I__3829 (
            .O(N__19136),
            .I(N__19122));
    SRMux I__3828 (
            .O(N__19135),
            .I(N__19119));
    LocalMux I__3827 (
            .O(N__19132),
            .I(N__19115));
    SRMux I__3826 (
            .O(N__19131),
            .I(N__19111));
    SRMux I__3825 (
            .O(N__19130),
            .I(N__19108));
    LocalMux I__3824 (
            .O(N__19127),
            .I(N__19105));
    Span4Mux_v I__3823 (
            .O(N__19122),
            .I(N__19100));
    LocalMux I__3822 (
            .O(N__19119),
            .I(N__19100));
    SRMux I__3821 (
            .O(N__19118),
            .I(N__19097));
    Span4Mux_h I__3820 (
            .O(N__19115),
            .I(N__19093));
    SRMux I__3819 (
            .O(N__19114),
            .I(N__19090));
    LocalMux I__3818 (
            .O(N__19111),
            .I(N__19087));
    LocalMux I__3817 (
            .O(N__19108),
            .I(N__19083));
    Span4Mux_v I__3816 (
            .O(N__19105),
            .I(N__19076));
    Span4Mux_v I__3815 (
            .O(N__19100),
            .I(N__19076));
    LocalMux I__3814 (
            .O(N__19097),
            .I(N__19076));
    SRMux I__3813 (
            .O(N__19096),
            .I(N__19073));
    Span4Mux_v I__3812 (
            .O(N__19093),
            .I(N__19070));
    LocalMux I__3811 (
            .O(N__19090),
            .I(N__19067));
    Span4Mux_v I__3810 (
            .O(N__19087),
            .I(N__19063));
    SRMux I__3809 (
            .O(N__19086),
            .I(N__19060));
    Span4Mux_h I__3808 (
            .O(N__19083),
            .I(N__19053));
    Span4Mux_h I__3807 (
            .O(N__19076),
            .I(N__19053));
    LocalMux I__3806 (
            .O(N__19073),
            .I(N__19053));
    IoSpan4Mux I__3805 (
            .O(N__19070),
            .I(N__19050));
    Span4Mux_v I__3804 (
            .O(N__19067),
            .I(N__19047));
    SRMux I__3803 (
            .O(N__19066),
            .I(N__19044));
    Span4Mux_v I__3802 (
            .O(N__19063),
            .I(N__19039));
    LocalMux I__3801 (
            .O(N__19060),
            .I(N__19039));
    Span4Mux_v I__3800 (
            .O(N__19053),
            .I(N__19036));
    IoSpan4Mux I__3799 (
            .O(N__19050),
            .I(N__19033));
    Span4Mux_h I__3798 (
            .O(N__19047),
            .I(N__19030));
    LocalMux I__3797 (
            .O(N__19044),
            .I(N__19027));
    Span4Mux_v I__3796 (
            .O(N__19039),
            .I(N__19022));
    Span4Mux_h I__3795 (
            .O(N__19036),
            .I(N__19022));
    Span4Mux_s0_v I__3794 (
            .O(N__19033),
            .I(N__19017));
    Span4Mux_v I__3793 (
            .O(N__19030),
            .I(N__19017));
    Span4Mux_v I__3792 (
            .O(N__19027),
            .I(N__19012));
    Span4Mux_s0_v I__3791 (
            .O(N__19022),
            .I(N__19012));
    Odrv4 I__3790 (
            .O(N__19017),
            .I(\tok.reset_N_2 ));
    Odrv4 I__3789 (
            .O(N__19012),
            .I(\tok.reset_N_2 ));
    InMux I__3788 (
            .O(N__19007),
            .I(N__18998));
    InMux I__3787 (
            .O(N__19006),
            .I(N__18998));
    InMux I__3786 (
            .O(N__19005),
            .I(N__18998));
    LocalMux I__3785 (
            .O(N__18998),
            .I(\tok.uart_stall ));
    CascadeMux I__3784 (
            .O(N__18995),
            .I(N__18992));
    InMux I__3783 (
            .O(N__18992),
            .I(N__18980));
    InMux I__3782 (
            .O(N__18991),
            .I(N__18980));
    InMux I__3781 (
            .O(N__18990),
            .I(N__18980));
    InMux I__3780 (
            .O(N__18989),
            .I(N__18980));
    LocalMux I__3779 (
            .O(N__18980),
            .I(N__18977));
    Odrv4 I__3778 (
            .O(N__18977),
            .I(\tok.n2724 ));
    InMux I__3777 (
            .O(N__18974),
            .I(N__18964));
    InMux I__3776 (
            .O(N__18973),
            .I(N__18964));
    InMux I__3775 (
            .O(N__18972),
            .I(N__18955));
    InMux I__3774 (
            .O(N__18971),
            .I(N__18955));
    InMux I__3773 (
            .O(N__18970),
            .I(N__18955));
    InMux I__3772 (
            .O(N__18969),
            .I(N__18955));
    LocalMux I__3771 (
            .O(N__18964),
            .I(N__18949));
    LocalMux I__3770 (
            .O(N__18955),
            .I(N__18949));
    InMux I__3769 (
            .O(N__18954),
            .I(N__18946));
    Span4Mux_s3_v I__3768 (
            .O(N__18949),
            .I(N__18941));
    LocalMux I__3767 (
            .O(N__18946),
            .I(N__18941));
    Span4Mux_v I__3766 (
            .O(N__18941),
            .I(N__18937));
    InMux I__3765 (
            .O(N__18940),
            .I(N__18934));
    Odrv4 I__3764 (
            .O(N__18937),
            .I(\tok.n4431 ));
    LocalMux I__3763 (
            .O(N__18934),
            .I(\tok.n4431 ));
    InMux I__3762 (
            .O(N__18929),
            .I(N__18926));
    LocalMux I__3761 (
            .O(N__18926),
            .I(N__18923));
    Span4Mux_h I__3760 (
            .O(N__18923),
            .I(N__18920));
    Odrv4 I__3759 (
            .O(N__18920),
            .I(\tok.n5_adj_682 ));
    InMux I__3758 (
            .O(N__18917),
            .I(N__18914));
    LocalMux I__3757 (
            .O(N__18914),
            .I(N__18908));
    InMux I__3756 (
            .O(N__18913),
            .I(N__18901));
    InMux I__3755 (
            .O(N__18912),
            .I(N__18901));
    InMux I__3754 (
            .O(N__18911),
            .I(N__18901));
    Odrv4 I__3753 (
            .O(N__18908),
            .I(\tok.tc_plus_1_6 ));
    LocalMux I__3752 (
            .O(N__18901),
            .I(\tok.tc_plus_1_6 ));
    InMux I__3751 (
            .O(N__18896),
            .I(\tok.n3900 ));
    InMux I__3750 (
            .O(N__18893),
            .I(\tok.n3901 ));
    InMux I__3749 (
            .O(N__18890),
            .I(N__18887));
    LocalMux I__3748 (
            .O(N__18887),
            .I(N__18884));
    Span4Mux_v I__3747 (
            .O(N__18884),
            .I(N__18881));
    Span4Mux_h I__3746 (
            .O(N__18881),
            .I(N__18875));
    InMux I__3745 (
            .O(N__18880),
            .I(N__18872));
    InMux I__3744 (
            .O(N__18879),
            .I(N__18867));
    InMux I__3743 (
            .O(N__18878),
            .I(N__18867));
    Odrv4 I__3742 (
            .O(N__18875),
            .I(\tok.tc_plus_1_7 ));
    LocalMux I__3741 (
            .O(N__18872),
            .I(\tok.tc_plus_1_7 ));
    LocalMux I__3740 (
            .O(N__18867),
            .I(\tok.tc_plus_1_7 ));
    InMux I__3739 (
            .O(N__18860),
            .I(N__18857));
    LocalMux I__3738 (
            .O(N__18857),
            .I(N__18853));
    InMux I__3737 (
            .O(N__18856),
            .I(N__18850));
    Odrv4 I__3736 (
            .O(N__18853),
            .I(n92_adj_872));
    LocalMux I__3735 (
            .O(N__18850),
            .I(n92_adj_872));
    CascadeMux I__3734 (
            .O(N__18845),
            .I(N__18842));
    InMux I__3733 (
            .O(N__18842),
            .I(N__18837));
    InMux I__3732 (
            .O(N__18841),
            .I(N__18833));
    InMux I__3731 (
            .O(N__18840),
            .I(N__18830));
    LocalMux I__3730 (
            .O(N__18837),
            .I(N__18827));
    InMux I__3729 (
            .O(N__18836),
            .I(N__18824));
    LocalMux I__3728 (
            .O(N__18833),
            .I(c_stk_w_7_N_18_7));
    LocalMux I__3727 (
            .O(N__18830),
            .I(c_stk_w_7_N_18_7));
    Odrv4 I__3726 (
            .O(N__18827),
            .I(c_stk_w_7_N_18_7));
    LocalMux I__3725 (
            .O(N__18824),
            .I(c_stk_w_7_N_18_7));
    InMux I__3724 (
            .O(N__18815),
            .I(N__18811));
    InMux I__3723 (
            .O(N__18814),
            .I(N__18808));
    LocalMux I__3722 (
            .O(N__18811),
            .I(n92_adj_871));
    LocalMux I__3721 (
            .O(N__18808),
            .I(n92_adj_871));
    InMux I__3720 (
            .O(N__18803),
            .I(N__18798));
    InMux I__3719 (
            .O(N__18802),
            .I(N__18795));
    InMux I__3718 (
            .O(N__18801),
            .I(N__18791));
    LocalMux I__3717 (
            .O(N__18798),
            .I(N__18788));
    LocalMux I__3716 (
            .O(N__18795),
            .I(N__18785));
    InMux I__3715 (
            .O(N__18794),
            .I(N__18782));
    LocalMux I__3714 (
            .O(N__18791),
            .I(c_stk_w_7_N_18_6));
    Odrv4 I__3713 (
            .O(N__18788),
            .I(c_stk_w_7_N_18_6));
    Odrv4 I__3712 (
            .O(N__18785),
            .I(c_stk_w_7_N_18_6));
    LocalMux I__3711 (
            .O(N__18782),
            .I(c_stk_w_7_N_18_6));
    InMux I__3710 (
            .O(N__18773),
            .I(N__18770));
    LocalMux I__3709 (
            .O(N__18770),
            .I(n92));
    InMux I__3708 (
            .O(N__18767),
            .I(N__18761));
    InMux I__3707 (
            .O(N__18766),
            .I(N__18756));
    InMux I__3706 (
            .O(N__18765),
            .I(N__18756));
    InMux I__3705 (
            .O(N__18764),
            .I(N__18753));
    LocalMux I__3704 (
            .O(N__18761),
            .I(c_stk_w_7_N_18_1));
    LocalMux I__3703 (
            .O(N__18756),
            .I(c_stk_w_7_N_18_1));
    LocalMux I__3702 (
            .O(N__18753),
            .I(c_stk_w_7_N_18_1));
    InMux I__3701 (
            .O(N__18746),
            .I(N__18740));
    CascadeMux I__3700 (
            .O(N__18745),
            .I(N__18736));
    CascadeMux I__3699 (
            .O(N__18744),
            .I(N__18733));
    InMux I__3698 (
            .O(N__18743),
            .I(N__18730));
    LocalMux I__3697 (
            .O(N__18740),
            .I(N__18727));
    InMux I__3696 (
            .O(N__18739),
            .I(N__18722));
    InMux I__3695 (
            .O(N__18736),
            .I(N__18722));
    InMux I__3694 (
            .O(N__18733),
            .I(N__18719));
    LocalMux I__3693 (
            .O(N__18730),
            .I(\tok.c_stk_r_7 ));
    Odrv4 I__3692 (
            .O(N__18727),
            .I(\tok.c_stk_r_7 ));
    LocalMux I__3691 (
            .O(N__18722),
            .I(\tok.c_stk_r_7 ));
    LocalMux I__3690 (
            .O(N__18719),
            .I(\tok.c_stk_r_7 ));
    CascadeMux I__3689 (
            .O(N__18710),
            .I(\tok.ram.n4696_cascade_ ));
    InMux I__3688 (
            .O(N__18707),
            .I(N__18704));
    LocalMux I__3687 (
            .O(N__18704),
            .I(\tok.n4602 ));
    CascadeMux I__3686 (
            .O(N__18701),
            .I(\tok.n1_adj_798_cascade_ ));
    InMux I__3685 (
            .O(N__18698),
            .I(N__18695));
    LocalMux I__3684 (
            .O(N__18695),
            .I(\tok.n13_adj_799 ));
    CascadeMux I__3683 (
            .O(N__18692),
            .I(N__18689));
    InMux I__3682 (
            .O(N__18689),
            .I(N__18686));
    LocalMux I__3681 (
            .O(N__18686),
            .I(N__18683));
    Span4Mux_h I__3680 (
            .O(N__18683),
            .I(N__18680));
    Odrv4 I__3679 (
            .O(N__18680),
            .I(\tok.tc_0 ));
    InMux I__3678 (
            .O(N__18677),
            .I(N__18674));
    LocalMux I__3677 (
            .O(N__18674),
            .I(N__18668));
    InMux I__3676 (
            .O(N__18673),
            .I(N__18661));
    InMux I__3675 (
            .O(N__18672),
            .I(N__18661));
    InMux I__3674 (
            .O(N__18671),
            .I(N__18661));
    Span4Mux_v I__3673 (
            .O(N__18668),
            .I(N__18656));
    LocalMux I__3672 (
            .O(N__18661),
            .I(N__18656));
    Odrv4 I__3671 (
            .O(N__18656),
            .I(\tok.tc_plus_1_0 ));
    InMux I__3670 (
            .O(N__18653),
            .I(bfn_9_5_0_));
    InMux I__3669 (
            .O(N__18650),
            .I(N__18647));
    LocalMux I__3668 (
            .O(N__18647),
            .I(N__18644));
    Span12Mux_s9_v I__3667 (
            .O(N__18644),
            .I(N__18638));
    InMux I__3666 (
            .O(N__18643),
            .I(N__18631));
    InMux I__3665 (
            .O(N__18642),
            .I(N__18631));
    InMux I__3664 (
            .O(N__18641),
            .I(N__18631));
    Odrv12 I__3663 (
            .O(N__18638),
            .I(\tok.tc_plus_1_1 ));
    LocalMux I__3662 (
            .O(N__18631),
            .I(\tok.tc_plus_1_1 ));
    InMux I__3661 (
            .O(N__18626),
            .I(\tok.n3895 ));
    InMux I__3660 (
            .O(N__18623),
            .I(\tok.n3896 ));
    InMux I__3659 (
            .O(N__18620),
            .I(\tok.n3897 ));
    InMux I__3658 (
            .O(N__18617),
            .I(\tok.n3898 ));
    InMux I__3657 (
            .O(N__18614),
            .I(\tok.n3899 ));
    CascadeMux I__3656 (
            .O(N__18611),
            .I(\tok.n13_adj_713_cascade_ ));
    CascadeMux I__3655 (
            .O(N__18608),
            .I(\tok.C_stk.n4894_cascade_ ));
    CascadeMux I__3654 (
            .O(N__18605),
            .I(N__18599));
    InMux I__3653 (
            .O(N__18604),
            .I(N__18595));
    InMux I__3652 (
            .O(N__18603),
            .I(N__18592));
    InMux I__3651 (
            .O(N__18602),
            .I(N__18587));
    InMux I__3650 (
            .O(N__18599),
            .I(N__18587));
    InMux I__3649 (
            .O(N__18598),
            .I(N__18584));
    LocalMux I__3648 (
            .O(N__18595),
            .I(\tok.c_stk_r_0 ));
    LocalMux I__3647 (
            .O(N__18592),
            .I(\tok.c_stk_r_0 ));
    LocalMux I__3646 (
            .O(N__18587),
            .I(\tok.c_stk_r_0 ));
    LocalMux I__3645 (
            .O(N__18584),
            .I(\tok.c_stk_r_0 ));
    CascadeMux I__3644 (
            .O(N__18575),
            .I(\tok.ram.n4717_cascade_ ));
    InMux I__3643 (
            .O(N__18572),
            .I(N__18569));
    LocalMux I__3642 (
            .O(N__18569),
            .I(\tok.n1_adj_712 ));
    InMux I__3641 (
            .O(N__18566),
            .I(N__18563));
    LocalMux I__3640 (
            .O(N__18563),
            .I(N__18559));
    InMux I__3639 (
            .O(N__18562),
            .I(N__18556));
    Odrv4 I__3638 (
            .O(N__18559),
            .I(\tok.C_stk.tail_7 ));
    LocalMux I__3637 (
            .O(N__18556),
            .I(\tok.C_stk.tail_7 ));
    CascadeMux I__3636 (
            .O(N__18551),
            .I(\tok.C_stk.n4912_cascade_ ));
    CascadeMux I__3635 (
            .O(N__18548),
            .I(N__18545));
    InMux I__3634 (
            .O(N__18545),
            .I(N__18542));
    LocalMux I__3633 (
            .O(N__18542),
            .I(N__18539));
    Odrv4 I__3632 (
            .O(N__18539),
            .I(\tok.tc_6 ));
    InMux I__3631 (
            .O(N__18536),
            .I(N__18532));
    InMux I__3630 (
            .O(N__18535),
            .I(N__18529));
    LocalMux I__3629 (
            .O(N__18532),
            .I(\tok.tail_26 ));
    LocalMux I__3628 (
            .O(N__18529),
            .I(\tok.tail_26 ));
    InMux I__3627 (
            .O(N__18524),
            .I(N__18520));
    InMux I__3626 (
            .O(N__18523),
            .I(N__18517));
    LocalMux I__3625 (
            .O(N__18520),
            .I(\tok.tail_12 ));
    LocalMux I__3624 (
            .O(N__18517),
            .I(\tok.tail_12 ));
    InMux I__3623 (
            .O(N__18512),
            .I(N__18508));
    InMux I__3622 (
            .O(N__18511),
            .I(N__18505));
    LocalMux I__3621 (
            .O(N__18508),
            .I(\tok.C_stk.tail_36 ));
    LocalMux I__3620 (
            .O(N__18505),
            .I(\tok.C_stk.tail_36 ));
    InMux I__3619 (
            .O(N__18500),
            .I(N__18497));
    LocalMux I__3618 (
            .O(N__18497),
            .I(N__18494));
    Span4Mux_s2_v I__3617 (
            .O(N__18494),
            .I(N__18490));
    InMux I__3616 (
            .O(N__18493),
            .I(N__18487));
    Odrv4 I__3615 (
            .O(N__18490),
            .I(\tok.tail_56 ));
    LocalMux I__3614 (
            .O(N__18487),
            .I(\tok.tail_56 ));
    InMux I__3613 (
            .O(N__18482),
            .I(N__18478));
    InMux I__3612 (
            .O(N__18481),
            .I(N__18475));
    LocalMux I__3611 (
            .O(N__18478),
            .I(\tok.tail_40 ));
    LocalMux I__3610 (
            .O(N__18475),
            .I(\tok.tail_40 ));
    CascadeMux I__3609 (
            .O(N__18470),
            .I(N__18467));
    InMux I__3608 (
            .O(N__18467),
            .I(N__18464));
    LocalMux I__3607 (
            .O(N__18464),
            .I(N__18461));
    Span4Mux_v I__3606 (
            .O(N__18461),
            .I(N__18457));
    InMux I__3605 (
            .O(N__18460),
            .I(N__18454));
    Odrv4 I__3604 (
            .O(N__18457),
            .I(\tok.tail_48 ));
    LocalMux I__3603 (
            .O(N__18454),
            .I(\tok.tail_48 ));
    InMux I__3602 (
            .O(N__18449),
            .I(N__18446));
    LocalMux I__3601 (
            .O(N__18446),
            .I(N__18443));
    Odrv4 I__3600 (
            .O(N__18443),
            .I(\tok.n83_adj_704 ));
    CascadeMux I__3599 (
            .O(N__18440),
            .I(\tok.n4694_cascade_ ));
    CascadeMux I__3598 (
            .O(N__18437),
            .I(N__18433));
    CascadeMux I__3597 (
            .O(N__18436),
            .I(N__18430));
    CascadeBuf I__3596 (
            .O(N__18433),
            .I(N__18427));
    CascadeBuf I__3595 (
            .O(N__18430),
            .I(N__18424));
    CascadeMux I__3594 (
            .O(N__18427),
            .I(N__18421));
    CascadeMux I__3593 (
            .O(N__18424),
            .I(N__18418));
    InMux I__3592 (
            .O(N__18421),
            .I(N__18415));
    InMux I__3591 (
            .O(N__18418),
            .I(N__18412));
    LocalMux I__3590 (
            .O(N__18415),
            .I(N__18409));
    LocalMux I__3589 (
            .O(N__18412),
            .I(N__18403));
    Span4Mux_h I__3588 (
            .O(N__18409),
            .I(N__18400));
    InMux I__3587 (
            .O(N__18408),
            .I(N__18397));
    InMux I__3586 (
            .O(N__18407),
            .I(N__18394));
    InMux I__3585 (
            .O(N__18406),
            .I(N__18391));
    Span4Mux_v I__3584 (
            .O(N__18403),
            .I(N__18388));
    Span4Mux_h I__3583 (
            .O(N__18400),
            .I(N__18385));
    LocalMux I__3582 (
            .O(N__18397),
            .I(\tok.n50 ));
    LocalMux I__3581 (
            .O(N__18394),
            .I(\tok.n50 ));
    LocalMux I__3580 (
            .O(N__18391),
            .I(\tok.n50 ));
    Odrv4 I__3579 (
            .O(N__18388),
            .I(\tok.n50 ));
    Odrv4 I__3578 (
            .O(N__18385),
            .I(\tok.n50 ));
    InMux I__3577 (
            .O(N__18374),
            .I(N__18371));
    LocalMux I__3576 (
            .O(N__18371),
            .I(\tok.n33_adj_841 ));
    InMux I__3575 (
            .O(N__18368),
            .I(\tok.n3888 ));
    CascadeMux I__3574 (
            .O(N__18365),
            .I(N__18361));
    CascadeMux I__3573 (
            .O(N__18364),
            .I(N__18358));
    CascadeBuf I__3572 (
            .O(N__18361),
            .I(N__18355));
    CascadeBuf I__3571 (
            .O(N__18358),
            .I(N__18352));
    CascadeMux I__3570 (
            .O(N__18355),
            .I(N__18349));
    CascadeMux I__3569 (
            .O(N__18352),
            .I(N__18346));
    InMux I__3568 (
            .O(N__18349),
            .I(N__18343));
    InMux I__3567 (
            .O(N__18346),
            .I(N__18340));
    LocalMux I__3566 (
            .O(N__18343),
            .I(N__18335));
    LocalMux I__3565 (
            .O(N__18340),
            .I(N__18335));
    Span4Mux_v I__3564 (
            .O(N__18335),
            .I(N__18329));
    InMux I__3563 (
            .O(N__18334),
            .I(N__18326));
    InMux I__3562 (
            .O(N__18333),
            .I(N__18323));
    InMux I__3561 (
            .O(N__18332),
            .I(N__18320));
    Span4Mux_h I__3560 (
            .O(N__18329),
            .I(N__18317));
    LocalMux I__3559 (
            .O(N__18326),
            .I(\tok.n49 ));
    LocalMux I__3558 (
            .O(N__18323),
            .I(\tok.n49 ));
    LocalMux I__3557 (
            .O(N__18320),
            .I(\tok.n49 ));
    Odrv4 I__3556 (
            .O(N__18317),
            .I(\tok.n49 ));
    CascadeMux I__3555 (
            .O(N__18308),
            .I(N__18305));
    InMux I__3554 (
            .O(N__18305),
            .I(N__18302));
    LocalMux I__3553 (
            .O(N__18302),
            .I(\tok.n33_adj_665 ));
    InMux I__3552 (
            .O(N__18299),
            .I(\tok.n3889 ));
    CascadeMux I__3551 (
            .O(N__18296),
            .I(N__18292));
    CascadeMux I__3550 (
            .O(N__18295),
            .I(N__18289));
    CascadeBuf I__3549 (
            .O(N__18292),
            .I(N__18286));
    CascadeBuf I__3548 (
            .O(N__18289),
            .I(N__18283));
    CascadeMux I__3547 (
            .O(N__18286),
            .I(N__18280));
    CascadeMux I__3546 (
            .O(N__18283),
            .I(N__18277));
    InMux I__3545 (
            .O(N__18280),
            .I(N__18274));
    InMux I__3544 (
            .O(N__18277),
            .I(N__18270));
    LocalMux I__3543 (
            .O(N__18274),
            .I(N__18267));
    CascadeMux I__3542 (
            .O(N__18273),
            .I(N__18264));
    LocalMux I__3541 (
            .O(N__18270),
            .I(N__18257));
    Span4Mux_v I__3540 (
            .O(N__18267),
            .I(N__18257));
    InMux I__3539 (
            .O(N__18264),
            .I(N__18254));
    InMux I__3538 (
            .O(N__18263),
            .I(N__18251));
    InMux I__3537 (
            .O(N__18262),
            .I(N__18248));
    Span4Mux_h I__3536 (
            .O(N__18257),
            .I(N__18245));
    LocalMux I__3535 (
            .O(N__18254),
            .I(\tok.n47 ));
    LocalMux I__3534 (
            .O(N__18251),
            .I(\tok.n47 ));
    LocalMux I__3533 (
            .O(N__18248),
            .I(\tok.n47 ));
    Odrv4 I__3532 (
            .O(N__18245),
            .I(\tok.n47 ));
    InMux I__3531 (
            .O(N__18236),
            .I(N__18233));
    LocalMux I__3530 (
            .O(N__18233),
            .I(N__18230));
    Span4Mux_v I__3529 (
            .O(N__18230),
            .I(N__18227));
    Odrv4 I__3528 (
            .O(N__18227),
            .I(\tok.n33_adj_755 ));
    InMux I__3527 (
            .O(N__18224),
            .I(\tok.n3890 ));
    CascadeMux I__3526 (
            .O(N__18221),
            .I(N__18217));
    CascadeMux I__3525 (
            .O(N__18220),
            .I(N__18214));
    CascadeBuf I__3524 (
            .O(N__18217),
            .I(N__18209));
    CascadeBuf I__3523 (
            .O(N__18214),
            .I(N__18206));
    InMux I__3522 (
            .O(N__18213),
            .I(N__18203));
    InMux I__3521 (
            .O(N__18212),
            .I(N__18200));
    CascadeMux I__3520 (
            .O(N__18209),
            .I(N__18197));
    CascadeMux I__3519 (
            .O(N__18206),
            .I(N__18194));
    LocalMux I__3518 (
            .O(N__18203),
            .I(N__18189));
    LocalMux I__3517 (
            .O(N__18200),
            .I(N__18189));
    InMux I__3516 (
            .O(N__18197),
            .I(N__18186));
    InMux I__3515 (
            .O(N__18194),
            .I(N__18183));
    Span4Mux_s2_v I__3514 (
            .O(N__18189),
            .I(N__18180));
    LocalMux I__3513 (
            .O(N__18186),
            .I(N__18175));
    LocalMux I__3512 (
            .O(N__18183),
            .I(N__18175));
    Span4Mux_v I__3511 (
            .O(N__18180),
            .I(N__18171));
    Sp12to4 I__3510 (
            .O(N__18175),
            .I(N__18168));
    InMux I__3509 (
            .O(N__18174),
            .I(N__18165));
    Sp12to4 I__3508 (
            .O(N__18171),
            .I(N__18160));
    Span12Mux_s6_v I__3507 (
            .O(N__18168),
            .I(N__18160));
    LocalMux I__3506 (
            .O(N__18165),
            .I(\tok.n45 ));
    Odrv12 I__3505 (
            .O(N__18160),
            .I(\tok.n45 ));
    CascadeMux I__3504 (
            .O(N__18155),
            .I(N__18152));
    InMux I__3503 (
            .O(N__18152),
            .I(N__18149));
    LocalMux I__3502 (
            .O(N__18149),
            .I(N__18146));
    Span4Mux_v I__3501 (
            .O(N__18146),
            .I(N__18143));
    Odrv4 I__3500 (
            .O(N__18143),
            .I(\tok.n33_adj_852 ));
    InMux I__3499 (
            .O(N__18140),
            .I(\tok.n3891 ));
    CascadeMux I__3498 (
            .O(N__18137),
            .I(N__18133));
    CascadeMux I__3497 (
            .O(N__18136),
            .I(N__18130));
    CascadeBuf I__3496 (
            .O(N__18133),
            .I(N__18127));
    CascadeBuf I__3495 (
            .O(N__18130),
            .I(N__18124));
    CascadeMux I__3494 (
            .O(N__18127),
            .I(N__18121));
    CascadeMux I__3493 (
            .O(N__18124),
            .I(N__18118));
    InMux I__3492 (
            .O(N__18121),
            .I(N__18115));
    InMux I__3491 (
            .O(N__18118),
            .I(N__18109));
    LocalMux I__3490 (
            .O(N__18115),
            .I(N__18106));
    CascadeMux I__3489 (
            .O(N__18114),
            .I(N__18103));
    InMux I__3488 (
            .O(N__18113),
            .I(N__18100));
    InMux I__3487 (
            .O(N__18112),
            .I(N__18097));
    LocalMux I__3486 (
            .O(N__18109),
            .I(N__18092));
    Span4Mux_h I__3485 (
            .O(N__18106),
            .I(N__18092));
    InMux I__3484 (
            .O(N__18103),
            .I(N__18089));
    LocalMux I__3483 (
            .O(N__18100),
            .I(N__18084));
    LocalMux I__3482 (
            .O(N__18097),
            .I(N__18084));
    Span4Mux_v I__3481 (
            .O(N__18092),
            .I(N__18081));
    LocalMux I__3480 (
            .O(N__18089),
            .I(\tok.n44 ));
    Odrv12 I__3479 (
            .O(N__18084),
            .I(\tok.n44 ));
    Odrv4 I__3478 (
            .O(N__18081),
            .I(\tok.n44 ));
    InMux I__3477 (
            .O(N__18074),
            .I(\tok.n3892 ));
    InMux I__3476 (
            .O(N__18071),
            .I(\tok.n3893 ));
    CascadeMux I__3475 (
            .O(N__18068),
            .I(N__18064));
    CascadeMux I__3474 (
            .O(N__18067),
            .I(N__18061));
    CascadeBuf I__3473 (
            .O(N__18064),
            .I(N__18058));
    CascadeBuf I__3472 (
            .O(N__18061),
            .I(N__18055));
    CascadeMux I__3471 (
            .O(N__18058),
            .I(N__18052));
    CascadeMux I__3470 (
            .O(N__18055),
            .I(N__18049));
    InMux I__3469 (
            .O(N__18052),
            .I(N__18046));
    InMux I__3468 (
            .O(N__18049),
            .I(N__18041));
    LocalMux I__3467 (
            .O(N__18046),
            .I(N__18038));
    InMux I__3466 (
            .O(N__18045),
            .I(N__18034));
    InMux I__3465 (
            .O(N__18044),
            .I(N__18031));
    LocalMux I__3464 (
            .O(N__18041),
            .I(N__18028));
    Span4Mux_h I__3463 (
            .O(N__18038),
            .I(N__18025));
    InMux I__3462 (
            .O(N__18037),
            .I(N__18022));
    LocalMux I__3461 (
            .O(N__18034),
            .I(N__18017));
    LocalMux I__3460 (
            .O(N__18031),
            .I(N__18017));
    Span4Mux_v I__3459 (
            .O(N__18028),
            .I(N__18014));
    Span4Mux_v I__3458 (
            .O(N__18025),
            .I(N__18011));
    LocalMux I__3457 (
            .O(N__18022),
            .I(\tok.n39 ));
    Odrv4 I__3456 (
            .O(N__18017),
            .I(\tok.n39 ));
    Odrv4 I__3455 (
            .O(N__18014),
            .I(\tok.n39 ));
    Odrv4 I__3454 (
            .O(N__18011),
            .I(\tok.n39 ));
    InMux I__3453 (
            .O(N__18002),
            .I(\tok.n3894 ));
    InMux I__3452 (
            .O(N__17999),
            .I(N__17996));
    LocalMux I__3451 (
            .O(N__17996),
            .I(N__17993));
    Odrv4 I__3450 (
            .O(N__17993),
            .I(\tok.n33_adj_643 ));
    InMux I__3449 (
            .O(N__17990),
            .I(N__17986));
    InMux I__3448 (
            .O(N__17989),
            .I(N__17983));
    LocalMux I__3447 (
            .O(N__17986),
            .I(\tok.C_stk.tail_20 ));
    LocalMux I__3446 (
            .O(N__17983),
            .I(\tok.C_stk.tail_20 ));
    InMux I__3445 (
            .O(N__17978),
            .I(N__17975));
    LocalMux I__3444 (
            .O(N__17975),
            .I(N__17972));
    Span4Mux_v I__3443 (
            .O(N__17972),
            .I(N__17969));
    Span4Mux_s2_v I__3442 (
            .O(N__17969),
            .I(N__17966));
    Odrv4 I__3441 (
            .O(N__17966),
            .I(\tok.n9_adj_689 ));
    CascadeMux I__3440 (
            .O(N__17963),
            .I(\tok.n181_cascade_ ));
    CascadeMux I__3439 (
            .O(N__17960),
            .I(\tok.n12_cascade_ ));
    InMux I__3438 (
            .O(N__17957),
            .I(N__17954));
    LocalMux I__3437 (
            .O(N__17954),
            .I(N__17951));
    Odrv12 I__3436 (
            .O(N__17951),
            .I(\tok.n6_adj_653 ));
    CascadeMux I__3435 (
            .O(N__17948),
            .I(\tok.n20_cascade_ ));
    InMux I__3434 (
            .O(N__17945),
            .I(N__17942));
    LocalMux I__3433 (
            .O(N__17942),
            .I(N__17939));
    Odrv4 I__3432 (
            .O(N__17939),
            .I(\tok.n16 ));
    InMux I__3431 (
            .O(N__17936),
            .I(N__17933));
    LocalMux I__3430 (
            .O(N__17933),
            .I(N__17930));
    Span4Mux_h I__3429 (
            .O(N__17930),
            .I(N__17927));
    Odrv4 I__3428 (
            .O(N__17927),
            .I(\tok.n4684 ));
    InMux I__3427 (
            .O(N__17924),
            .I(N__17916));
    InMux I__3426 (
            .O(N__17923),
            .I(N__17916));
    InMux I__3425 (
            .O(N__17922),
            .I(N__17913));
    InMux I__3424 (
            .O(N__17921),
            .I(N__17910));
    LocalMux I__3423 (
            .O(N__17916),
            .I(N__17905));
    LocalMux I__3422 (
            .O(N__17913),
            .I(N__17899));
    LocalMux I__3421 (
            .O(N__17910),
            .I(N__17899));
    InMux I__3420 (
            .O(N__17909),
            .I(N__17894));
    InMux I__3419 (
            .O(N__17908),
            .I(N__17894));
    Span4Mux_h I__3418 (
            .O(N__17905),
            .I(N__17885));
    InMux I__3417 (
            .O(N__17904),
            .I(N__17882));
    Span4Mux_h I__3416 (
            .O(N__17899),
            .I(N__17875));
    LocalMux I__3415 (
            .O(N__17894),
            .I(N__17875));
    InMux I__3414 (
            .O(N__17893),
            .I(N__17870));
    InMux I__3413 (
            .O(N__17892),
            .I(N__17870));
    InMux I__3412 (
            .O(N__17891),
            .I(N__17865));
    InMux I__3411 (
            .O(N__17890),
            .I(N__17865));
    InMux I__3410 (
            .O(N__17889),
            .I(N__17862));
    InMux I__3409 (
            .O(N__17888),
            .I(N__17859));
    Span4Mux_h I__3408 (
            .O(N__17885),
            .I(N__17854));
    LocalMux I__3407 (
            .O(N__17882),
            .I(N__17854));
    InMux I__3406 (
            .O(N__17881),
            .I(N__17849));
    InMux I__3405 (
            .O(N__17880),
            .I(N__17849));
    Odrv4 I__3404 (
            .O(N__17875),
            .I(\tok.n892 ));
    LocalMux I__3403 (
            .O(N__17870),
            .I(\tok.n892 ));
    LocalMux I__3402 (
            .O(N__17865),
            .I(\tok.n892 ));
    LocalMux I__3401 (
            .O(N__17862),
            .I(\tok.n892 ));
    LocalMux I__3400 (
            .O(N__17859),
            .I(\tok.n892 ));
    Odrv4 I__3399 (
            .O(N__17854),
            .I(\tok.n892 ));
    LocalMux I__3398 (
            .O(N__17849),
            .I(\tok.n892 ));
    CascadeMux I__3397 (
            .O(N__17834),
            .I(\tok.n177_cascade_ ));
    CascadeMux I__3396 (
            .O(N__17831),
            .I(\tok.n12_adj_696_cascade_ ));
    InMux I__3395 (
            .O(N__17828),
            .I(N__17825));
    LocalMux I__3394 (
            .O(N__17825),
            .I(N__17822));
    Odrv12 I__3393 (
            .O(N__17822),
            .I(\tok.n20_adj_700 ));
    CascadeMux I__3392 (
            .O(N__17819),
            .I(N__17815));
    CascadeMux I__3391 (
            .O(N__17818),
            .I(N__17812));
    CascadeBuf I__3390 (
            .O(N__17815),
            .I(N__17809));
    CascadeBuf I__3389 (
            .O(N__17812),
            .I(N__17806));
    CascadeMux I__3388 (
            .O(N__17809),
            .I(N__17803));
    CascadeMux I__3387 (
            .O(N__17806),
            .I(N__17800));
    InMux I__3386 (
            .O(N__17803),
            .I(N__17797));
    InMux I__3385 (
            .O(N__17800),
            .I(N__17793));
    LocalMux I__3384 (
            .O(N__17797),
            .I(N__17790));
    CascadeMux I__3383 (
            .O(N__17796),
            .I(N__17787));
    LocalMux I__3382 (
            .O(N__17793),
            .I(N__17780));
    Span4Mux_h I__3381 (
            .O(N__17790),
            .I(N__17780));
    InMux I__3380 (
            .O(N__17787),
            .I(N__17777));
    InMux I__3379 (
            .O(N__17786),
            .I(N__17774));
    InMux I__3378 (
            .O(N__17785),
            .I(N__17771));
    Span4Mux_v I__3377 (
            .O(N__17780),
            .I(N__17768));
    LocalMux I__3376 (
            .O(N__17777),
            .I(\tok.n52 ));
    LocalMux I__3375 (
            .O(N__17774),
            .I(\tok.n52 ));
    LocalMux I__3374 (
            .O(N__17771),
            .I(\tok.n52 ));
    Odrv4 I__3373 (
            .O(N__17768),
            .I(\tok.n52 ));
    InMux I__3372 (
            .O(N__17759),
            .I(N__17756));
    LocalMux I__3371 (
            .O(N__17756),
            .I(\tok.n33_adj_663 ));
    InMux I__3370 (
            .O(N__17753),
            .I(bfn_8_13_0_));
    InMux I__3369 (
            .O(N__17750),
            .I(N__17745));
    InMux I__3368 (
            .O(N__17749),
            .I(N__17742));
    InMux I__3367 (
            .O(N__17748),
            .I(N__17739));
    LocalMux I__3366 (
            .O(N__17745),
            .I(N__17732));
    LocalMux I__3365 (
            .O(N__17742),
            .I(N__17729));
    LocalMux I__3364 (
            .O(N__17739),
            .I(N__17726));
    InMux I__3363 (
            .O(N__17738),
            .I(N__17723));
    InMux I__3362 (
            .O(N__17737),
            .I(N__17716));
    InMux I__3361 (
            .O(N__17736),
            .I(N__17716));
    InMux I__3360 (
            .O(N__17735),
            .I(N__17716));
    Span4Mux_h I__3359 (
            .O(N__17732),
            .I(N__17710));
    Span4Mux_v I__3358 (
            .O(N__17729),
            .I(N__17710));
    Span4Mux_h I__3357 (
            .O(N__17726),
            .I(N__17703));
    LocalMux I__3356 (
            .O(N__17723),
            .I(N__17703));
    LocalMux I__3355 (
            .O(N__17716),
            .I(N__17703));
    InMux I__3354 (
            .O(N__17715),
            .I(N__17700));
    Odrv4 I__3353 (
            .O(N__17710),
            .I(\tok.A__15__N_129 ));
    Odrv4 I__3352 (
            .O(N__17703),
            .I(\tok.A__15__N_129 ));
    LocalMux I__3351 (
            .O(N__17700),
            .I(\tok.A__15__N_129 ));
    InMux I__3350 (
            .O(N__17693),
            .I(N__17687));
    InMux I__3349 (
            .O(N__17692),
            .I(N__17687));
    LocalMux I__3348 (
            .O(N__17687),
            .I(\tok.A_15_N_113_3 ));
    InMux I__3347 (
            .O(N__17684),
            .I(N__17681));
    LocalMux I__3346 (
            .O(N__17681),
            .I(\tok.A_3 ));
    CascadeMux I__3345 (
            .O(N__17678),
            .I(\tok.n4528_cascade_ ));
    CascadeMux I__3344 (
            .O(N__17675),
            .I(\tok.n892_cascade_ ));
    InMux I__3343 (
            .O(N__17672),
            .I(N__17669));
    LocalMux I__3342 (
            .O(N__17669),
            .I(N__17666));
    Span4Mux_h I__3341 (
            .O(N__17666),
            .I(N__17663));
    Odrv4 I__3340 (
            .O(N__17663),
            .I(\tok.n10_adj_818 ));
    InMux I__3339 (
            .O(N__17660),
            .I(N__17657));
    LocalMux I__3338 (
            .O(N__17657),
            .I(N__17654));
    Odrv4 I__3337 (
            .O(N__17654),
            .I(\tok.n13_adj_842 ));
    InMux I__3336 (
            .O(N__17651),
            .I(N__17648));
    LocalMux I__3335 (
            .O(N__17648),
            .I(\tok.n8_adj_666 ));
    InMux I__3334 (
            .O(N__17645),
            .I(N__17639));
    InMux I__3333 (
            .O(N__17644),
            .I(N__17636));
    InMux I__3332 (
            .O(N__17643),
            .I(N__17631));
    InMux I__3331 (
            .O(N__17642),
            .I(N__17631));
    LocalMux I__3330 (
            .O(N__17639),
            .I(N__17628));
    LocalMux I__3329 (
            .O(N__17636),
            .I(N__17625));
    LocalMux I__3328 (
            .O(N__17631),
            .I(N__17622));
    Span4Mux_s3_v I__3327 (
            .O(N__17628),
            .I(N__17617));
    Span4Mux_v I__3326 (
            .O(N__17625),
            .I(N__17617));
    Span4Mux_h I__3325 (
            .O(N__17622),
            .I(N__17614));
    Odrv4 I__3324 (
            .O(N__17617),
            .I(\tok.n8_adj_777 ));
    Odrv4 I__3323 (
            .O(N__17614),
            .I(\tok.n8_adj_777 ));
    CascadeMux I__3322 (
            .O(N__17609),
            .I(\tok.n4502_cascade_ ));
    InMux I__3321 (
            .O(N__17606),
            .I(N__17603));
    LocalMux I__3320 (
            .O(N__17603),
            .I(\tok.n12_adj_830 ));
    InMux I__3319 (
            .O(N__17600),
            .I(N__17597));
    LocalMux I__3318 (
            .O(N__17597),
            .I(N__17594));
    Span4Mux_s3_v I__3317 (
            .O(N__17594),
            .I(N__17591));
    Span4Mux_v I__3316 (
            .O(N__17591),
            .I(N__17588));
    Odrv4 I__3315 (
            .O(N__17588),
            .I(\tok.n4607 ));
    CascadeMux I__3314 (
            .O(N__17585),
            .I(\tok.n2616_cascade_ ));
    InMux I__3313 (
            .O(N__17582),
            .I(N__17579));
    LocalMux I__3312 (
            .O(N__17579),
            .I(N__17576));
    Odrv4 I__3311 (
            .O(N__17576),
            .I(\tok.n10_adj_849 ));
    InMux I__3310 (
            .O(N__17573),
            .I(N__17570));
    LocalMux I__3309 (
            .O(N__17570),
            .I(N__17567));
    Odrv4 I__3308 (
            .O(N__17567),
            .I(\tok.n12_adj_851 ));
    InMux I__3307 (
            .O(N__17564),
            .I(N__17560));
    CascadeMux I__3306 (
            .O(N__17563),
            .I(N__17557));
    LocalMux I__3305 (
            .O(N__17560),
            .I(N__17554));
    InMux I__3304 (
            .O(N__17557),
            .I(N__17551));
    Span4Mux_h I__3303 (
            .O(N__17554),
            .I(N__17548));
    LocalMux I__3302 (
            .O(N__17551),
            .I(N__17545));
    Span4Mux_h I__3301 (
            .O(N__17548),
            .I(N__17540));
    Span4Mux_h I__3300 (
            .O(N__17545),
            .I(N__17540));
    Span4Mux_v I__3299 (
            .O(N__17540),
            .I(N__17537));
    Odrv4 I__3298 (
            .O(N__17537),
            .I(\tok.table_rd_1 ));
    InMux I__3297 (
            .O(N__17534),
            .I(N__17531));
    LocalMux I__3296 (
            .O(N__17531),
            .I(\tok.n8_adj_850 ));
    InMux I__3295 (
            .O(N__17528),
            .I(N__17525));
    LocalMux I__3294 (
            .O(N__17525),
            .I(\tok.A_4 ));
    InMux I__3293 (
            .O(N__17522),
            .I(N__17513));
    InMux I__3292 (
            .O(N__17521),
            .I(N__17510));
    CascadeMux I__3291 (
            .O(N__17520),
            .I(N__17505));
    CascadeMux I__3290 (
            .O(N__17519),
            .I(N__17502));
    InMux I__3289 (
            .O(N__17518),
            .I(N__17490));
    InMux I__3288 (
            .O(N__17517),
            .I(N__17490));
    InMux I__3287 (
            .O(N__17516),
            .I(N__17490));
    LocalMux I__3286 (
            .O(N__17513),
            .I(N__17483));
    LocalMux I__3285 (
            .O(N__17510),
            .I(N__17483));
    InMux I__3284 (
            .O(N__17509),
            .I(N__17480));
    InMux I__3283 (
            .O(N__17508),
            .I(N__17475));
    InMux I__3282 (
            .O(N__17505),
            .I(N__17475));
    InMux I__3281 (
            .O(N__17502),
            .I(N__17472));
    InMux I__3280 (
            .O(N__17501),
            .I(N__17463));
    InMux I__3279 (
            .O(N__17500),
            .I(N__17463));
    InMux I__3278 (
            .O(N__17499),
            .I(N__17463));
    InMux I__3277 (
            .O(N__17498),
            .I(N__17463));
    InMux I__3276 (
            .O(N__17497),
            .I(N__17460));
    LocalMux I__3275 (
            .O(N__17490),
            .I(N__17457));
    InMux I__3274 (
            .O(N__17489),
            .I(N__17454));
    InMux I__3273 (
            .O(N__17488),
            .I(N__17451));
    Span4Mux_v I__3272 (
            .O(N__17483),
            .I(N__17442));
    LocalMux I__3271 (
            .O(N__17480),
            .I(N__17442));
    LocalMux I__3270 (
            .O(N__17475),
            .I(N__17442));
    LocalMux I__3269 (
            .O(N__17472),
            .I(N__17442));
    LocalMux I__3268 (
            .O(N__17463),
            .I(N__17439));
    LocalMux I__3267 (
            .O(N__17460),
            .I(N__17436));
    Span4Mux_v I__3266 (
            .O(N__17457),
            .I(N__17431));
    LocalMux I__3265 (
            .O(N__17454),
            .I(N__17431));
    LocalMux I__3264 (
            .O(N__17451),
            .I(N__17428));
    Span4Mux_v I__3263 (
            .O(N__17442),
            .I(N__17425));
    Span4Mux_v I__3262 (
            .O(N__17439),
            .I(N__17416));
    Span4Mux_v I__3261 (
            .O(N__17436),
            .I(N__17416));
    Span4Mux_h I__3260 (
            .O(N__17431),
            .I(N__17416));
    Span4Mux_h I__3259 (
            .O(N__17428),
            .I(N__17416));
    Odrv4 I__3258 (
            .O(N__17425),
            .I(\tok.n4051 ));
    Odrv4 I__3257 (
            .O(N__17416),
            .I(\tok.n4051 ));
    InMux I__3256 (
            .O(N__17411),
            .I(N__17408));
    LocalMux I__3255 (
            .O(N__17408),
            .I(\tok.A_15_N_113_4 ));
    CascadeMux I__3254 (
            .O(N__17405),
            .I(\tok.A_15_N_113_4_cascade_ ));
    InMux I__3253 (
            .O(N__17402),
            .I(N__17399));
    LocalMux I__3252 (
            .O(N__17399),
            .I(\tok.A_15_N_113_0 ));
    InMux I__3251 (
            .O(N__17396),
            .I(N__17393));
    LocalMux I__3250 (
            .O(N__17393),
            .I(\tok.A_15_N_113_6 ));
    InMux I__3249 (
            .O(N__17390),
            .I(N__17386));
    CascadeMux I__3248 (
            .O(N__17389),
            .I(N__17382));
    LocalMux I__3247 (
            .O(N__17386),
            .I(N__17375));
    CascadeMux I__3246 (
            .O(N__17385),
            .I(N__17371));
    InMux I__3245 (
            .O(N__17382),
            .I(N__17361));
    InMux I__3244 (
            .O(N__17381),
            .I(N__17361));
    InMux I__3243 (
            .O(N__17380),
            .I(N__17361));
    InMux I__3242 (
            .O(N__17379),
            .I(N__17356));
    InMux I__3241 (
            .O(N__17378),
            .I(N__17356));
    Span4Mux_h I__3240 (
            .O(N__17375),
            .I(N__17353));
    CascadeMux I__3239 (
            .O(N__17374),
            .I(N__17350));
    InMux I__3238 (
            .O(N__17371),
            .I(N__17335));
    InMux I__3237 (
            .O(N__17370),
            .I(N__17335));
    InMux I__3236 (
            .O(N__17369),
            .I(N__17335));
    InMux I__3235 (
            .O(N__17368),
            .I(N__17335));
    LocalMux I__3234 (
            .O(N__17361),
            .I(N__17332));
    LocalMux I__3233 (
            .O(N__17356),
            .I(N__17329));
    Span4Mux_h I__3232 (
            .O(N__17353),
            .I(N__17326));
    InMux I__3231 (
            .O(N__17350),
            .I(N__17315));
    InMux I__3230 (
            .O(N__17349),
            .I(N__17315));
    InMux I__3229 (
            .O(N__17348),
            .I(N__17315));
    InMux I__3228 (
            .O(N__17347),
            .I(N__17315));
    InMux I__3227 (
            .O(N__17346),
            .I(N__17315));
    InMux I__3226 (
            .O(N__17345),
            .I(N__17312));
    InMux I__3225 (
            .O(N__17344),
            .I(N__17309));
    LocalMux I__3224 (
            .O(N__17335),
            .I(N__17304));
    Span4Mux_h I__3223 (
            .O(N__17332),
            .I(N__17304));
    Span4Mux_h I__3222 (
            .O(N__17329),
            .I(N__17297));
    Span4Mux_h I__3221 (
            .O(N__17326),
            .I(N__17297));
    LocalMux I__3220 (
            .O(N__17315),
            .I(N__17297));
    LocalMux I__3219 (
            .O(N__17312),
            .I(N__17294));
    LocalMux I__3218 (
            .O(N__17309),
            .I(N__17289));
    Span4Mux_v I__3217 (
            .O(N__17304),
            .I(N__17289));
    Span4Mux_v I__3216 (
            .O(N__17297),
            .I(N__17286));
    Odrv12 I__3215 (
            .O(N__17294),
            .I(\tok.n23 ));
    Odrv4 I__3214 (
            .O(N__17289),
            .I(\tok.n23 ));
    Odrv4 I__3213 (
            .O(N__17286),
            .I(\tok.n23 ));
    CEMux I__3212 (
            .O(N__17279),
            .I(N__17276));
    LocalMux I__3211 (
            .O(N__17276),
            .I(N__17272));
    CEMux I__3210 (
            .O(N__17275),
            .I(N__17269));
    Span4Mux_v I__3209 (
            .O(N__17272),
            .I(N__17262));
    LocalMux I__3208 (
            .O(N__17269),
            .I(N__17262));
    CEMux I__3207 (
            .O(N__17268),
            .I(N__17259));
    CEMux I__3206 (
            .O(N__17267),
            .I(N__17256));
    Span4Mux_v I__3205 (
            .O(N__17262),
            .I(N__17253));
    LocalMux I__3204 (
            .O(N__17259),
            .I(N__17249));
    LocalMux I__3203 (
            .O(N__17256),
            .I(N__17246));
    Span4Mux_h I__3202 (
            .O(N__17253),
            .I(N__17243));
    CEMux I__3201 (
            .O(N__17252),
            .I(N__17240));
    Span4Mux_v I__3200 (
            .O(N__17249),
            .I(N__17236));
    Span4Mux_v I__3199 (
            .O(N__17246),
            .I(N__17233));
    Sp12to4 I__3198 (
            .O(N__17243),
            .I(N__17228));
    LocalMux I__3197 (
            .O(N__17240),
            .I(N__17228));
    CEMux I__3196 (
            .O(N__17239),
            .I(N__17225));
    Odrv4 I__3195 (
            .O(N__17236),
            .I(\tok.n950 ));
    Odrv4 I__3194 (
            .O(N__17233),
            .I(\tok.n950 ));
    Odrv12 I__3193 (
            .O(N__17228),
            .I(\tok.n950 ));
    LocalMux I__3192 (
            .O(N__17225),
            .I(\tok.n950 ));
    InMux I__3191 (
            .O(N__17216),
            .I(N__17213));
    LocalMux I__3190 (
            .O(N__17213),
            .I(\tok.n15_adj_847 ));
    CascadeMux I__3189 (
            .O(N__17210),
            .I(N__17207));
    InMux I__3188 (
            .O(N__17207),
            .I(N__17204));
    LocalMux I__3187 (
            .O(N__17204),
            .I(N__17201));
    Span4Mux_h I__3186 (
            .O(N__17201),
            .I(N__17197));
    InMux I__3185 (
            .O(N__17200),
            .I(N__17194));
    Span4Mux_v I__3184 (
            .O(N__17197),
            .I(N__17191));
    LocalMux I__3183 (
            .O(N__17194),
            .I(uart_rx_data_2));
    Odrv4 I__3182 (
            .O(N__17191),
            .I(uart_rx_data_2));
    InMux I__3181 (
            .O(N__17186),
            .I(N__17183));
    LocalMux I__3180 (
            .O(N__17183),
            .I(\tok.n12_adj_843 ));
    InMux I__3179 (
            .O(N__17180),
            .I(N__17177));
    LocalMux I__3178 (
            .O(N__17177),
            .I(N__17174));
    Span4Mux_h I__3177 (
            .O(N__17174),
            .I(N__17169));
    InMux I__3176 (
            .O(N__17173),
            .I(N__17166));
    InMux I__3175 (
            .O(N__17172),
            .I(N__17163));
    Odrv4 I__3174 (
            .O(N__17169),
            .I(capture_1));
    LocalMux I__3173 (
            .O(N__17166),
            .I(capture_1));
    LocalMux I__3172 (
            .O(N__17163),
            .I(capture_1));
    InMux I__3171 (
            .O(N__17156),
            .I(N__17152));
    InMux I__3170 (
            .O(N__17155),
            .I(N__17149));
    LocalMux I__3169 (
            .O(N__17152),
            .I(uart_rx_data_0));
    LocalMux I__3168 (
            .O(N__17149),
            .I(uart_rx_data_0));
    InMux I__3167 (
            .O(N__17144),
            .I(N__17141));
    LocalMux I__3166 (
            .O(N__17141),
            .I(N__17138));
    Span4Mux_h I__3165 (
            .O(N__17138),
            .I(N__17135));
    Odrv4 I__3164 (
            .O(N__17135),
            .I(\tok.table_rd_14 ));
    InMux I__3163 (
            .O(N__17132),
            .I(N__17129));
    LocalMux I__3162 (
            .O(N__17129),
            .I(N__17126));
    Span4Mux_h I__3161 (
            .O(N__17126),
            .I(N__17123));
    Span4Mux_h I__3160 (
            .O(N__17123),
            .I(N__17120));
    Odrv4 I__3159 (
            .O(N__17120),
            .I(\tok.n16_adj_730 ));
    CascadeMux I__3158 (
            .O(N__17117),
            .I(N__17114));
    InMux I__3157 (
            .O(N__17114),
            .I(N__17105));
    InMux I__3156 (
            .O(N__17113),
            .I(N__17100));
    InMux I__3155 (
            .O(N__17112),
            .I(N__17100));
    InMux I__3154 (
            .O(N__17111),
            .I(N__17091));
    InMux I__3153 (
            .O(N__17110),
            .I(N__17091));
    InMux I__3152 (
            .O(N__17109),
            .I(N__17091));
    InMux I__3151 (
            .O(N__17108),
            .I(N__17091));
    LocalMux I__3150 (
            .O(N__17105),
            .I(N__17079));
    LocalMux I__3149 (
            .O(N__17100),
            .I(N__17079));
    LocalMux I__3148 (
            .O(N__17091),
            .I(N__17079));
    InMux I__3147 (
            .O(N__17090),
            .I(N__17074));
    InMux I__3146 (
            .O(N__17089),
            .I(N__17074));
    InMux I__3145 (
            .O(N__17088),
            .I(N__17067));
    InMux I__3144 (
            .O(N__17087),
            .I(N__17067));
    InMux I__3143 (
            .O(N__17086),
            .I(N__17067));
    Span4Mux_s3_v I__3142 (
            .O(N__17079),
            .I(N__17060));
    LocalMux I__3141 (
            .O(N__17074),
            .I(N__17060));
    LocalMux I__3140 (
            .O(N__17067),
            .I(N__17060));
    Span4Mux_h I__3139 (
            .O(N__17060),
            .I(N__17057));
    Odrv4 I__3138 (
            .O(N__17057),
            .I(\tok.n400 ));
    InMux I__3137 (
            .O(N__17054),
            .I(N__17051));
    LocalMux I__3136 (
            .O(N__17051),
            .I(N__17048));
    Span4Mux_v I__3135 (
            .O(N__17048),
            .I(N__17045));
    Span4Mux_h I__3134 (
            .O(N__17045),
            .I(N__17042));
    Sp12to4 I__3133 (
            .O(N__17042),
            .I(N__17039));
    Odrv12 I__3132 (
            .O(N__17039),
            .I(\tok.table_wr_data_0 ));
    InMux I__3131 (
            .O(N__17036),
            .I(N__17033));
    LocalMux I__3130 (
            .O(N__17033),
            .I(\tok.n2614 ));
    CascadeMux I__3129 (
            .O(N__17030),
            .I(\tok.n2614_cascade_ ));
    InMux I__3128 (
            .O(N__17027),
            .I(N__17024));
    LocalMux I__3127 (
            .O(N__17024),
            .I(N__17021));
    Span4Mux_h I__3126 (
            .O(N__17021),
            .I(N__17018));
    Odrv4 I__3125 (
            .O(N__17018),
            .I(\tok.n10_adj_786 ));
    CascadeMux I__3124 (
            .O(N__17015),
            .I(\tok.n6_adj_848_cascade_ ));
    CascadeMux I__3123 (
            .O(N__17012),
            .I(\tok.n32_cascade_ ));
    InMux I__3122 (
            .O(N__17009),
            .I(N__17003));
    InMux I__3121 (
            .O(N__17008),
            .I(N__17003));
    LocalMux I__3120 (
            .O(N__17003),
            .I(uart_rx_data_1));
    InMux I__3119 (
            .O(N__17000),
            .I(N__16997));
    LocalMux I__3118 (
            .O(N__16997),
            .I(N__16994));
    Span4Mux_v I__3117 (
            .O(N__16994),
            .I(N__16991));
    Sp12to4 I__3116 (
            .O(N__16991),
            .I(N__16988));
    Odrv12 I__3115 (
            .O(N__16988),
            .I(\tok.table_wr_data_6 ));
    CascadeMux I__3114 (
            .O(N__16985),
            .I(N__16982));
    InMux I__3113 (
            .O(N__16982),
            .I(N__16976));
    InMux I__3112 (
            .O(N__16981),
            .I(N__16976));
    LocalMux I__3111 (
            .O(N__16976),
            .I(N__16972));
    InMux I__3110 (
            .O(N__16975),
            .I(N__16969));
    Odrv12 I__3109 (
            .O(N__16972),
            .I(capture_2));
    LocalMux I__3108 (
            .O(N__16969),
            .I(capture_2));
    InMux I__3107 (
            .O(N__16964),
            .I(N__16961));
    LocalMux I__3106 (
            .O(N__16961),
            .I(N__16957));
    InMux I__3105 (
            .O(N__16960),
            .I(N__16954));
    Span4Mux_h I__3104 (
            .O(N__16957),
            .I(N__16948));
    LocalMux I__3103 (
            .O(N__16954),
            .I(N__16948));
    InMux I__3102 (
            .O(N__16953),
            .I(N__16945));
    Span4Mux_h I__3101 (
            .O(N__16948),
            .I(N__16939));
    LocalMux I__3100 (
            .O(N__16945),
            .I(N__16936));
    InMux I__3099 (
            .O(N__16944),
            .I(N__16929));
    InMux I__3098 (
            .O(N__16943),
            .I(N__16929));
    InMux I__3097 (
            .O(N__16942),
            .I(N__16929));
    Span4Mux_v I__3096 (
            .O(N__16939),
            .I(N__16923));
    Span4Mux_v I__3095 (
            .O(N__16936),
            .I(N__16917));
    LocalMux I__3094 (
            .O(N__16929),
            .I(N__16917));
    InMux I__3093 (
            .O(N__16928),
            .I(N__16910));
    InMux I__3092 (
            .O(N__16927),
            .I(N__16910));
    InMux I__3091 (
            .O(N__16926),
            .I(N__16910));
    Span4Mux_h I__3090 (
            .O(N__16923),
            .I(N__16907));
    InMux I__3089 (
            .O(N__16922),
            .I(N__16904));
    Span4Mux_h I__3088 (
            .O(N__16917),
            .I(N__16899));
    LocalMux I__3087 (
            .O(N__16910),
            .I(N__16899));
    Odrv4 I__3086 (
            .O(N__16907),
            .I(n4005));
    LocalMux I__3085 (
            .O(N__16904),
            .I(n4005));
    Odrv4 I__3084 (
            .O(N__16899),
            .I(n4005));
    InMux I__3083 (
            .O(N__16892),
            .I(N__16889));
    LocalMux I__3082 (
            .O(N__16889),
            .I(N__16886));
    Span4Mux_v I__3081 (
            .O(N__16886),
            .I(N__16883));
    Span4Mux_h I__3080 (
            .O(N__16883),
            .I(N__16880));
    Sp12to4 I__3079 (
            .O(N__16880),
            .I(N__16877));
    Odrv12 I__3078 (
            .O(N__16877),
            .I(\tok.table_wr_data_2 ));
    CascadeMux I__3077 (
            .O(N__16874),
            .I(\tok.n18_adj_844_cascade_ ));
    InMux I__3076 (
            .O(N__16871),
            .I(N__16868));
    LocalMux I__3075 (
            .O(N__16868),
            .I(N__16865));
    Span12Mux_s10_v I__3074 (
            .O(N__16865),
            .I(N__16862));
    Odrv12 I__3073 (
            .O(N__16862),
            .I(\tok.n16_adj_845 ));
    CascadeMux I__3072 (
            .O(N__16859),
            .I(\tok.n20_adj_846_cascade_ ));
    InMux I__3071 (
            .O(N__16856),
            .I(N__16852));
    InMux I__3070 (
            .O(N__16855),
            .I(N__16849));
    LocalMux I__3069 (
            .O(N__16852),
            .I(\tok.A_15_N_113_2 ));
    LocalMux I__3068 (
            .O(N__16849),
            .I(\tok.A_15_N_113_2 ));
    CascadeMux I__3067 (
            .O(N__16844),
            .I(N__16841));
    InMux I__3066 (
            .O(N__16841),
            .I(N__16838));
    LocalMux I__3065 (
            .O(N__16838),
            .I(N__16835));
    Span4Mux_v I__3064 (
            .O(N__16835),
            .I(N__16832));
    Odrv4 I__3063 (
            .O(N__16832),
            .I(\tok.tc_7 ));
    InMux I__3062 (
            .O(N__16829),
            .I(N__16826));
    LocalMux I__3061 (
            .O(N__16826),
            .I(N__16823));
    Span4Mux_v I__3060 (
            .O(N__16823),
            .I(N__16819));
    InMux I__3059 (
            .O(N__16822),
            .I(N__16816));
    Odrv4 I__3058 (
            .O(N__16819),
            .I(\tok.C_stk.tail_1 ));
    LocalMux I__3057 (
            .O(N__16816),
            .I(\tok.C_stk.tail_1 ));
    CascadeMux I__3056 (
            .O(N__16811),
            .I(\tok.C_stk.n4870_cascade_ ));
    CascadeMux I__3055 (
            .O(N__16808),
            .I(\tok.ram.n4714_cascade_ ));
    InMux I__3054 (
            .O(N__16805),
            .I(N__16802));
    LocalMux I__3053 (
            .O(N__16802),
            .I(N__16798));
    InMux I__3052 (
            .O(N__16801),
            .I(N__16795));
    Span4Mux_s1_v I__3051 (
            .O(N__16798),
            .I(N__16789));
    LocalMux I__3050 (
            .O(N__16795),
            .I(N__16789));
    CascadeMux I__3049 (
            .O(N__16794),
            .I(N__16784));
    Span4Mux_v I__3048 (
            .O(N__16789),
            .I(N__16781));
    InMux I__3047 (
            .O(N__16788),
            .I(N__16774));
    InMux I__3046 (
            .O(N__16787),
            .I(N__16774));
    InMux I__3045 (
            .O(N__16784),
            .I(N__16774));
    Span4Mux_h I__3044 (
            .O(N__16781),
            .I(N__16771));
    LocalMux I__3043 (
            .O(N__16774),
            .I(\tok.c_stk_r_1 ));
    Odrv4 I__3042 (
            .O(N__16771),
            .I(\tok.c_stk_r_1 ));
    InMux I__3041 (
            .O(N__16766),
            .I(N__16763));
    LocalMux I__3040 (
            .O(N__16763),
            .I(N__16760));
    Span4Mux_h I__3039 (
            .O(N__16760),
            .I(N__16757));
    Odrv4 I__3038 (
            .O(N__16757),
            .I(\tok.n4690 ));
    CascadeMux I__3037 (
            .O(N__16754),
            .I(\tok.n1_adj_717_cascade_ ));
    CascadeMux I__3036 (
            .O(N__16751),
            .I(\tok.n5_adj_718_cascade_ ));
    CascadeMux I__3035 (
            .O(N__16748),
            .I(n92_cascade_));
    CascadeMux I__3034 (
            .O(N__16745),
            .I(N__16742));
    InMux I__3033 (
            .O(N__16742),
            .I(N__16739));
    LocalMux I__3032 (
            .O(N__16739),
            .I(N__16736));
    Span4Mux_h I__3031 (
            .O(N__16736),
            .I(N__16733));
    Odrv4 I__3030 (
            .O(N__16733),
            .I(\tok.tc_1 ));
    InMux I__3029 (
            .O(N__16730),
            .I(N__16727));
    LocalMux I__3028 (
            .O(N__16727),
            .I(N__16724));
    Span4Mux_v I__3027 (
            .O(N__16724),
            .I(N__16721));
    Odrv4 I__3026 (
            .O(N__16721),
            .I(\tok.n28_adj_821 ));
    InMux I__3025 (
            .O(N__16718),
            .I(N__16715));
    LocalMux I__3024 (
            .O(N__16715),
            .I(N__16712));
    Span4Mux_v I__3023 (
            .O(N__16712),
            .I(N__16709));
    Span4Mux_h I__3022 (
            .O(N__16709),
            .I(N__16705));
    InMux I__3021 (
            .O(N__16708),
            .I(N__16702));
    Span4Mux_h I__3020 (
            .O(N__16705),
            .I(N__16698));
    LocalMux I__3019 (
            .O(N__16702),
            .I(N__16695));
    InMux I__3018 (
            .O(N__16701),
            .I(N__16692));
    Odrv4 I__3017 (
            .O(N__16698),
            .I(capture_3));
    Odrv12 I__3016 (
            .O(N__16695),
            .I(capture_3));
    LocalMux I__3015 (
            .O(N__16692),
            .I(capture_3));
    CascadeMux I__3014 (
            .O(N__16685),
            .I(N__16682));
    InMux I__3013 (
            .O(N__16682),
            .I(N__16673));
    InMux I__3012 (
            .O(N__16681),
            .I(N__16673));
    InMux I__3011 (
            .O(N__16680),
            .I(N__16673));
    LocalMux I__3010 (
            .O(N__16673),
            .I(\tok.n847 ));
    InMux I__3009 (
            .O(N__16670),
            .I(N__16667));
    LocalMux I__3008 (
            .O(N__16667),
            .I(N__16664));
    Odrv4 I__3007 (
            .O(N__16664),
            .I(\tok.n31 ));
    CascadeMux I__3006 (
            .O(N__16661),
            .I(\tok.C_stk.n4906_cascade_ ));
    CascadeMux I__3005 (
            .O(N__16658),
            .I(\tok.ram.n4699_cascade_ ));
    InMux I__3004 (
            .O(N__16655),
            .I(N__16652));
    LocalMux I__3003 (
            .O(N__16652),
            .I(N__16649));
    Span4Mux_h I__3002 (
            .O(N__16649),
            .I(N__16646));
    Odrv4 I__3001 (
            .O(N__16646),
            .I(\tok.n4649 ));
    CascadeMux I__3000 (
            .O(N__16643),
            .I(\tok.n1_adj_760_cascade_ ));
    CascadeMux I__2999 (
            .O(N__16640),
            .I(\tok.n13_adj_761_cascade_ ));
    CascadeMux I__2998 (
            .O(N__16637),
            .I(\tok.n28_adj_834_cascade_ ));
    CascadeMux I__2997 (
            .O(N__16634),
            .I(\tok.n4604_cascade_ ));
    CascadeMux I__2996 (
            .O(N__16631),
            .I(N__16628));
    InMux I__2995 (
            .O(N__16628),
            .I(N__16625));
    LocalMux I__2994 (
            .O(N__16625),
            .I(N__16622));
    Odrv4 I__2993 (
            .O(N__16622),
            .I(\tok.n34_adj_719 ));
    CascadeMux I__2992 (
            .O(N__16619),
            .I(\tok.n4610_cascade_ ));
    InMux I__2991 (
            .O(N__16616),
            .I(N__16610));
    InMux I__2990 (
            .O(N__16615),
            .I(N__16610));
    LocalMux I__2989 (
            .O(N__16610),
            .I(\tok.n37 ));
    InMux I__2988 (
            .O(N__16607),
            .I(N__16604));
    LocalMux I__2987 (
            .O(N__16604),
            .I(N__16601));
    Span4Mux_h I__2986 (
            .O(N__16601),
            .I(N__16598));
    Span4Mux_v I__2985 (
            .O(N__16598),
            .I(N__16594));
    InMux I__2984 (
            .O(N__16597),
            .I(N__16591));
    Span4Mux_h I__2983 (
            .O(N__16594),
            .I(N__16588));
    LocalMux I__2982 (
            .O(N__16591),
            .I(\tok.table_rd_7 ));
    Odrv4 I__2981 (
            .O(N__16588),
            .I(\tok.table_rd_7 ));
    CascadeMux I__2980 (
            .O(N__16583),
            .I(\tok.n83_adj_796_cascade_ ));
    CascadeMux I__2979 (
            .O(N__16580),
            .I(N__16577));
    InMux I__2978 (
            .O(N__16577),
            .I(N__16573));
    CascadeMux I__2977 (
            .O(N__16576),
            .I(N__16570));
    LocalMux I__2976 (
            .O(N__16573),
            .I(N__16567));
    InMux I__2975 (
            .O(N__16570),
            .I(N__16564));
    Odrv4 I__2974 (
            .O(N__16567),
            .I(\tok.tail_50 ));
    LocalMux I__2973 (
            .O(N__16564),
            .I(\tok.tail_50 ));
    InMux I__2972 (
            .O(N__16559),
            .I(N__16553));
    InMux I__2971 (
            .O(N__16558),
            .I(N__16553));
    LocalMux I__2970 (
            .O(N__16553),
            .I(\tok.C_stk.tail_34 ));
    CascadeMux I__2969 (
            .O(N__16550),
            .I(N__16546));
    CascadeMux I__2968 (
            .O(N__16549),
            .I(N__16543));
    InMux I__2967 (
            .O(N__16546),
            .I(N__16540));
    InMux I__2966 (
            .O(N__16543),
            .I(N__16537));
    LocalMux I__2965 (
            .O(N__16540),
            .I(\tok.tail_42 ));
    LocalMux I__2964 (
            .O(N__16537),
            .I(\tok.tail_42 ));
    InMux I__2963 (
            .O(N__16532),
            .I(N__16526));
    InMux I__2962 (
            .O(N__16531),
            .I(N__16526));
    LocalMux I__2961 (
            .O(N__16526),
            .I(\tok.tail_28 ));
    CascadeMux I__2960 (
            .O(N__16523),
            .I(\tok.n127_cascade_ ));
    InMux I__2959 (
            .O(N__16520),
            .I(N__16517));
    LocalMux I__2958 (
            .O(N__16517),
            .I(N__16513));
    InMux I__2957 (
            .O(N__16516),
            .I(N__16510));
    Odrv12 I__2956 (
            .O(N__16513),
            .I(\tok.n4446 ));
    LocalMux I__2955 (
            .O(N__16510),
            .I(\tok.n4446 ));
    CascadeMux I__2954 (
            .O(N__16505),
            .I(\tok.n4394_cascade_ ));
    CascadeMux I__2953 (
            .O(N__16502),
            .I(\tok.n27_adj_863_cascade_ ));
    CascadeMux I__2952 (
            .O(N__16499),
            .I(\tok.n27_adj_865_cascade_ ));
    InMux I__2951 (
            .O(N__16496),
            .I(N__16493));
    LocalMux I__2950 (
            .O(N__16493),
            .I(\tok.n27_adj_664 ));
    InMux I__2949 (
            .O(N__16490),
            .I(N__16487));
    LocalMux I__2948 (
            .O(N__16487),
            .I(N__16484));
    Span4Mux_s3_v I__2947 (
            .O(N__16484),
            .I(N__16481));
    Odrv4 I__2946 (
            .O(N__16481),
            .I(\tok.n27_adj_866 ));
    InMux I__2945 (
            .O(N__16478),
            .I(N__16475));
    LocalMux I__2944 (
            .O(N__16475),
            .I(\tok.uart.sender_6 ));
    InMux I__2943 (
            .O(N__16472),
            .I(N__16456));
    InMux I__2942 (
            .O(N__16471),
            .I(N__16456));
    InMux I__2941 (
            .O(N__16470),
            .I(N__16456));
    InMux I__2940 (
            .O(N__16469),
            .I(N__16456));
    InMux I__2939 (
            .O(N__16468),
            .I(N__16449));
    InMux I__2938 (
            .O(N__16467),
            .I(N__16449));
    InMux I__2937 (
            .O(N__16466),
            .I(N__16449));
    SRMux I__2936 (
            .O(N__16465),
            .I(N__16444));
    LocalMux I__2935 (
            .O(N__16456),
            .I(N__16439));
    LocalMux I__2934 (
            .O(N__16449),
            .I(N__16439));
    InMux I__2933 (
            .O(N__16448),
            .I(N__16434));
    InMux I__2932 (
            .O(N__16447),
            .I(N__16434));
    LocalMux I__2931 (
            .O(N__16444),
            .I(N__16431));
    Span4Mux_v I__2930 (
            .O(N__16439),
            .I(N__16428));
    LocalMux I__2929 (
            .O(N__16434),
            .I(N__16424));
    Span4Mux_v I__2928 (
            .O(N__16431),
            .I(N__16420));
    Span4Mux_h I__2927 (
            .O(N__16428),
            .I(N__16417));
    InMux I__2926 (
            .O(N__16427),
            .I(N__16414));
    Span4Mux_h I__2925 (
            .O(N__16424),
            .I(N__16411));
    InMux I__2924 (
            .O(N__16423),
            .I(N__16408));
    Odrv4 I__2923 (
            .O(N__16420),
            .I(n23));
    Odrv4 I__2922 (
            .O(N__16417),
            .I(n23));
    LocalMux I__2921 (
            .O(N__16414),
            .I(n23));
    Odrv4 I__2920 (
            .O(N__16411),
            .I(n23));
    LocalMux I__2919 (
            .O(N__16408),
            .I(n23));
    InMux I__2918 (
            .O(N__16397),
            .I(N__16394));
    LocalMux I__2917 (
            .O(N__16394),
            .I(N__16391));
    Odrv4 I__2916 (
            .O(N__16391),
            .I(\tok.uart.sender_5 ));
    CEMux I__2915 (
            .O(N__16388),
            .I(N__16383));
    CEMux I__2914 (
            .O(N__16387),
            .I(N__16380));
    CEMux I__2913 (
            .O(N__16386),
            .I(N__16377));
    LocalMux I__2912 (
            .O(N__16383),
            .I(N__16374));
    LocalMux I__2911 (
            .O(N__16380),
            .I(N__16371));
    LocalMux I__2910 (
            .O(N__16377),
            .I(N__16368));
    Span4Mux_h I__2909 (
            .O(N__16374),
            .I(N__16364));
    Span4Mux_h I__2908 (
            .O(N__16371),
            .I(N__16359));
    Span4Mux_s3_v I__2907 (
            .O(N__16368),
            .I(N__16359));
    CEMux I__2906 (
            .O(N__16367),
            .I(N__16356));
    Span4Mux_h I__2905 (
            .O(N__16364),
            .I(N__16353));
    Span4Mux_v I__2904 (
            .O(N__16359),
            .I(N__16348));
    LocalMux I__2903 (
            .O(N__16356),
            .I(N__16348));
    Span4Mux_s1_h I__2902 (
            .O(N__16353),
            .I(N__16345));
    Span4Mux_h I__2901 (
            .O(N__16348),
            .I(N__16342));
    Odrv4 I__2900 (
            .O(N__16345),
            .I(\tok.uart.n964 ));
    Odrv4 I__2899 (
            .O(N__16342),
            .I(\tok.uart.n964 ));
    InMux I__2898 (
            .O(N__16337),
            .I(N__16334));
    LocalMux I__2897 (
            .O(N__16334),
            .I(N__16331));
    Span4Mux_v I__2896 (
            .O(N__16331),
            .I(N__16328));
    Odrv4 I__2895 (
            .O(N__16328),
            .I(\tok.n16_adj_706 ));
    InMux I__2894 (
            .O(N__16325),
            .I(N__16322));
    LocalMux I__2893 (
            .O(N__16322),
            .I(\tok.n14_adj_707 ));
    CascadeMux I__2892 (
            .O(N__16319),
            .I(\tok.n20_adj_708_cascade_ ));
    CascadeMux I__2891 (
            .O(N__16316),
            .I(\tok.n22_adj_709_cascade_ ));
    InMux I__2890 (
            .O(N__16313),
            .I(N__16310));
    LocalMux I__2889 (
            .O(N__16310),
            .I(\tok.A_15_N_113_5 ));
    InMux I__2888 (
            .O(N__16307),
            .I(N__16304));
    LocalMux I__2887 (
            .O(N__16304),
            .I(N__16301));
    Span4Mux_v I__2886 (
            .O(N__16301),
            .I(N__16298));
    Odrv4 I__2885 (
            .O(N__16298),
            .I(\tok.n10_adj_806 ));
    CascadeMux I__2884 (
            .O(N__16295),
            .I(\tok.n13_adj_813_cascade_ ));
    InMux I__2883 (
            .O(N__16292),
            .I(N__16289));
    LocalMux I__2882 (
            .O(N__16289),
            .I(\tok.n18_adj_819 ));
    InMux I__2881 (
            .O(N__16286),
            .I(N__16283));
    LocalMux I__2880 (
            .O(N__16283),
            .I(\tok.n15_adj_823 ));
    InMux I__2879 (
            .O(N__16280),
            .I(N__16277));
    LocalMux I__2878 (
            .O(N__16277),
            .I(\tok.uart.sender_3 ));
    InMux I__2877 (
            .O(N__16274),
            .I(N__16271));
    LocalMux I__2876 (
            .O(N__16271),
            .I(\tok.A_0 ));
    CascadeMux I__2875 (
            .O(N__16268),
            .I(N__16265));
    InMux I__2874 (
            .O(N__16265),
            .I(N__16262));
    LocalMux I__2873 (
            .O(N__16262),
            .I(N__16259));
    Odrv12 I__2872 (
            .O(N__16259),
            .I(sender_2));
    InMux I__2871 (
            .O(N__16256),
            .I(N__16253));
    LocalMux I__2870 (
            .O(N__16253),
            .I(N__16250));
    Odrv4 I__2869 (
            .O(N__16250),
            .I(\tok.A_2 ));
    InMux I__2868 (
            .O(N__16247),
            .I(N__16244));
    LocalMux I__2867 (
            .O(N__16244),
            .I(\tok.uart.sender_4 ));
    InMux I__2866 (
            .O(N__16241),
            .I(N__16238));
    LocalMux I__2865 (
            .O(N__16238),
            .I(N__16235));
    Span4Mux_h I__2864 (
            .O(N__16235),
            .I(N__16232));
    Odrv4 I__2863 (
            .O(N__16232),
            .I(\tok.n10_adj_783 ));
    CascadeMux I__2862 (
            .O(N__16229),
            .I(\tok.n14_adj_779_cascade_ ));
    InMux I__2861 (
            .O(N__16226),
            .I(N__16223));
    LocalMux I__2860 (
            .O(N__16223),
            .I(N__16220));
    Span4Mux_h I__2859 (
            .O(N__16220),
            .I(N__16217));
    Odrv4 I__2858 (
            .O(N__16217),
            .I(\tok.n20_adj_781 ));
    CascadeMux I__2857 (
            .O(N__16214),
            .I(\tok.n22_adj_784_cascade_ ));
    CascadeMux I__2856 (
            .O(N__16211),
            .I(\tok.A_15_N_113_6_cascade_ ));
    CascadeMux I__2855 (
            .O(N__16208),
            .I(\tok.A_6_cascade_ ));
    InMux I__2854 (
            .O(N__16205),
            .I(N__16202));
    LocalMux I__2853 (
            .O(N__16202),
            .I(N__16199));
    Span4Mux_h I__2852 (
            .O(N__16199),
            .I(N__16196));
    Span4Mux_v I__2851 (
            .O(N__16196),
            .I(N__16193));
    Span4Mux_h I__2850 (
            .O(N__16193),
            .I(N__16190));
    Odrv4 I__2849 (
            .O(N__16190),
            .I(\tok.uart.sender_9 ));
    InMux I__2848 (
            .O(N__16187),
            .I(N__16184));
    LocalMux I__2847 (
            .O(N__16184),
            .I(\tok.uart.sender_8 ));
    InMux I__2846 (
            .O(N__16181),
            .I(N__16178));
    LocalMux I__2845 (
            .O(N__16178),
            .I(\tok.A_5 ));
    InMux I__2844 (
            .O(N__16175),
            .I(N__16172));
    LocalMux I__2843 (
            .O(N__16172),
            .I(\tok.uart.sender_7 ));
    InMux I__2842 (
            .O(N__16169),
            .I(N__16166));
    LocalMux I__2841 (
            .O(N__16166),
            .I(\tok.n2 ));
    CascadeMux I__2840 (
            .O(N__16163),
            .I(\tok.n19_cascade_ ));
    InMux I__2839 (
            .O(N__16160),
            .I(N__16157));
    LocalMux I__2838 (
            .O(N__16157),
            .I(N__16154));
    Span4Mux_h I__2837 (
            .O(N__16154),
            .I(N__16151));
    Odrv4 I__2836 (
            .O(N__16151),
            .I(\tok.n6_adj_684 ));
    CascadeMux I__2835 (
            .O(N__16148),
            .I(\tok.n22_adj_683_cascade_ ));
    InMux I__2834 (
            .O(N__16145),
            .I(N__16142));
    LocalMux I__2833 (
            .O(N__16142),
            .I(\tok.n4544 ));
    CascadeMux I__2832 (
            .O(N__16139),
            .I(\tok.A_15_N_113_0_cascade_ ));
    InMux I__2831 (
            .O(N__16136),
            .I(N__16133));
    LocalMux I__2830 (
            .O(N__16133),
            .I(\tok.n4520 ));
    CascadeMux I__2829 (
            .O(N__16130),
            .I(\tok.n46_cascade_ ));
    InMux I__2828 (
            .O(N__16127),
            .I(N__16124));
    LocalMux I__2827 (
            .O(N__16124),
            .I(N__16121));
    Odrv4 I__2826 (
            .O(N__16121),
            .I(\tok.A_15_N_113_1 ));
    CascadeMux I__2825 (
            .O(N__16118),
            .I(\tok.A_15_N_113_1_cascade_ ));
    CascadeMux I__2824 (
            .O(N__16115),
            .I(\tok.A_1_cascade_ ));
    CascadeMux I__2823 (
            .O(N__16112),
            .I(\tok.A__15__N_129_cascade_ ));
    CascadeMux I__2822 (
            .O(N__16109),
            .I(\tok.n27_adj_867_cascade_ ));
    CascadeMux I__2821 (
            .O(N__16106),
            .I(N__16103));
    InMux I__2820 (
            .O(N__16103),
            .I(N__16100));
    LocalMux I__2819 (
            .O(N__16100),
            .I(\tok.n1 ));
    CascadeMux I__2818 (
            .O(N__16097),
            .I(\tok.n14_adj_678_cascade_ ));
    InMux I__2817 (
            .O(N__16094),
            .I(N__16091));
    LocalMux I__2816 (
            .O(N__16091),
            .I(\tok.n18_adj_859 ));
    InMux I__2815 (
            .O(N__16088),
            .I(N__16085));
    LocalMux I__2814 (
            .O(N__16085),
            .I(N__16082));
    Odrv4 I__2813 (
            .O(N__16082),
            .I(\tok.n22_adj_855 ));
    InMux I__2812 (
            .O(N__16079),
            .I(N__16076));
    LocalMux I__2811 (
            .O(N__16076),
            .I(N__16072));
    InMux I__2810 (
            .O(N__16075),
            .I(N__16069));
    Span4Mux_h I__2809 (
            .O(N__16072),
            .I(N__16066));
    LocalMux I__2808 (
            .O(N__16069),
            .I(\tok.n880 ));
    Odrv4 I__2807 (
            .O(N__16066),
            .I(\tok.n880 ));
    CascadeMux I__2806 (
            .O(N__16061),
            .I(\tok.n23_cascade_ ));
    InMux I__2805 (
            .O(N__16058),
            .I(N__16055));
    LocalMux I__2804 (
            .O(N__16055),
            .I(\tok.n23_adj_856 ));
    CascadeMux I__2803 (
            .O(N__16052),
            .I(N__16043));
    CascadeMux I__2802 (
            .O(N__16051),
            .I(N__16040));
    InMux I__2801 (
            .O(N__16050),
            .I(N__16034));
    InMux I__2800 (
            .O(N__16049),
            .I(N__16034));
    InMux I__2799 (
            .O(N__16048),
            .I(N__16025));
    InMux I__2798 (
            .O(N__16047),
            .I(N__16025));
    InMux I__2797 (
            .O(N__16046),
            .I(N__16025));
    InMux I__2796 (
            .O(N__16043),
            .I(N__16025));
    InMux I__2795 (
            .O(N__16040),
            .I(N__16020));
    InMux I__2794 (
            .O(N__16039),
            .I(N__16020));
    LocalMux I__2793 (
            .O(N__16034),
            .I(N__16015));
    LocalMux I__2792 (
            .O(N__16025),
            .I(N__16015));
    LocalMux I__2791 (
            .O(N__16020),
            .I(\tok.n64 ));
    Odrv12 I__2790 (
            .O(N__16015),
            .I(\tok.n64 ));
    InMux I__2789 (
            .O(N__16010),
            .I(N__16003));
    InMux I__2788 (
            .O(N__16009),
            .I(N__16003));
    InMux I__2787 (
            .O(N__16008),
            .I(N__15998));
    LocalMux I__2786 (
            .O(N__16003),
            .I(N__15995));
    InMux I__2785 (
            .O(N__16002),
            .I(N__15990));
    InMux I__2784 (
            .O(N__16001),
            .I(N__15990));
    LocalMux I__2783 (
            .O(N__15998),
            .I(\tok.n1_adj_802 ));
    Odrv4 I__2782 (
            .O(N__15995),
            .I(\tok.n1_adj_802 ));
    LocalMux I__2781 (
            .O(N__15990),
            .I(\tok.n1_adj_802 ));
    InMux I__2780 (
            .O(N__15983),
            .I(N__15980));
    LocalMux I__2779 (
            .O(N__15980),
            .I(N__15977));
    Odrv12 I__2778 (
            .O(N__15977),
            .I(\tok.depth_2 ));
    CascadeMux I__2777 (
            .O(N__15974),
            .I(\tok.depth_0_cascade_ ));
    InMux I__2776 (
            .O(N__15971),
            .I(N__15968));
    LocalMux I__2775 (
            .O(N__15968),
            .I(N__15965));
    Odrv12 I__2774 (
            .O(N__15965),
            .I(\tok.n6_adj_853 ));
    InMux I__2773 (
            .O(N__15962),
            .I(N__15956));
    InMux I__2772 (
            .O(N__15961),
            .I(N__15956));
    LocalMux I__2771 (
            .O(N__15956),
            .I(\tok.n6_adj_832 ));
    InMux I__2770 (
            .O(N__15953),
            .I(N__15950));
    LocalMux I__2769 (
            .O(N__15950),
            .I(\tok.n4504 ));
    CascadeMux I__2768 (
            .O(N__15947),
            .I(\tok.n4432_cascade_ ));
    CascadeMux I__2767 (
            .O(N__15944),
            .I(N__15936));
    InMux I__2766 (
            .O(N__15943),
            .I(N__15931));
    InMux I__2765 (
            .O(N__15942),
            .I(N__15931));
    InMux I__2764 (
            .O(N__15941),
            .I(N__15928));
    InMux I__2763 (
            .O(N__15940),
            .I(N__15921));
    InMux I__2762 (
            .O(N__15939),
            .I(N__15921));
    InMux I__2761 (
            .O(N__15936),
            .I(N__15921));
    LocalMux I__2760 (
            .O(N__15931),
            .I(\tok.A_stk_delta_1__N_4 ));
    LocalMux I__2759 (
            .O(N__15928),
            .I(\tok.A_stk_delta_1__N_4 ));
    LocalMux I__2758 (
            .O(N__15921),
            .I(\tok.A_stk_delta_1__N_4 ));
    CascadeMux I__2757 (
            .O(N__15914),
            .I(\tok.n1_adj_802_cascade_ ));
    InMux I__2756 (
            .O(N__15911),
            .I(N__15902));
    InMux I__2755 (
            .O(N__15910),
            .I(N__15902));
    InMux I__2754 (
            .O(N__15909),
            .I(N__15902));
    LocalMux I__2753 (
            .O(N__15902),
            .I(\tok.n189 ));
    CascadeMux I__2752 (
            .O(N__15899),
            .I(N__15891));
    InMux I__2751 (
            .O(N__15898),
            .I(N__15886));
    InMux I__2750 (
            .O(N__15897),
            .I(N__15879));
    InMux I__2749 (
            .O(N__15896),
            .I(N__15879));
    InMux I__2748 (
            .O(N__15895),
            .I(N__15879));
    InMux I__2747 (
            .O(N__15894),
            .I(N__15870));
    InMux I__2746 (
            .O(N__15891),
            .I(N__15870));
    InMux I__2745 (
            .O(N__15890),
            .I(N__15870));
    InMux I__2744 (
            .O(N__15889),
            .I(N__15870));
    LocalMux I__2743 (
            .O(N__15886),
            .I(\tok.n62 ));
    LocalMux I__2742 (
            .O(N__15879),
            .I(\tok.n62 ));
    LocalMux I__2741 (
            .O(N__15870),
            .I(\tok.n62 ));
    CascadeMux I__2740 (
            .O(N__15863),
            .I(\tok.n189_cascade_ ));
    InMux I__2739 (
            .O(N__15860),
            .I(N__15853));
    InMux I__2738 (
            .O(N__15859),
            .I(N__15853));
    InMux I__2737 (
            .O(N__15858),
            .I(N__15850));
    LocalMux I__2736 (
            .O(N__15853),
            .I(\tok.n4_adj_809 ));
    LocalMux I__2735 (
            .O(N__15850),
            .I(\tok.n4_adj_809 ));
    CascadeMux I__2734 (
            .O(N__15845),
            .I(\tok.n27_adj_793_cascade_ ));
    InMux I__2733 (
            .O(N__15842),
            .I(N__15839));
    LocalMux I__2732 (
            .O(N__15839),
            .I(\tok.n25_adj_794 ));
    InMux I__2731 (
            .O(N__15836),
            .I(N__15833));
    LocalMux I__2730 (
            .O(N__15833),
            .I(\tok.n26_adj_792 ));
    InMux I__2729 (
            .O(N__15830),
            .I(N__15827));
    LocalMux I__2728 (
            .O(N__15827),
            .I(\tok.n28_adj_791 ));
    CascadeMux I__2727 (
            .O(N__15824),
            .I(N__15820));
    CascadeMux I__2726 (
            .O(N__15823),
            .I(N__15814));
    InMux I__2725 (
            .O(N__15820),
            .I(N__15808));
    InMux I__2724 (
            .O(N__15819),
            .I(N__15808));
    InMux I__2723 (
            .O(N__15818),
            .I(N__15803));
    InMux I__2722 (
            .O(N__15817),
            .I(N__15803));
    InMux I__2721 (
            .O(N__15814),
            .I(N__15798));
    InMux I__2720 (
            .O(N__15813),
            .I(N__15798));
    LocalMux I__2719 (
            .O(N__15808),
            .I(\tok.n63 ));
    LocalMux I__2718 (
            .O(N__15803),
            .I(\tok.n63 ));
    LocalMux I__2717 (
            .O(N__15798),
            .I(\tok.n63 ));
    CascadeMux I__2716 (
            .O(N__15791),
            .I(\tok.A_stk_delta_1__N_4_cascade_ ));
    InMux I__2715 (
            .O(N__15788),
            .I(N__15778));
    InMux I__2714 (
            .O(N__15787),
            .I(N__15778));
    InMux I__2713 (
            .O(N__15786),
            .I(N__15771));
    InMux I__2712 (
            .O(N__15785),
            .I(N__15771));
    InMux I__2711 (
            .O(N__15784),
            .I(N__15771));
    InMux I__2710 (
            .O(N__15783),
            .I(N__15768));
    LocalMux I__2709 (
            .O(N__15778),
            .I(\tok.n61 ));
    LocalMux I__2708 (
            .O(N__15771),
            .I(\tok.n61 ));
    LocalMux I__2707 (
            .O(N__15768),
            .I(\tok.n61 ));
    CascadeMux I__2706 (
            .O(N__15761),
            .I(\tok.n4_adj_809_cascade_ ));
    CascadeMux I__2705 (
            .O(N__15758),
            .I(\tok.depth_3_cascade_ ));
    InMux I__2704 (
            .O(N__15755),
            .I(N__15752));
    LocalMux I__2703 (
            .O(N__15752),
            .I(\tok.depth_1 ));
    CascadeMux I__2702 (
            .O(N__15749),
            .I(\tok.n4554_cascade_ ));
    InMux I__2701 (
            .O(N__15746),
            .I(N__15736));
    InMux I__2700 (
            .O(N__15745),
            .I(N__15733));
    InMux I__2699 (
            .O(N__15744),
            .I(N__15728));
    InMux I__2698 (
            .O(N__15743),
            .I(N__15725));
    InMux I__2697 (
            .O(N__15742),
            .I(N__15721));
    InMux I__2696 (
            .O(N__15741),
            .I(N__15716));
    InMux I__2695 (
            .O(N__15740),
            .I(N__15713));
    InMux I__2694 (
            .O(N__15739),
            .I(N__15709));
    LocalMux I__2693 (
            .O(N__15736),
            .I(N__15706));
    LocalMux I__2692 (
            .O(N__15733),
            .I(N__15703));
    InMux I__2691 (
            .O(N__15732),
            .I(N__15700));
    InMux I__2690 (
            .O(N__15731),
            .I(N__15697));
    LocalMux I__2689 (
            .O(N__15728),
            .I(N__15692));
    LocalMux I__2688 (
            .O(N__15725),
            .I(N__15692));
    InMux I__2687 (
            .O(N__15724),
            .I(N__15689));
    LocalMux I__2686 (
            .O(N__15721),
            .I(N__15686));
    InMux I__2685 (
            .O(N__15720),
            .I(N__15683));
    InMux I__2684 (
            .O(N__15719),
            .I(N__15678));
    LocalMux I__2683 (
            .O(N__15716),
            .I(N__15673));
    LocalMux I__2682 (
            .O(N__15713),
            .I(N__15673));
    InMux I__2681 (
            .O(N__15712),
            .I(N__15670));
    LocalMux I__2680 (
            .O(N__15709),
            .I(N__15667));
    Span4Mux_s3_h I__2679 (
            .O(N__15706),
            .I(N__15658));
    Span4Mux_v I__2678 (
            .O(N__15703),
            .I(N__15658));
    LocalMux I__2677 (
            .O(N__15700),
            .I(N__15658));
    LocalMux I__2676 (
            .O(N__15697),
            .I(N__15658));
    Span4Mux_s3_h I__2675 (
            .O(N__15692),
            .I(N__15653));
    LocalMux I__2674 (
            .O(N__15689),
            .I(N__15653));
    Span4Mux_v I__2673 (
            .O(N__15686),
            .I(N__15650));
    LocalMux I__2672 (
            .O(N__15683),
            .I(N__15647));
    InMux I__2671 (
            .O(N__15682),
            .I(N__15644));
    InMux I__2670 (
            .O(N__15681),
            .I(N__15641));
    LocalMux I__2669 (
            .O(N__15678),
            .I(N__15638));
    Span12Mux_s7_h I__2668 (
            .O(N__15673),
            .I(N__15635));
    LocalMux I__2667 (
            .O(N__15670),
            .I(N__15632));
    Span4Mux_h I__2666 (
            .O(N__15667),
            .I(N__15627));
    Span4Mux_h I__2665 (
            .O(N__15658),
            .I(N__15627));
    Span4Mux_h I__2664 (
            .O(N__15653),
            .I(N__15624));
    Span4Mux_h I__2663 (
            .O(N__15650),
            .I(N__15615));
    Span4Mux_v I__2662 (
            .O(N__15647),
            .I(N__15615));
    LocalMux I__2661 (
            .O(N__15644),
            .I(N__15615));
    LocalMux I__2660 (
            .O(N__15641),
            .I(N__15615));
    Odrv12 I__2659 (
            .O(N__15638),
            .I(\tok.n237 ));
    Odrv12 I__2658 (
            .O(N__15635),
            .I(\tok.n237 ));
    Odrv4 I__2657 (
            .O(N__15632),
            .I(\tok.n237 ));
    Odrv4 I__2656 (
            .O(N__15627),
            .I(\tok.n237 ));
    Odrv4 I__2655 (
            .O(N__15624),
            .I(\tok.n237 ));
    Odrv4 I__2654 (
            .O(N__15615),
            .I(\tok.n237 ));
    CascadeMux I__2653 (
            .O(N__15602),
            .I(\tok.n875_cascade_ ));
    InMux I__2652 (
            .O(N__15599),
            .I(N__15594));
    InMux I__2651 (
            .O(N__15598),
            .I(N__15591));
    InMux I__2650 (
            .O(N__15597),
            .I(N__15588));
    LocalMux I__2649 (
            .O(N__15594),
            .I(N__15585));
    LocalMux I__2648 (
            .O(N__15591),
            .I(\tok.n2562 ));
    LocalMux I__2647 (
            .O(N__15588),
            .I(\tok.n2562 ));
    Odrv4 I__2646 (
            .O(N__15585),
            .I(\tok.n2562 ));
    InMux I__2645 (
            .O(N__15578),
            .I(N__15572));
    InMux I__2644 (
            .O(N__15577),
            .I(N__15572));
    LocalMux I__2643 (
            .O(N__15572),
            .I(\tok.n2503 ));
    CascadeMux I__2642 (
            .O(N__15569),
            .I(\tok.n2562_cascade_ ));
    CascadeMux I__2641 (
            .O(N__15566),
            .I(\tok.n4474_cascade_ ));
    InMux I__2640 (
            .O(N__15563),
            .I(N__15560));
    LocalMux I__2639 (
            .O(N__15560),
            .I(\tok.n875 ));
    CascadeMux I__2638 (
            .O(N__15557),
            .I(\tok.n20_adj_772_cascade_ ));
    InMux I__2637 (
            .O(N__15554),
            .I(N__15548));
    InMux I__2636 (
            .O(N__15553),
            .I(N__15548));
    LocalMux I__2635 (
            .O(N__15548),
            .I(\tok.tail_9 ));
    InMux I__2634 (
            .O(N__15545),
            .I(N__15539));
    InMux I__2633 (
            .O(N__15544),
            .I(N__15539));
    LocalMux I__2632 (
            .O(N__15539),
            .I(\tok.C_stk.tail_17 ));
    CascadeMux I__2631 (
            .O(N__15536),
            .I(N__15533));
    InMux I__2630 (
            .O(N__15533),
            .I(N__15527));
    InMux I__2629 (
            .O(N__15532),
            .I(N__15527));
    LocalMux I__2628 (
            .O(N__15527),
            .I(N__15524));
    Odrv4 I__2627 (
            .O(N__15524),
            .I(\tok.tail_25 ));
    InMux I__2626 (
            .O(N__15521),
            .I(N__15515));
    InMux I__2625 (
            .O(N__15520),
            .I(N__15515));
    LocalMux I__2624 (
            .O(N__15515),
            .I(\tok.C_stk.tail_33 ));
    InMux I__2623 (
            .O(N__15512),
            .I(N__15508));
    InMux I__2622 (
            .O(N__15511),
            .I(N__15505));
    LocalMux I__2621 (
            .O(N__15508),
            .I(\tok.tail_57 ));
    LocalMux I__2620 (
            .O(N__15505),
            .I(\tok.tail_57 ));
    InMux I__2619 (
            .O(N__15500),
            .I(N__15494));
    InMux I__2618 (
            .O(N__15499),
            .I(N__15494));
    LocalMux I__2617 (
            .O(N__15494),
            .I(\tok.tail_41 ));
    InMux I__2616 (
            .O(N__15491),
            .I(N__15487));
    InMux I__2615 (
            .O(N__15490),
            .I(N__15484));
    LocalMux I__2614 (
            .O(N__15487),
            .I(\tok.tail_49 ));
    LocalMux I__2613 (
            .O(N__15484),
            .I(\tok.tail_49 ));
    InMux I__2612 (
            .O(N__15479),
            .I(N__15475));
    InMux I__2611 (
            .O(N__15478),
            .I(N__15472));
    LocalMux I__2610 (
            .O(N__15475),
            .I(\tok.tail_58 ));
    LocalMux I__2609 (
            .O(N__15472),
            .I(\tok.tail_58 ));
    InMux I__2608 (
            .O(N__15467),
            .I(N__15464));
    LocalMux I__2607 (
            .O(N__15464),
            .I(N__15461));
    Odrv4 I__2606 (
            .O(N__15461),
            .I(\tok.n16_adj_820 ));
    CascadeMux I__2605 (
            .O(N__15458),
            .I(\tok.n20_adj_822_cascade_ ));
    CascadeMux I__2604 (
            .O(N__15455),
            .I(\tok.A_15_N_113_5_cascade_ ));
    InMux I__2603 (
            .O(N__15452),
            .I(N__15449));
    LocalMux I__2602 (
            .O(N__15449),
            .I(N__15446));
    Span4Mux_v I__2601 (
            .O(N__15446),
            .I(N__15443));
    Odrv4 I__2600 (
            .O(N__15443),
            .I(\tok.n297 ));
    CascadeMux I__2599 (
            .O(N__15440),
            .I(N__15437));
    InMux I__2598 (
            .O(N__15437),
            .I(N__15434));
    LocalMux I__2597 (
            .O(N__15434),
            .I(\tok.n208 ));
    InMux I__2596 (
            .O(N__15431),
            .I(N__15428));
    LocalMux I__2595 (
            .O(N__15428),
            .I(N__15425));
    Span4Mux_v I__2594 (
            .O(N__15425),
            .I(N__15422));
    Odrv4 I__2593 (
            .O(N__15422),
            .I(\tok.n20_adj_858 ));
    InMux I__2592 (
            .O(N__15419),
            .I(N__15416));
    LocalMux I__2591 (
            .O(N__15416),
            .I(N__15413));
    Span4Mux_h I__2590 (
            .O(N__15413),
            .I(N__15410));
    Odrv4 I__2589 (
            .O(N__15410),
            .I(\tok.n299 ));
    CascadeMux I__2588 (
            .O(N__15407),
            .I(\tok.n27_adj_644_cascade_ ));
    CascadeMux I__2587 (
            .O(N__15404),
            .I(\tok.n2_adj_720_cascade_ ));
    InMux I__2586 (
            .O(N__15401),
            .I(N__15398));
    LocalMux I__2585 (
            .O(N__15398),
            .I(\tok.n14_adj_722 ));
    InMux I__2584 (
            .O(N__15395),
            .I(N__15392));
    LocalMux I__2583 (
            .O(N__15392),
            .I(N__15389));
    Span12Mux_s11_v I__2582 (
            .O(N__15389),
            .I(N__15386));
    Odrv12 I__2581 (
            .O(N__15386),
            .I(\tok.n6_adj_731 ));
    CascadeMux I__2580 (
            .O(N__15383),
            .I(\tok.n13_adj_726_cascade_ ));
    InMux I__2579 (
            .O(N__15380),
            .I(N__15377));
    LocalMux I__2578 (
            .O(N__15377),
            .I(N__15374));
    Odrv12 I__2577 (
            .O(N__15374),
            .I(\tok.n12_adj_723 ));
    InMux I__2576 (
            .O(N__15371),
            .I(N__15368));
    LocalMux I__2575 (
            .O(N__15368),
            .I(N__15365));
    Span4Mux_v I__2574 (
            .O(N__15365),
            .I(N__15362));
    Odrv4 I__2573 (
            .O(N__15362),
            .I(\tok.n4661 ));
    CascadeMux I__2572 (
            .O(N__15359),
            .I(\tok.n20_adj_732_cascade_ ));
    InMux I__2571 (
            .O(N__15356),
            .I(N__15353));
    LocalMux I__2570 (
            .O(N__15353),
            .I(N__15350));
    Odrv12 I__2569 (
            .O(N__15350),
            .I(\tok.n4658 ));
    InMux I__2568 (
            .O(N__15347),
            .I(N__15344));
    LocalMux I__2567 (
            .O(N__15344),
            .I(\tok.n9_adj_728 ));
    InMux I__2566 (
            .O(N__15341),
            .I(N__15338));
    LocalMux I__2565 (
            .O(N__15338),
            .I(N__15335));
    Span4Mux_v I__2564 (
            .O(N__15335),
            .I(N__15332));
    Odrv4 I__2563 (
            .O(N__15332),
            .I(\tok.n184 ));
    CascadeMux I__2562 (
            .O(N__15329),
            .I(N__15326));
    InMux I__2561 (
            .O(N__15326),
            .I(N__15323));
    LocalMux I__2560 (
            .O(N__15323),
            .I(N__15319));
    InMux I__2559 (
            .O(N__15322),
            .I(N__15316));
    Span4Mux_h I__2558 (
            .O(N__15319),
            .I(N__15313));
    LocalMux I__2557 (
            .O(N__15316),
            .I(uart_rx_data_5));
    Odrv4 I__2556 (
            .O(N__15313),
            .I(uart_rx_data_5));
    CascadeMux I__2555 (
            .O(N__15308),
            .I(\tok.n12_adj_815_cascade_ ));
    InMux I__2554 (
            .O(N__15305),
            .I(N__15302));
    LocalMux I__2553 (
            .O(N__15302),
            .I(\tok.n4653 ));
    InMux I__2552 (
            .O(N__15299),
            .I(N__15296));
    LocalMux I__2551 (
            .O(N__15296),
            .I(\tok.n4671 ));
    CascadeMux I__2550 (
            .O(N__15293),
            .I(N__15290));
    InMux I__2549 (
            .O(N__15290),
            .I(N__15287));
    LocalMux I__2548 (
            .O(N__15287),
            .I(\tok.n18_adj_672 ));
    InMux I__2547 (
            .O(N__15284),
            .I(N__15281));
    LocalMux I__2546 (
            .O(N__15281),
            .I(N__15278));
    Span4Mux_v I__2545 (
            .O(N__15278),
            .I(N__15275));
    Odrv4 I__2544 (
            .O(N__15275),
            .I(\tok.n6_adj_676 ));
    CascadeMux I__2543 (
            .O(N__15272),
            .I(\tok.n20_adj_674_cascade_ ));
    InMux I__2542 (
            .O(N__15269),
            .I(N__15266));
    LocalMux I__2541 (
            .O(N__15266),
            .I(N__15263));
    Span4Mux_v I__2540 (
            .O(N__15263),
            .I(N__15260));
    Odrv4 I__2539 (
            .O(N__15260),
            .I(\tok.n16_adj_673 ));
    CascadeMux I__2538 (
            .O(N__15257),
            .I(\tok.n4676_cascade_ ));
    InMux I__2537 (
            .O(N__15254),
            .I(N__15251));
    LocalMux I__2536 (
            .O(N__15251),
            .I(\tok.n12_adj_744 ));
    InMux I__2535 (
            .O(N__15248),
            .I(N__15245));
    LocalMux I__2534 (
            .O(N__15245),
            .I(\tok.n4524 ));
    InMux I__2533 (
            .O(N__15242),
            .I(N__15239));
    LocalMux I__2532 (
            .O(N__15239),
            .I(\tok.n12_adj_670 ));
    CascadeMux I__2531 (
            .O(N__15236),
            .I(\tok.n15_cascade_ ));
    CascadeMux I__2530 (
            .O(N__15233),
            .I(N__15230));
    InMux I__2529 (
            .O(N__15230),
            .I(N__15227));
    LocalMux I__2528 (
            .O(N__15227),
            .I(\tok.n183 ));
    CascadeMux I__2527 (
            .O(N__15224),
            .I(N__15221));
    InMux I__2526 (
            .O(N__15221),
            .I(N__15217));
    InMux I__2525 (
            .O(N__15220),
            .I(N__15214));
    LocalMux I__2524 (
            .O(N__15217),
            .I(N__15211));
    LocalMux I__2523 (
            .O(N__15214),
            .I(N__15208));
    Span4Mux_h I__2522 (
            .O(N__15211),
            .I(N__15205));
    Span4Mux_v I__2521 (
            .O(N__15208),
            .I(N__15202));
    Span4Mux_v I__2520 (
            .O(N__15205),
            .I(N__15199));
    Odrv4 I__2519 (
            .O(N__15202),
            .I(\tok.table_rd_6 ));
    Odrv4 I__2518 (
            .O(N__15199),
            .I(\tok.table_rd_6 ));
    CascadeMux I__2517 (
            .O(N__15194),
            .I(\tok.n16_adj_778_cascade_ ));
    InMux I__2516 (
            .O(N__15191),
            .I(N__15188));
    LocalMux I__2515 (
            .O(N__15188),
            .I(N__15185));
    Span4Mux_h I__2514 (
            .O(N__15185),
            .I(N__15182));
    Odrv4 I__2513 (
            .O(N__15182),
            .I(\tok.n6_adj_780 ));
    CascadeMux I__2512 (
            .O(N__15179),
            .I(N__15176));
    InMux I__2511 (
            .O(N__15176),
            .I(N__15173));
    LocalMux I__2510 (
            .O(N__15173),
            .I(N__15170));
    Odrv4 I__2509 (
            .O(N__15170),
            .I(\tok.table_rd_13 ));
    InMux I__2508 (
            .O(N__15167),
            .I(N__15164));
    LocalMux I__2507 (
            .O(N__15164),
            .I(N__15161));
    Span4Mux_h I__2506 (
            .O(N__15161),
            .I(N__15158));
    Odrv4 I__2505 (
            .O(N__15158),
            .I(\tok.table_rd_10 ));
    InMux I__2504 (
            .O(N__15155),
            .I(N__15152));
    LocalMux I__2503 (
            .O(N__15152),
            .I(\tok.n10_adj_671 ));
    CascadeMux I__2502 (
            .O(N__15149),
            .I(\tok.n14_adj_669_cascade_ ));
    InMux I__2501 (
            .O(N__15146),
            .I(N__15143));
    LocalMux I__2500 (
            .O(N__15143),
            .I(N__15140));
    Span4Mux_h I__2499 (
            .O(N__15140),
            .I(N__15137));
    Odrv4 I__2498 (
            .O(N__15137),
            .I(\tok.table_rd_11 ));
    InMux I__2497 (
            .O(N__15134),
            .I(N__15131));
    LocalMux I__2496 (
            .O(N__15131),
            .I(N__15128));
    Span4Mux_h I__2495 (
            .O(N__15128),
            .I(N__15125));
    Odrv4 I__2494 (
            .O(N__15125),
            .I(\tok.n16_adj_691 ));
    InMux I__2493 (
            .O(N__15122),
            .I(N__15118));
    CascadeMux I__2492 (
            .O(N__15121),
            .I(N__15115));
    LocalMux I__2491 (
            .O(N__15118),
            .I(N__15112));
    InMux I__2490 (
            .O(N__15115),
            .I(N__15109));
    Span4Mux_h I__2489 (
            .O(N__15112),
            .I(N__15106));
    LocalMux I__2488 (
            .O(N__15109),
            .I(\tok.key_rd_4 ));
    Odrv4 I__2487 (
            .O(N__15106),
            .I(\tok.key_rd_4 ));
    CascadeMux I__2486 (
            .O(N__15101),
            .I(N__15098));
    InMux I__2485 (
            .O(N__15098),
            .I(N__15095));
    LocalMux I__2484 (
            .O(N__15095),
            .I(N__15091));
    InMux I__2483 (
            .O(N__15094),
            .I(N__15088));
    Span4Mux_h I__2482 (
            .O(N__15091),
            .I(N__15085));
    LocalMux I__2481 (
            .O(N__15088),
            .I(\tok.key_rd_1 ));
    Odrv4 I__2480 (
            .O(N__15085),
            .I(\tok.key_rd_1 ));
    InMux I__2479 (
            .O(N__15080),
            .I(N__15077));
    LocalMux I__2478 (
            .O(N__15077),
            .I(\tok.n18_adj_756 ));
    InMux I__2477 (
            .O(N__15074),
            .I(N__15071));
    LocalMux I__2476 (
            .O(N__15071),
            .I(N__15068));
    Span4Mux_h I__2475 (
            .O(N__15068),
            .I(N__15064));
    InMux I__2474 (
            .O(N__15067),
            .I(N__15061));
    Span4Mux_s3_h I__2473 (
            .O(N__15064),
            .I(N__15058));
    LocalMux I__2472 (
            .O(N__15061),
            .I(\tok.key_rd_0 ));
    Odrv4 I__2471 (
            .O(N__15058),
            .I(\tok.key_rd_0 ));
    CascadeMux I__2470 (
            .O(N__15053),
            .I(N__15050));
    InMux I__2469 (
            .O(N__15050),
            .I(N__15047));
    LocalMux I__2468 (
            .O(N__15047),
            .I(N__15044));
    Span4Mux_v I__2467 (
            .O(N__15044),
            .I(N__15040));
    InMux I__2466 (
            .O(N__15043),
            .I(N__15037));
    Span4Mux_h I__2465 (
            .O(N__15040),
            .I(N__15034));
    LocalMux I__2464 (
            .O(N__15037),
            .I(\tok.key_rd_6 ));
    Odrv4 I__2463 (
            .O(N__15034),
            .I(\tok.key_rd_6 ));
    InMux I__2462 (
            .O(N__15029),
            .I(N__15026));
    LocalMux I__2461 (
            .O(N__15026),
            .I(N__15023));
    Odrv4 I__2460 (
            .O(N__15023),
            .I(\tok.n4645 ));
    InMux I__2459 (
            .O(N__15020),
            .I(N__15017));
    LocalMux I__2458 (
            .O(N__15017),
            .I(N__15014));
    Span4Mux_h I__2457 (
            .O(N__15014),
            .I(N__15011));
    Odrv4 I__2456 (
            .O(N__15011),
            .I(\tok.n13_adj_657 ));
    InMux I__2455 (
            .O(N__15008),
            .I(N__15005));
    LocalMux I__2454 (
            .O(N__15005),
            .I(\tok.n10_adj_656 ));
    InMux I__2453 (
            .O(N__15002),
            .I(N__14999));
    LocalMux I__2452 (
            .O(N__14999),
            .I(N__14996));
    Span4Mux_h I__2451 (
            .O(N__14996),
            .I(N__14993));
    Odrv4 I__2450 (
            .O(N__14993),
            .I(\tok.table_rd_9 ));
    CascadeMux I__2449 (
            .O(N__14990),
            .I(\tok.n30_cascade_ ));
    InMux I__2448 (
            .O(N__14987),
            .I(N__14984));
    LocalMux I__2447 (
            .O(N__14984),
            .I(N__14981));
    Span4Mux_v I__2446 (
            .O(N__14981),
            .I(N__14978));
    Span4Mux_h I__2445 (
            .O(N__14978),
            .I(N__14975));
    Odrv4 I__2444 (
            .O(N__14975),
            .I(\tok.n12_adj_659 ));
    CEMux I__2443 (
            .O(N__14972),
            .I(N__14969));
    LocalMux I__2442 (
            .O(N__14969),
            .I(N__14966));
    Odrv12 I__2441 (
            .O(N__14966),
            .I(\tok.uart.n922 ));
    InMux I__2440 (
            .O(N__14963),
            .I(N__14960));
    LocalMux I__2439 (
            .O(N__14960),
            .I(N__14957));
    Span4Mux_h I__2438 (
            .O(N__14957),
            .I(N__14954));
    Odrv4 I__2437 (
            .O(N__14954),
            .I(\tok.n301 ));
    CascadeMux I__2436 (
            .O(N__14951),
            .I(\tok.n19_adj_860_cascade_ ));
    InMux I__2435 (
            .O(N__14948),
            .I(N__14945));
    LocalMux I__2434 (
            .O(N__14945),
            .I(\tok.n17_adj_861 ));
    InMux I__2433 (
            .O(N__14942),
            .I(N__14939));
    LocalMux I__2432 (
            .O(N__14939),
            .I(\tok.n29_adj_864 ));
    InMux I__2431 (
            .O(N__14936),
            .I(N__14933));
    LocalMux I__2430 (
            .O(N__14933),
            .I(N__14930));
    Span4Mux_h I__2429 (
            .O(N__14930),
            .I(N__14926));
    InMux I__2428 (
            .O(N__14929),
            .I(N__14923));
    Span4Mux_v I__2427 (
            .O(N__14926),
            .I(N__14918));
    LocalMux I__2426 (
            .O(N__14923),
            .I(N__14918));
    Span4Mux_h I__2425 (
            .O(N__14918),
            .I(N__14915));
    Span4Mux_s2_h I__2424 (
            .O(N__14915),
            .I(N__14911));
    InMux I__2423 (
            .O(N__14914),
            .I(N__14908));
    Odrv4 I__2422 (
            .O(N__14911),
            .I(capture_8));
    LocalMux I__2421 (
            .O(N__14908),
            .I(capture_8));
    CascadeMux I__2420 (
            .O(N__14903),
            .I(N__14900));
    InMux I__2419 (
            .O(N__14900),
            .I(N__14896));
    InMux I__2418 (
            .O(N__14899),
            .I(N__14893));
    LocalMux I__2417 (
            .O(N__14896),
            .I(uart_rx_data_7));
    LocalMux I__2416 (
            .O(N__14893),
            .I(uart_rx_data_7));
    InMux I__2415 (
            .O(N__14888),
            .I(N__14885));
    LocalMux I__2414 (
            .O(N__14885),
            .I(N__14882));
    Span4Mux_v I__2413 (
            .O(N__14882),
            .I(N__14879));
    Span4Mux_h I__2412 (
            .O(N__14879),
            .I(N__14876));
    Odrv4 I__2411 (
            .O(N__14876),
            .I(\tok.table_wr_data_10 ));
    CascadeMux I__2410 (
            .O(N__14873),
            .I(N__14870));
    InMux I__2409 (
            .O(N__14870),
            .I(N__14867));
    LocalMux I__2408 (
            .O(N__14867),
            .I(N__14864));
    Span4Mux_h I__2407 (
            .O(N__14864),
            .I(N__14861));
    Span4Mux_v I__2406 (
            .O(N__14861),
            .I(N__14858));
    Odrv4 I__2405 (
            .O(N__14858),
            .I(\tok.n293 ));
    InMux I__2404 (
            .O(N__14855),
            .I(N__14852));
    LocalMux I__2403 (
            .O(N__14852),
            .I(N__14849));
    Odrv4 I__2402 (
            .O(N__14849),
            .I(\tok.n2634 ));
    SRMux I__2401 (
            .O(N__14846),
            .I(N__14842));
    SRMux I__2400 (
            .O(N__14845),
            .I(N__14839));
    LocalMux I__2399 (
            .O(N__14842),
            .I(N__14834));
    LocalMux I__2398 (
            .O(N__14839),
            .I(N__14834));
    Span4Mux_v I__2397 (
            .O(N__14834),
            .I(N__14831));
    Span4Mux_s3_h I__2396 (
            .O(N__14831),
            .I(N__14828));
    Span4Mux_h I__2395 (
            .O(N__14828),
            .I(N__14825));
    Odrv4 I__2394 (
            .O(N__14825),
            .I(\tok.write_slot ));
    InMux I__2393 (
            .O(N__14822),
            .I(N__14819));
    LocalMux I__2392 (
            .O(N__14819),
            .I(N__14816));
    Span4Mux_h I__2391 (
            .O(N__14816),
            .I(N__14813));
    Span4Mux_s3_h I__2390 (
            .O(N__14813),
            .I(N__14810));
    Span4Mux_h I__2389 (
            .O(N__14810),
            .I(N__14807));
    Odrv4 I__2388 (
            .O(N__14807),
            .I(\tok.table_wr_data_5 ));
    CascadeMux I__2387 (
            .O(N__14804),
            .I(\tok.n83_adj_716_cascade_ ));
    CascadeMux I__2386 (
            .O(N__14801),
            .I(\tok.n12_adj_740_cascade_ ));
    CascadeMux I__2385 (
            .O(N__14798),
            .I(\tok.n12_adj_801_cascade_ ));
    InMux I__2384 (
            .O(N__14795),
            .I(N__14792));
    LocalMux I__2383 (
            .O(N__14792),
            .I(\tok.n284 ));
    CascadeMux I__2382 (
            .O(N__14789),
            .I(\tok.n284_cascade_ ));
    CascadeMux I__2381 (
            .O(N__14786),
            .I(\tok.n182_cascade_ ));
    InMux I__2380 (
            .O(N__14783),
            .I(N__14780));
    LocalMux I__2379 (
            .O(N__14780),
            .I(N__14777));
    Span4Mux_h I__2378 (
            .O(N__14777),
            .I(N__14774));
    Odrv4 I__2377 (
            .O(N__14774),
            .I(\tok.n12_adj_766 ));
    CascadeMux I__2376 (
            .O(N__14771),
            .I(N__14768));
    InMux I__2375 (
            .O(N__14768),
            .I(N__14765));
    LocalMux I__2374 (
            .O(N__14765),
            .I(N__14762));
    Span4Mux_h I__2373 (
            .O(N__14762),
            .I(N__14759));
    Odrv4 I__2372 (
            .O(N__14759),
            .I(\tok.n24_adj_854 ));
    InMux I__2371 (
            .O(N__14756),
            .I(N__14753));
    LocalMux I__2370 (
            .O(N__14753),
            .I(N__14750));
    Span12Mux_s9_h I__2369 (
            .O(N__14750),
            .I(N__14747));
    Odrv12 I__2368 (
            .O(N__14747),
            .I(\tok.n21_adj_857 ));
    CascadeMux I__2367 (
            .O(N__14744),
            .I(\tok.n30_adj_862_cascade_ ));
    CascadeMux I__2366 (
            .O(N__14741),
            .I(n29_cascade_));
    CEMux I__2365 (
            .O(N__14738),
            .I(N__14733));
    CEMux I__2364 (
            .O(N__14737),
            .I(N__14730));
    CEMux I__2363 (
            .O(N__14736),
            .I(N__14723));
    LocalMux I__2362 (
            .O(N__14733),
            .I(N__14717));
    LocalMux I__2361 (
            .O(N__14730),
            .I(N__14717));
    CEMux I__2360 (
            .O(N__14729),
            .I(N__14714));
    CEMux I__2359 (
            .O(N__14728),
            .I(N__14709));
    CEMux I__2358 (
            .O(N__14727),
            .I(N__14704));
    CEMux I__2357 (
            .O(N__14726),
            .I(N__14700));
    LocalMux I__2356 (
            .O(N__14723),
            .I(N__14697));
    CEMux I__2355 (
            .O(N__14722),
            .I(N__14694));
    Span4Mux_v I__2354 (
            .O(N__14717),
            .I(N__14689));
    LocalMux I__2353 (
            .O(N__14714),
            .I(N__14689));
    CEMux I__2352 (
            .O(N__14713),
            .I(N__14686));
    CEMux I__2351 (
            .O(N__14712),
            .I(N__14683));
    LocalMux I__2350 (
            .O(N__14709),
            .I(N__14677));
    CEMux I__2349 (
            .O(N__14708),
            .I(N__14674));
    CEMux I__2348 (
            .O(N__14707),
            .I(N__14671));
    LocalMux I__2347 (
            .O(N__14704),
            .I(N__14668));
    CEMux I__2346 (
            .O(N__14703),
            .I(N__14665));
    LocalMux I__2345 (
            .O(N__14700),
            .I(N__14661));
    Span4Mux_s3_h I__2344 (
            .O(N__14697),
            .I(N__14656));
    LocalMux I__2343 (
            .O(N__14694),
            .I(N__14656));
    Span4Mux_s2_h I__2342 (
            .O(N__14689),
            .I(N__14651));
    LocalMux I__2341 (
            .O(N__14686),
            .I(N__14651));
    LocalMux I__2340 (
            .O(N__14683),
            .I(N__14648));
    CEMux I__2339 (
            .O(N__14682),
            .I(N__14645));
    CEMux I__2338 (
            .O(N__14681),
            .I(N__14642));
    CEMux I__2337 (
            .O(N__14680),
            .I(N__14639));
    Span4Mux_h I__2336 (
            .O(N__14677),
            .I(N__14634));
    LocalMux I__2335 (
            .O(N__14674),
            .I(N__14634));
    LocalMux I__2334 (
            .O(N__14671),
            .I(N__14631));
    Span4Mux_v I__2333 (
            .O(N__14668),
            .I(N__14626));
    LocalMux I__2332 (
            .O(N__14665),
            .I(N__14626));
    CEMux I__2331 (
            .O(N__14664),
            .I(N__14623));
    Span4Mux_h I__2330 (
            .O(N__14661),
            .I(N__14620));
    Span4Mux_h I__2329 (
            .O(N__14656),
            .I(N__14617));
    Span4Mux_h I__2328 (
            .O(N__14651),
            .I(N__14606));
    Span4Mux_v I__2327 (
            .O(N__14648),
            .I(N__14606));
    LocalMux I__2326 (
            .O(N__14645),
            .I(N__14606));
    LocalMux I__2325 (
            .O(N__14642),
            .I(N__14606));
    LocalMux I__2324 (
            .O(N__14639),
            .I(N__14606));
    Span4Mux_v I__2323 (
            .O(N__14634),
            .I(N__14597));
    Span4Mux_h I__2322 (
            .O(N__14631),
            .I(N__14597));
    Span4Mux_s2_v I__2321 (
            .O(N__14626),
            .I(N__14597));
    LocalMux I__2320 (
            .O(N__14623),
            .I(N__14597));
    Odrv4 I__2319 (
            .O(N__14620),
            .I(\tok.A_stk.rd_15__N_301 ));
    Odrv4 I__2318 (
            .O(N__14617),
            .I(\tok.A_stk.rd_15__N_301 ));
    Odrv4 I__2317 (
            .O(N__14606),
            .I(\tok.A_stk.rd_15__N_301 ));
    Odrv4 I__2316 (
            .O(N__14597),
            .I(\tok.A_stk.rd_15__N_301 ));
    CascadeMux I__2315 (
            .O(N__14588),
            .I(\tok.n83_adj_735_cascade_ ));
    CascadeMux I__2314 (
            .O(N__14585),
            .I(\tok.n7_cascade_ ));
    InMux I__2313 (
            .O(N__14582),
            .I(N__14579));
    LocalMux I__2312 (
            .O(N__14579),
            .I(\tok.n4516 ));
    InMux I__2311 (
            .O(N__14576),
            .I(N__14573));
    LocalMux I__2310 (
            .O(N__14573),
            .I(N__14569));
    InMux I__2309 (
            .O(N__14572),
            .I(N__14566));
    Span12Mux_s6_h I__2308 (
            .O(N__14569),
            .I(N__14563));
    LocalMux I__2307 (
            .O(N__14566),
            .I(capture_0));
    Odrv12 I__2306 (
            .O(N__14563),
            .I(capture_0));
    InMux I__2305 (
            .O(N__14558),
            .I(N__14554));
    InMux I__2304 (
            .O(N__14557),
            .I(N__14551));
    LocalMux I__2303 (
            .O(N__14554),
            .I(\tok.n17 ));
    LocalMux I__2302 (
            .O(N__14551),
            .I(\tok.n17 ));
    CascadeMux I__2301 (
            .O(N__14546),
            .I(\tok.n4_adj_654_cascade_ ));
    InMux I__2300 (
            .O(N__14543),
            .I(N__14491));
    InMux I__2299 (
            .O(N__14542),
            .I(N__14491));
    InMux I__2298 (
            .O(N__14541),
            .I(N__14491));
    InMux I__2297 (
            .O(N__14540),
            .I(N__14491));
    InMux I__2296 (
            .O(N__14539),
            .I(N__14491));
    InMux I__2295 (
            .O(N__14538),
            .I(N__14491));
    InMux I__2294 (
            .O(N__14537),
            .I(N__14491));
    InMux I__2293 (
            .O(N__14536),
            .I(N__14469));
    InMux I__2292 (
            .O(N__14535),
            .I(N__14469));
    InMux I__2291 (
            .O(N__14534),
            .I(N__14469));
    InMux I__2290 (
            .O(N__14533),
            .I(N__14469));
    InMux I__2289 (
            .O(N__14532),
            .I(N__14469));
    InMux I__2288 (
            .O(N__14531),
            .I(N__14469));
    InMux I__2287 (
            .O(N__14530),
            .I(N__14469));
    CascadeMux I__2286 (
            .O(N__14529),
            .I(N__14451));
    CascadeMux I__2285 (
            .O(N__14528),
            .I(N__14448));
    InMux I__2284 (
            .O(N__14527),
            .I(N__14431));
    InMux I__2283 (
            .O(N__14526),
            .I(N__14431));
    InMux I__2282 (
            .O(N__14525),
            .I(N__14431));
    InMux I__2281 (
            .O(N__14524),
            .I(N__14431));
    InMux I__2280 (
            .O(N__14523),
            .I(N__14431));
    InMux I__2279 (
            .O(N__14522),
            .I(N__14431));
    InMux I__2278 (
            .O(N__14521),
            .I(N__14388));
    InMux I__2277 (
            .O(N__14520),
            .I(N__14388));
    InMux I__2276 (
            .O(N__14519),
            .I(N__14388));
    InMux I__2275 (
            .O(N__14518),
            .I(N__14388));
    InMux I__2274 (
            .O(N__14517),
            .I(N__14388));
    InMux I__2273 (
            .O(N__14516),
            .I(N__14388));
    InMux I__2272 (
            .O(N__14515),
            .I(N__14388));
    InMux I__2271 (
            .O(N__14514),
            .I(N__14378));
    InMux I__2270 (
            .O(N__14513),
            .I(N__14375));
    InMux I__2269 (
            .O(N__14512),
            .I(N__14360));
    InMux I__2268 (
            .O(N__14511),
            .I(N__14360));
    InMux I__2267 (
            .O(N__14510),
            .I(N__14360));
    InMux I__2266 (
            .O(N__14509),
            .I(N__14360));
    InMux I__2265 (
            .O(N__14508),
            .I(N__14360));
    InMux I__2264 (
            .O(N__14507),
            .I(N__14360));
    InMux I__2263 (
            .O(N__14506),
            .I(N__14360));
    LocalMux I__2262 (
            .O(N__14491),
            .I(N__14357));
    InMux I__2261 (
            .O(N__14490),
            .I(N__14342));
    InMux I__2260 (
            .O(N__14489),
            .I(N__14342));
    InMux I__2259 (
            .O(N__14488),
            .I(N__14342));
    InMux I__2258 (
            .O(N__14487),
            .I(N__14342));
    InMux I__2257 (
            .O(N__14486),
            .I(N__14342));
    InMux I__2256 (
            .O(N__14485),
            .I(N__14342));
    InMux I__2255 (
            .O(N__14484),
            .I(N__14342));
    LocalMux I__2254 (
            .O(N__14469),
            .I(N__14339));
    InMux I__2253 (
            .O(N__14468),
            .I(N__14330));
    InMux I__2252 (
            .O(N__14467),
            .I(N__14315));
    InMux I__2251 (
            .O(N__14466),
            .I(N__14315));
    InMux I__2250 (
            .O(N__14465),
            .I(N__14315));
    InMux I__2249 (
            .O(N__14464),
            .I(N__14315));
    InMux I__2248 (
            .O(N__14463),
            .I(N__14315));
    InMux I__2247 (
            .O(N__14462),
            .I(N__14315));
    InMux I__2246 (
            .O(N__14461),
            .I(N__14315));
    InMux I__2245 (
            .O(N__14460),
            .I(N__14300));
    InMux I__2244 (
            .O(N__14459),
            .I(N__14300));
    InMux I__2243 (
            .O(N__14458),
            .I(N__14300));
    InMux I__2242 (
            .O(N__14457),
            .I(N__14300));
    InMux I__2241 (
            .O(N__14456),
            .I(N__14300));
    InMux I__2240 (
            .O(N__14455),
            .I(N__14300));
    InMux I__2239 (
            .O(N__14454),
            .I(N__14300));
    InMux I__2238 (
            .O(N__14451),
            .I(N__14295));
    InMux I__2237 (
            .O(N__14448),
            .I(N__14295));
    InMux I__2236 (
            .O(N__14447),
            .I(N__14286));
    InMux I__2235 (
            .O(N__14446),
            .I(N__14286));
    InMux I__2234 (
            .O(N__14445),
            .I(N__14286));
    InMux I__2233 (
            .O(N__14444),
            .I(N__14286));
    LocalMux I__2232 (
            .O(N__14431),
            .I(N__14283));
    InMux I__2231 (
            .O(N__14430),
            .I(N__14268));
    InMux I__2230 (
            .O(N__14429),
            .I(N__14268));
    InMux I__2229 (
            .O(N__14428),
            .I(N__14268));
    InMux I__2228 (
            .O(N__14427),
            .I(N__14268));
    InMux I__2227 (
            .O(N__14426),
            .I(N__14268));
    InMux I__2226 (
            .O(N__14425),
            .I(N__14268));
    InMux I__2225 (
            .O(N__14424),
            .I(N__14268));
    InMux I__2224 (
            .O(N__14423),
            .I(N__14253));
    InMux I__2223 (
            .O(N__14422),
            .I(N__14253));
    InMux I__2222 (
            .O(N__14421),
            .I(N__14253));
    InMux I__2221 (
            .O(N__14420),
            .I(N__14253));
    InMux I__2220 (
            .O(N__14419),
            .I(N__14253));
    InMux I__2219 (
            .O(N__14418),
            .I(N__14253));
    InMux I__2218 (
            .O(N__14417),
            .I(N__14253));
    InMux I__2217 (
            .O(N__14416),
            .I(N__14217));
    InMux I__2216 (
            .O(N__14415),
            .I(N__14217));
    InMux I__2215 (
            .O(N__14414),
            .I(N__14217));
    InMux I__2214 (
            .O(N__14413),
            .I(N__14217));
    InMux I__2213 (
            .O(N__14412),
            .I(N__14217));
    InMux I__2212 (
            .O(N__14411),
            .I(N__14217));
    InMux I__2211 (
            .O(N__14410),
            .I(N__14217));
    InMux I__2210 (
            .O(N__14409),
            .I(N__14202));
    InMux I__2209 (
            .O(N__14408),
            .I(N__14202));
    InMux I__2208 (
            .O(N__14407),
            .I(N__14202));
    InMux I__2207 (
            .O(N__14406),
            .I(N__14202));
    InMux I__2206 (
            .O(N__14405),
            .I(N__14202));
    InMux I__2205 (
            .O(N__14404),
            .I(N__14202));
    InMux I__2204 (
            .O(N__14403),
            .I(N__14202));
    LocalMux I__2203 (
            .O(N__14388),
            .I(N__14199));
    InMux I__2202 (
            .O(N__14387),
            .I(N__14184));
    InMux I__2201 (
            .O(N__14386),
            .I(N__14184));
    InMux I__2200 (
            .O(N__14385),
            .I(N__14184));
    InMux I__2199 (
            .O(N__14384),
            .I(N__14184));
    InMux I__2198 (
            .O(N__14383),
            .I(N__14184));
    InMux I__2197 (
            .O(N__14382),
            .I(N__14184));
    InMux I__2196 (
            .O(N__14381),
            .I(N__14184));
    LocalMux I__2195 (
            .O(N__14378),
            .I(N__14179));
    LocalMux I__2194 (
            .O(N__14375),
            .I(N__14179));
    LocalMux I__2193 (
            .O(N__14360),
            .I(N__14174));
    Span4Mux_s2_h I__2192 (
            .O(N__14357),
            .I(N__14174));
    LocalMux I__2191 (
            .O(N__14342),
            .I(N__14171));
    Span4Mux_s2_h I__2190 (
            .O(N__14339),
            .I(N__14168));
    InMux I__2189 (
            .O(N__14338),
            .I(N__14155));
    InMux I__2188 (
            .O(N__14337),
            .I(N__14155));
    InMux I__2187 (
            .O(N__14336),
            .I(N__14155));
    InMux I__2186 (
            .O(N__14335),
            .I(N__14155));
    InMux I__2185 (
            .O(N__14334),
            .I(N__14155));
    InMux I__2184 (
            .O(N__14333),
            .I(N__14155));
    LocalMux I__2183 (
            .O(N__14330),
            .I(N__14148));
    LocalMux I__2182 (
            .O(N__14315),
            .I(N__14148));
    LocalMux I__2181 (
            .O(N__14300),
            .I(N__14148));
    LocalMux I__2180 (
            .O(N__14295),
            .I(N__14137));
    LocalMux I__2179 (
            .O(N__14286),
            .I(N__14137));
    Span4Mux_s3_v I__2178 (
            .O(N__14283),
            .I(N__14137));
    LocalMux I__2177 (
            .O(N__14268),
            .I(N__14137));
    LocalMux I__2176 (
            .O(N__14253),
            .I(N__14137));
    InMux I__2175 (
            .O(N__14252),
            .I(N__14119));
    InMux I__2174 (
            .O(N__14251),
            .I(N__14119));
    InMux I__2173 (
            .O(N__14250),
            .I(N__14119));
    InMux I__2172 (
            .O(N__14249),
            .I(N__14119));
    InMux I__2171 (
            .O(N__14248),
            .I(N__14119));
    InMux I__2170 (
            .O(N__14247),
            .I(N__14119));
    InMux I__2169 (
            .O(N__14246),
            .I(N__14119));
    InMux I__2168 (
            .O(N__14245),
            .I(N__14104));
    InMux I__2167 (
            .O(N__14244),
            .I(N__14104));
    InMux I__2166 (
            .O(N__14243),
            .I(N__14104));
    InMux I__2165 (
            .O(N__14242),
            .I(N__14104));
    InMux I__2164 (
            .O(N__14241),
            .I(N__14104));
    InMux I__2163 (
            .O(N__14240),
            .I(N__14104));
    InMux I__2162 (
            .O(N__14239),
            .I(N__14104));
    InMux I__2161 (
            .O(N__14238),
            .I(N__14089));
    InMux I__2160 (
            .O(N__14237),
            .I(N__14089));
    InMux I__2159 (
            .O(N__14236),
            .I(N__14089));
    InMux I__2158 (
            .O(N__14235),
            .I(N__14089));
    InMux I__2157 (
            .O(N__14234),
            .I(N__14089));
    InMux I__2156 (
            .O(N__14233),
            .I(N__14089));
    InMux I__2155 (
            .O(N__14232),
            .I(N__14089));
    LocalMux I__2154 (
            .O(N__14217),
            .I(N__14082));
    LocalMux I__2153 (
            .O(N__14202),
            .I(N__14082));
    Span4Mux_h I__2152 (
            .O(N__14199),
            .I(N__14082));
    LocalMux I__2151 (
            .O(N__14184),
            .I(N__14075));
    Span4Mux_h I__2150 (
            .O(N__14179),
            .I(N__14075));
    Span4Mux_h I__2149 (
            .O(N__14174),
            .I(N__14075));
    Span4Mux_h I__2148 (
            .O(N__14171),
            .I(N__14070));
    Span4Mux_h I__2147 (
            .O(N__14168),
            .I(N__14070));
    LocalMux I__2146 (
            .O(N__14155),
            .I(N__14063));
    Span4Mux_s3_h I__2145 (
            .O(N__14148),
            .I(N__14063));
    Span4Mux_v I__2144 (
            .O(N__14137),
            .I(N__14063));
    InMux I__2143 (
            .O(N__14136),
            .I(N__14056));
    InMux I__2142 (
            .O(N__14135),
            .I(N__14056));
    InMux I__2141 (
            .O(N__14134),
            .I(N__14056));
    LocalMux I__2140 (
            .O(N__14119),
            .I(n786));
    LocalMux I__2139 (
            .O(N__14104),
            .I(n786));
    LocalMux I__2138 (
            .O(N__14089),
            .I(n786));
    Odrv4 I__2137 (
            .O(N__14082),
            .I(n786));
    Odrv4 I__2136 (
            .O(N__14075),
            .I(n786));
    Odrv4 I__2135 (
            .O(N__14070),
            .I(n786));
    Odrv4 I__2134 (
            .O(N__14063),
            .I(n786));
    LocalMux I__2133 (
            .O(N__14056),
            .I(n786));
    CascadeMux I__2132 (
            .O(N__14039),
            .I(N__14035));
    InMux I__2131 (
            .O(N__14038),
            .I(N__14030));
    InMux I__2130 (
            .O(N__14035),
            .I(N__14030));
    LocalMux I__2129 (
            .O(N__14030),
            .I(\tok.A_stk.tail_31 ));
    InMux I__2128 (
            .O(N__14027),
            .I(N__14021));
    InMux I__2127 (
            .O(N__14026),
            .I(N__14021));
    LocalMux I__2126 (
            .O(N__14021),
            .I(\tok.A_stk.tail_15 ));
    InMux I__2125 (
            .O(N__14018),
            .I(N__14012));
    InMux I__2124 (
            .O(N__14017),
            .I(N__14012));
    LocalMux I__2123 (
            .O(N__14012),
            .I(\tok.A_stk.tail_79 ));
    CascadeMux I__2122 (
            .O(N__14009),
            .I(N__14006));
    InMux I__2121 (
            .O(N__14006),
            .I(N__14000));
    InMux I__2120 (
            .O(N__14005),
            .I(N__14000));
    LocalMux I__2119 (
            .O(N__14000),
            .I(\tok.A_stk.tail_95 ));
    InMux I__2118 (
            .O(N__13997),
            .I(N__13993));
    InMux I__2117 (
            .O(N__13996),
            .I(N__13990));
    LocalMux I__2116 (
            .O(N__13993),
            .I(tail_111));
    LocalMux I__2115 (
            .O(N__13990),
            .I(tail_111));
    CascadeMux I__2114 (
            .O(N__13985),
            .I(N__13982));
    InMux I__2113 (
            .O(N__13982),
            .I(N__13978));
    InMux I__2112 (
            .O(N__13981),
            .I(N__13975));
    LocalMux I__2111 (
            .O(N__13978),
            .I(N__13972));
    LocalMux I__2110 (
            .O(N__13975),
            .I(N__13969));
    Odrv4 I__2109 (
            .O(N__13972),
            .I(tail_127));
    Odrv4 I__2108 (
            .O(N__13969),
            .I(tail_127));
    CascadeMux I__2107 (
            .O(N__13964),
            .I(N__13961));
    InMux I__2106 (
            .O(N__13961),
            .I(N__13957));
    InMux I__2105 (
            .O(N__13960),
            .I(N__13954));
    LocalMux I__2104 (
            .O(N__13957),
            .I(tail_97));
    LocalMux I__2103 (
            .O(N__13954),
            .I(tail_97));
    CascadeMux I__2102 (
            .O(N__13949),
            .I(N__13946));
    InMux I__2101 (
            .O(N__13946),
            .I(N__13942));
    InMux I__2100 (
            .O(N__13945),
            .I(N__13939));
    LocalMux I__2099 (
            .O(N__13942),
            .I(tail_113));
    LocalMux I__2098 (
            .O(N__13939),
            .I(tail_113));
    CascadeMux I__2097 (
            .O(N__13934),
            .I(N__13918));
    CascadeMux I__2096 (
            .O(N__13933),
            .I(N__13915));
    CascadeMux I__2095 (
            .O(N__13932),
            .I(N__13912));
    CascadeMux I__2094 (
            .O(N__13931),
            .I(N__13901));
    CascadeMux I__2093 (
            .O(N__13930),
            .I(N__13898));
    CascadeMux I__2092 (
            .O(N__13929),
            .I(N__13895));
    CascadeMux I__2091 (
            .O(N__13928),
            .I(N__13867));
    CascadeMux I__2090 (
            .O(N__13927),
            .I(N__13864));
    CascadeMux I__2089 (
            .O(N__13926),
            .I(N__13861));
    CascadeMux I__2088 (
            .O(N__13925),
            .I(N__13854));
    CascadeMux I__2087 (
            .O(N__13924),
            .I(N__13851));
    CascadeMux I__2086 (
            .O(N__13923),
            .I(N__13848));
    CascadeMux I__2085 (
            .O(N__13922),
            .I(N__13843));
    InMux I__2084 (
            .O(N__13921),
            .I(N__13821));
    InMux I__2083 (
            .O(N__13918),
            .I(N__13821));
    InMux I__2082 (
            .O(N__13915),
            .I(N__13821));
    InMux I__2081 (
            .O(N__13912),
            .I(N__13821));
    InMux I__2080 (
            .O(N__13911),
            .I(N__13821));
    InMux I__2079 (
            .O(N__13910),
            .I(N__13821));
    InMux I__2078 (
            .O(N__13909),
            .I(N__13821));
    InMux I__2077 (
            .O(N__13908),
            .I(N__13818));
    CascadeMux I__2076 (
            .O(N__13907),
            .I(N__13810));
    CascadeMux I__2075 (
            .O(N__13906),
            .I(N__13807));
    CascadeMux I__2074 (
            .O(N__13905),
            .I(N__13804));
    InMux I__2073 (
            .O(N__13904),
            .I(N__13785));
    InMux I__2072 (
            .O(N__13901),
            .I(N__13785));
    InMux I__2071 (
            .O(N__13898),
            .I(N__13785));
    InMux I__2070 (
            .O(N__13895),
            .I(N__13785));
    InMux I__2069 (
            .O(N__13894),
            .I(N__13785));
    InMux I__2068 (
            .O(N__13893),
            .I(N__13785));
    InMux I__2067 (
            .O(N__13892),
            .I(N__13785));
    InMux I__2066 (
            .O(N__13891),
            .I(N__13772));
    InMux I__2065 (
            .O(N__13890),
            .I(N__13772));
    InMux I__2064 (
            .O(N__13889),
            .I(N__13772));
    CascadeMux I__2063 (
            .O(N__13888),
            .I(N__13764));
    CascadeMux I__2062 (
            .O(N__13887),
            .I(N__13761));
    CascadeMux I__2061 (
            .O(N__13886),
            .I(N__13758));
    CascadeMux I__2060 (
            .O(N__13885),
            .I(N__13752));
    CascadeMux I__2059 (
            .O(N__13884),
            .I(N__13749));
    InMux I__2058 (
            .O(N__13883),
            .I(N__13730));
    InMux I__2057 (
            .O(N__13882),
            .I(N__13730));
    InMux I__2056 (
            .O(N__13881),
            .I(N__13730));
    InMux I__2055 (
            .O(N__13880),
            .I(N__13730));
    InMux I__2054 (
            .O(N__13879),
            .I(N__13730));
    InMux I__2053 (
            .O(N__13878),
            .I(N__13730));
    InMux I__2052 (
            .O(N__13877),
            .I(N__13730));
    CascadeMux I__2051 (
            .O(N__13876),
            .I(N__13716));
    CascadeMux I__2050 (
            .O(N__13875),
            .I(N__13712));
    CascadeMux I__2049 (
            .O(N__13874),
            .I(N__13709));
    CascadeMux I__2048 (
            .O(N__13873),
            .I(N__13706));
    InMux I__2047 (
            .O(N__13872),
            .I(N__13696));
    InMux I__2046 (
            .O(N__13871),
            .I(N__13696));
    InMux I__2045 (
            .O(N__13870),
            .I(N__13696));
    InMux I__2044 (
            .O(N__13867),
            .I(N__13683));
    InMux I__2043 (
            .O(N__13864),
            .I(N__13683));
    InMux I__2042 (
            .O(N__13861),
            .I(N__13683));
    InMux I__2041 (
            .O(N__13860),
            .I(N__13683));
    InMux I__2040 (
            .O(N__13859),
            .I(N__13683));
    InMux I__2039 (
            .O(N__13858),
            .I(N__13683));
    InMux I__2038 (
            .O(N__13857),
            .I(N__13670));
    InMux I__2037 (
            .O(N__13854),
            .I(N__13670));
    InMux I__2036 (
            .O(N__13851),
            .I(N__13670));
    InMux I__2035 (
            .O(N__13848),
            .I(N__13670));
    InMux I__2034 (
            .O(N__13847),
            .I(N__13670));
    InMux I__2033 (
            .O(N__13846),
            .I(N__13670));
    InMux I__2032 (
            .O(N__13843),
            .I(N__13667));
    InMux I__2031 (
            .O(N__13842),
            .I(N__13660));
    InMux I__2030 (
            .O(N__13841),
            .I(N__13660));
    InMux I__2029 (
            .O(N__13840),
            .I(N__13660));
    InMux I__2028 (
            .O(N__13839),
            .I(N__13651));
    InMux I__2027 (
            .O(N__13838),
            .I(N__13651));
    InMux I__2026 (
            .O(N__13837),
            .I(N__13651));
    InMux I__2025 (
            .O(N__13836),
            .I(N__13651));
    LocalMux I__2024 (
            .O(N__13821),
            .I(N__13646));
    LocalMux I__2023 (
            .O(N__13818),
            .I(N__13646));
    InMux I__2022 (
            .O(N__13817),
            .I(N__13635));
    InMux I__2021 (
            .O(N__13816),
            .I(N__13632));
    InMux I__2020 (
            .O(N__13815),
            .I(N__13619));
    InMux I__2019 (
            .O(N__13814),
            .I(N__13619));
    InMux I__2018 (
            .O(N__13813),
            .I(N__13619));
    InMux I__2017 (
            .O(N__13810),
            .I(N__13619));
    InMux I__2016 (
            .O(N__13807),
            .I(N__13619));
    InMux I__2015 (
            .O(N__13804),
            .I(N__13619));
    InMux I__2014 (
            .O(N__13803),
            .I(N__13610));
    InMux I__2013 (
            .O(N__13802),
            .I(N__13610));
    InMux I__2012 (
            .O(N__13801),
            .I(N__13610));
    InMux I__2011 (
            .O(N__13800),
            .I(N__13610));
    LocalMux I__2010 (
            .O(N__13785),
            .I(N__13607));
    InMux I__2009 (
            .O(N__13784),
            .I(N__13594));
    InMux I__2008 (
            .O(N__13783),
            .I(N__13594));
    InMux I__2007 (
            .O(N__13782),
            .I(N__13594));
    InMux I__2006 (
            .O(N__13781),
            .I(N__13594));
    InMux I__2005 (
            .O(N__13780),
            .I(N__13594));
    InMux I__2004 (
            .O(N__13779),
            .I(N__13594));
    LocalMux I__2003 (
            .O(N__13772),
            .I(N__13591));
    InMux I__2002 (
            .O(N__13771),
            .I(N__13582));
    InMux I__2001 (
            .O(N__13770),
            .I(N__13582));
    InMux I__2000 (
            .O(N__13769),
            .I(N__13582));
    InMux I__1999 (
            .O(N__13768),
            .I(N__13582));
    InMux I__1998 (
            .O(N__13767),
            .I(N__13567));
    InMux I__1997 (
            .O(N__13764),
            .I(N__13567));
    InMux I__1996 (
            .O(N__13761),
            .I(N__13567));
    InMux I__1995 (
            .O(N__13758),
            .I(N__13567));
    InMux I__1994 (
            .O(N__13757),
            .I(N__13567));
    InMux I__1993 (
            .O(N__13756),
            .I(N__13567));
    InMux I__1992 (
            .O(N__13755),
            .I(N__13567));
    InMux I__1991 (
            .O(N__13752),
            .I(N__13554));
    InMux I__1990 (
            .O(N__13749),
            .I(N__13554));
    InMux I__1989 (
            .O(N__13748),
            .I(N__13554));
    InMux I__1988 (
            .O(N__13747),
            .I(N__13554));
    InMux I__1987 (
            .O(N__13746),
            .I(N__13554));
    InMux I__1986 (
            .O(N__13745),
            .I(N__13554));
    LocalMux I__1985 (
            .O(N__13730),
            .I(N__13551));
    CascadeMux I__1984 (
            .O(N__13729),
            .I(N__13548));
    CascadeMux I__1983 (
            .O(N__13728),
            .I(N__13545));
    CascadeMux I__1982 (
            .O(N__13727),
            .I(N__13542));
    CascadeMux I__1981 (
            .O(N__13726),
            .I(N__13539));
    CascadeMux I__1980 (
            .O(N__13725),
            .I(N__13533));
    CascadeMux I__1979 (
            .O(N__13724),
            .I(N__13530));
    CascadeMux I__1978 (
            .O(N__13723),
            .I(N__13527));
    CascadeMux I__1977 (
            .O(N__13722),
            .I(N__13520));
    CascadeMux I__1976 (
            .O(N__13721),
            .I(N__13517));
    CascadeMux I__1975 (
            .O(N__13720),
            .I(N__13514));
    CascadeMux I__1974 (
            .O(N__13719),
            .I(N__13508));
    InMux I__1973 (
            .O(N__13716),
            .I(N__13497));
    InMux I__1972 (
            .O(N__13715),
            .I(N__13482));
    InMux I__1971 (
            .O(N__13712),
            .I(N__13482));
    InMux I__1970 (
            .O(N__13709),
            .I(N__13482));
    InMux I__1969 (
            .O(N__13706),
            .I(N__13482));
    InMux I__1968 (
            .O(N__13705),
            .I(N__13482));
    InMux I__1967 (
            .O(N__13704),
            .I(N__13482));
    InMux I__1966 (
            .O(N__13703),
            .I(N__13482));
    LocalMux I__1965 (
            .O(N__13696),
            .I(N__13473));
    LocalMux I__1964 (
            .O(N__13683),
            .I(N__13473));
    LocalMux I__1963 (
            .O(N__13670),
            .I(N__13473));
    LocalMux I__1962 (
            .O(N__13667),
            .I(N__13473));
    LocalMux I__1961 (
            .O(N__13660),
            .I(N__13466));
    LocalMux I__1960 (
            .O(N__13651),
            .I(N__13466));
    Span4Mux_s2_h I__1959 (
            .O(N__13646),
            .I(N__13466));
    InMux I__1958 (
            .O(N__13645),
            .I(N__13463));
    InMux I__1957 (
            .O(N__13644),
            .I(N__13448));
    InMux I__1956 (
            .O(N__13643),
            .I(N__13448));
    InMux I__1955 (
            .O(N__13642),
            .I(N__13448));
    InMux I__1954 (
            .O(N__13641),
            .I(N__13448));
    InMux I__1953 (
            .O(N__13640),
            .I(N__13448));
    InMux I__1952 (
            .O(N__13639),
            .I(N__13448));
    InMux I__1951 (
            .O(N__13638),
            .I(N__13448));
    LocalMux I__1950 (
            .O(N__13635),
            .I(N__13443));
    LocalMux I__1949 (
            .O(N__13632),
            .I(N__13443));
    LocalMux I__1948 (
            .O(N__13619),
            .I(N__13436));
    LocalMux I__1947 (
            .O(N__13610),
            .I(N__13436));
    Span4Mux_s2_h I__1946 (
            .O(N__13607),
            .I(N__13436));
    LocalMux I__1945 (
            .O(N__13594),
            .I(N__13433));
    Span4Mux_s3_h I__1944 (
            .O(N__13591),
            .I(N__13426));
    LocalMux I__1943 (
            .O(N__13582),
            .I(N__13426));
    LocalMux I__1942 (
            .O(N__13567),
            .I(N__13426));
    LocalMux I__1941 (
            .O(N__13554),
            .I(N__13421));
    Span4Mux_s3_h I__1940 (
            .O(N__13551),
            .I(N__13421));
    InMux I__1939 (
            .O(N__13548),
            .I(N__13406));
    InMux I__1938 (
            .O(N__13545),
            .I(N__13406));
    InMux I__1937 (
            .O(N__13542),
            .I(N__13406));
    InMux I__1936 (
            .O(N__13539),
            .I(N__13406));
    InMux I__1935 (
            .O(N__13538),
            .I(N__13406));
    InMux I__1934 (
            .O(N__13537),
            .I(N__13406));
    InMux I__1933 (
            .O(N__13536),
            .I(N__13406));
    InMux I__1932 (
            .O(N__13533),
            .I(N__13393));
    InMux I__1931 (
            .O(N__13530),
            .I(N__13393));
    InMux I__1930 (
            .O(N__13527),
            .I(N__13393));
    InMux I__1929 (
            .O(N__13526),
            .I(N__13393));
    InMux I__1928 (
            .O(N__13525),
            .I(N__13393));
    InMux I__1927 (
            .O(N__13524),
            .I(N__13393));
    InMux I__1926 (
            .O(N__13523),
            .I(N__13378));
    InMux I__1925 (
            .O(N__13520),
            .I(N__13378));
    InMux I__1924 (
            .O(N__13517),
            .I(N__13378));
    InMux I__1923 (
            .O(N__13514),
            .I(N__13378));
    InMux I__1922 (
            .O(N__13513),
            .I(N__13378));
    InMux I__1921 (
            .O(N__13512),
            .I(N__13378));
    InMux I__1920 (
            .O(N__13511),
            .I(N__13378));
    InMux I__1919 (
            .O(N__13508),
            .I(N__13373));
    InMux I__1918 (
            .O(N__13507),
            .I(N__13373));
    InMux I__1917 (
            .O(N__13506),
            .I(N__13358));
    InMux I__1916 (
            .O(N__13505),
            .I(N__13358));
    InMux I__1915 (
            .O(N__13504),
            .I(N__13358));
    InMux I__1914 (
            .O(N__13503),
            .I(N__13358));
    InMux I__1913 (
            .O(N__13502),
            .I(N__13358));
    InMux I__1912 (
            .O(N__13501),
            .I(N__13358));
    InMux I__1911 (
            .O(N__13500),
            .I(N__13358));
    LocalMux I__1910 (
            .O(N__13497),
            .I(N__13351));
    LocalMux I__1909 (
            .O(N__13482),
            .I(N__13351));
    Span4Mux_v I__1908 (
            .O(N__13473),
            .I(N__13351));
    Span4Mux_h I__1907 (
            .O(N__13466),
            .I(N__13348));
    LocalMux I__1906 (
            .O(N__13463),
            .I(N__13339));
    LocalMux I__1905 (
            .O(N__13448),
            .I(N__13339));
    Span4Mux_h I__1904 (
            .O(N__13443),
            .I(N__13339));
    Span4Mux_h I__1903 (
            .O(N__13436),
            .I(N__13339));
    Span4Mux_s3_h I__1902 (
            .O(N__13433),
            .I(N__13332));
    Span4Mux_v I__1901 (
            .O(N__13426),
            .I(N__13332));
    Span4Mux_v I__1900 (
            .O(N__13421),
            .I(N__13332));
    LocalMux I__1899 (
            .O(N__13406),
            .I(n29));
    LocalMux I__1898 (
            .O(N__13393),
            .I(n29));
    LocalMux I__1897 (
            .O(N__13378),
            .I(n29));
    LocalMux I__1896 (
            .O(N__13373),
            .I(n29));
    LocalMux I__1895 (
            .O(N__13358),
            .I(n29));
    Odrv4 I__1894 (
            .O(N__13351),
            .I(n29));
    Odrv4 I__1893 (
            .O(N__13348),
            .I(n29));
    Odrv4 I__1892 (
            .O(N__13339),
            .I(n29));
    Odrv4 I__1891 (
            .O(N__13332),
            .I(n29));
    CascadeMux I__1890 (
            .O(N__13313),
            .I(\tok.n2_adj_685_cascade_ ));
    InMux I__1889 (
            .O(N__13310),
            .I(N__13307));
    LocalMux I__1888 (
            .O(N__13307),
            .I(\tok.n14_adj_686 ));
    InMux I__1887 (
            .O(N__13304),
            .I(N__13301));
    LocalMux I__1886 (
            .O(N__13301),
            .I(N__13297));
    InMux I__1885 (
            .O(N__13300),
            .I(N__13294));
    Odrv4 I__1884 (
            .O(N__13297),
            .I(sender_1));
    LocalMux I__1883 (
            .O(N__13294),
            .I(sender_1));
    IoInMux I__1882 (
            .O(N__13289),
            .I(N__13286));
    LocalMux I__1881 (
            .O(N__13286),
            .I(N__13283));
    Odrv4 I__1880 (
            .O(N__13283),
            .I(tx_c));
    InMux I__1879 (
            .O(N__13280),
            .I(N__13277));
    LocalMux I__1878 (
            .O(N__13277),
            .I(reset_c));
    InMux I__1877 (
            .O(N__13274),
            .I(N__13268));
    InMux I__1876 (
            .O(N__13273),
            .I(N__13268));
    LocalMux I__1875 (
            .O(N__13268),
            .I(\tok.A_stk.tail_63 ));
    InMux I__1874 (
            .O(N__13265),
            .I(N__13259));
    InMux I__1873 (
            .O(N__13264),
            .I(N__13259));
    LocalMux I__1872 (
            .O(N__13259),
            .I(\tok.A_stk.tail_47 ));
    InMux I__1871 (
            .O(N__13256),
            .I(N__13253));
    LocalMux I__1870 (
            .O(N__13253),
            .I(N__13250));
    Odrv4 I__1869 (
            .O(N__13250),
            .I(\tok.n6_adj_667 ));
    CascadeMux I__1868 (
            .O(N__13247),
            .I(N__13244));
    InMux I__1867 (
            .O(N__13244),
            .I(N__13241));
    LocalMux I__1866 (
            .O(N__13241),
            .I(\tok.n294 ));
    InMux I__1865 (
            .O(N__13238),
            .I(N__13235));
    LocalMux I__1864 (
            .O(N__13235),
            .I(N__13232));
    Span4Mux_h I__1863 (
            .O(N__13232),
            .I(N__13229));
    Span4Mux_h I__1862 (
            .O(N__13229),
            .I(N__13226));
    Sp12to4 I__1861 (
            .O(N__13226),
            .I(N__13223));
    Odrv12 I__1860 (
            .O(N__13223),
            .I(\tok.table_wr_data_3 ));
    CascadeMux I__1859 (
            .O(N__13220),
            .I(N__13217));
    InMux I__1858 (
            .O(N__13217),
            .I(N__13214));
    LocalMux I__1857 (
            .O(N__13214),
            .I(\tok.n298 ));
    CascadeMux I__1856 (
            .O(N__13211),
            .I(N__13208));
    InMux I__1855 (
            .O(N__13208),
            .I(N__13205));
    LocalMux I__1854 (
            .O(N__13205),
            .I(\tok.n289 ));
    InMux I__1853 (
            .O(N__13202),
            .I(N__13199));
    LocalMux I__1852 (
            .O(N__13199),
            .I(\tok.n6_adj_814 ));
    CascadeMux I__1851 (
            .O(N__13196),
            .I(\tok.n34_cascade_ ));
    InMux I__1850 (
            .O(N__13193),
            .I(N__13190));
    LocalMux I__1849 (
            .O(N__13190),
            .I(N__13187));
    Span4Mux_h I__1848 (
            .O(N__13187),
            .I(N__13184));
    Odrv4 I__1847 (
            .O(N__13184),
            .I(\tok.n13 ));
    InMux I__1846 (
            .O(N__13181),
            .I(N__13178));
    LocalMux I__1845 (
            .O(N__13178),
            .I(\tok.n4656 ));
    CascadeMux I__1844 (
            .O(N__13175),
            .I(\tok.n20_adj_754_cascade_ ));
    InMux I__1843 (
            .O(N__13172),
            .I(N__13169));
    LocalMux I__1842 (
            .O(N__13169),
            .I(N__13166));
    Odrv4 I__1841 (
            .O(N__13166),
            .I(\tok.n9_adj_749 ));
    InMux I__1840 (
            .O(N__13163),
            .I(N__13160));
    LocalMux I__1839 (
            .O(N__13160),
            .I(N__13157));
    Span4Mux_v I__1838 (
            .O(N__13157),
            .I(N__13154));
    Span4Mux_h I__1837 (
            .O(N__13154),
            .I(N__13151));
    Span4Mux_s1_h I__1836 (
            .O(N__13151),
            .I(N__13148));
    Odrv4 I__1835 (
            .O(N__13148),
            .I(\tok.table_rd_15 ));
    InMux I__1834 (
            .O(N__13145),
            .I(N__13142));
    LocalMux I__1833 (
            .O(N__13142),
            .I(\tok.n16_adj_751 ));
    InMux I__1832 (
            .O(N__13139),
            .I(N__13136));
    LocalMux I__1831 (
            .O(N__13136),
            .I(\tok.n17_adj_774 ));
    InMux I__1830 (
            .O(N__13133),
            .I(N__13130));
    LocalMux I__1829 (
            .O(N__13130),
            .I(N__13127));
    Odrv4 I__1828 (
            .O(N__13127),
            .I(\tok.n10_adj_705 ));
    InMux I__1827 (
            .O(N__13124),
            .I(N__13121));
    LocalMux I__1826 (
            .O(N__13121),
            .I(\tok.n6_adj_692 ));
    CascadeMux I__1825 (
            .O(N__13118),
            .I(\tok.n13_adj_688_cascade_ ));
    InMux I__1824 (
            .O(N__13115),
            .I(N__13112));
    LocalMux I__1823 (
            .O(N__13112),
            .I(\tok.n12_adj_687 ));
    InMux I__1822 (
            .O(N__13109),
            .I(N__13106));
    LocalMux I__1821 (
            .O(N__13106),
            .I(N__13103));
    Odrv4 I__1820 (
            .O(N__13103),
            .I(\tok.n4674 ));
    CascadeMux I__1819 (
            .O(N__13100),
            .I(\tok.n20_adj_693_cascade_ ));
    InMux I__1818 (
            .O(N__13097),
            .I(\tok.n3949 ));
    InMux I__1817 (
            .O(N__13094),
            .I(\tok.n3950 ));
    InMux I__1816 (
            .O(N__13091),
            .I(\tok.n3951 ));
    InMux I__1815 (
            .O(N__13088),
            .I(\tok.n3952 ));
    InMux I__1814 (
            .O(N__13085),
            .I(\tok.n3953 ));
    InMux I__1813 (
            .O(N__13082),
            .I(\tok.n3954 ));
    CascadeMux I__1812 (
            .O(N__13079),
            .I(\tok.n2_adj_739_cascade_ ));
    InMux I__1811 (
            .O(N__13076),
            .I(N__13073));
    LocalMux I__1810 (
            .O(N__13073),
            .I(N__13070));
    Span4Mux_v I__1809 (
            .O(N__13070),
            .I(N__13067));
    Odrv4 I__1808 (
            .O(N__13067),
            .I(\tok.n6_adj_753 ));
    CascadeMux I__1807 (
            .O(N__13064),
            .I(\tok.n14_adj_741_cascade_ ));
    InMux I__1806 (
            .O(N__13061),
            .I(N__13058));
    LocalMux I__1805 (
            .O(N__13058),
            .I(N__13055));
    Span4Mux_h I__1804 (
            .O(N__13055),
            .I(N__13052));
    Odrv4 I__1803 (
            .O(N__13052),
            .I(\tok.n13_adj_748 ));
    InMux I__1802 (
            .O(N__13049),
            .I(\tok.n3940 ));
    InMux I__1801 (
            .O(N__13046),
            .I(\tok.n3941 ));
    InMux I__1800 (
            .O(N__13043),
            .I(\tok.n3942 ));
    InMux I__1799 (
            .O(N__13040),
            .I(\tok.n3943 ));
    InMux I__1798 (
            .O(N__13037),
            .I(\tok.n3944 ));
    InMux I__1797 (
            .O(N__13034),
            .I(\tok.n3945 ));
    InMux I__1796 (
            .O(N__13031),
            .I(N__13028));
    LocalMux I__1795 (
            .O(N__13028),
            .I(N__13025));
    Odrv12 I__1794 (
            .O(N__13025),
            .I(\tok.n10_adj_764 ));
    InMux I__1793 (
            .O(N__13022),
            .I(\tok.n3946 ));
    InMux I__1792 (
            .O(N__13019),
            .I(bfn_5_9_0_));
    InMux I__1791 (
            .O(N__13016),
            .I(\tok.n3948 ));
    CascadeMux I__1790 (
            .O(N__13013),
            .I(N__13010));
    InMux I__1789 (
            .O(N__13010),
            .I(N__13004));
    InMux I__1788 (
            .O(N__13009),
            .I(N__13004));
    LocalMux I__1787 (
            .O(N__13004),
            .I(\tok.A_stk.tail_4 ));
    CascadeMux I__1786 (
            .O(N__13001),
            .I(N__12998));
    InMux I__1785 (
            .O(N__12998),
            .I(N__12995));
    LocalMux I__1784 (
            .O(N__12995),
            .I(\tok.n23_adj_677 ));
    InMux I__1783 (
            .O(N__12992),
            .I(N__12989));
    LocalMux I__1782 (
            .O(N__12989),
            .I(\tok.n24 ));
    InMux I__1781 (
            .O(N__12986),
            .I(N__12983));
    LocalMux I__1780 (
            .O(N__12983),
            .I(\tok.n26_adj_805 ));
    CascadeMux I__1779 (
            .O(N__12980),
            .I(\tok.n30_adj_824_cascade_ ));
    InMux I__1778 (
            .O(N__12977),
            .I(N__12974));
    LocalMux I__1777 (
            .O(N__12974),
            .I(\tok.found_slot_N_145 ));
    CascadeMux I__1776 (
            .O(N__12971),
            .I(\tok.n4642_cascade_ ));
    InMux I__1775 (
            .O(N__12968),
            .I(N__12964));
    InMux I__1774 (
            .O(N__12967),
            .I(N__12961));
    LocalMux I__1773 (
            .O(N__12964),
            .I(N__12958));
    LocalMux I__1772 (
            .O(N__12961),
            .I(\tok.key_rd_13 ));
    Odrv4 I__1771 (
            .O(N__12958),
            .I(\tok.key_rd_13 ));
    InMux I__1770 (
            .O(N__12953),
            .I(N__12950));
    LocalMux I__1769 (
            .O(N__12950),
            .I(\tok.n14_adj_804 ));
    InMux I__1768 (
            .O(N__12947),
            .I(N__12944));
    LocalMux I__1767 (
            .O(N__12944),
            .I(\tok.n27_adj_734 ));
    CascadeMux I__1766 (
            .O(N__12941),
            .I(N__12937));
    InMux I__1765 (
            .O(N__12940),
            .I(N__12934));
    InMux I__1764 (
            .O(N__12937),
            .I(N__12931));
    LocalMux I__1763 (
            .O(N__12934),
            .I(N__12926));
    LocalMux I__1762 (
            .O(N__12931),
            .I(N__12926));
    Odrv4 I__1761 (
            .O(N__12926),
            .I(\tok.key_rd_12 ));
    CascadeMux I__1760 (
            .O(N__12923),
            .I(N__12920));
    InMux I__1759 (
            .O(N__12920),
            .I(N__12916));
    InMux I__1758 (
            .O(N__12919),
            .I(N__12913));
    LocalMux I__1757 (
            .O(N__12916),
            .I(N__12910));
    LocalMux I__1756 (
            .O(N__12913),
            .I(N__12907));
    Odrv12 I__1755 (
            .O(N__12910),
            .I(\tok.key_rd_10 ));
    Odrv4 I__1754 (
            .O(N__12907),
            .I(\tok.key_rd_10 ));
    InMux I__1753 (
            .O(N__12902),
            .I(N__12899));
    LocalMux I__1752 (
            .O(N__12899),
            .I(\tok.n21_adj_714 ));
    InMux I__1751 (
            .O(N__12896),
            .I(N__12890));
    InMux I__1750 (
            .O(N__12895),
            .I(N__12890));
    LocalMux I__1749 (
            .O(N__12890),
            .I(N__12887));
    Span4Mux_h I__1748 (
            .O(N__12887),
            .I(N__12884));
    Odrv4 I__1747 (
            .O(N__12884),
            .I(\tok.key_rd_2 ));
    InMux I__1746 (
            .O(N__12881),
            .I(N__12878));
    LocalMux I__1745 (
            .O(N__12878),
            .I(N__12874));
    InMux I__1744 (
            .O(N__12877),
            .I(N__12871));
    Span4Mux_v I__1743 (
            .O(N__12874),
            .I(N__12868));
    LocalMux I__1742 (
            .O(N__12871),
            .I(N__12865));
    Span4Mux_h I__1741 (
            .O(N__12868),
            .I(N__12860));
    Span4Mux_v I__1740 (
            .O(N__12865),
            .I(N__12860));
    Odrv4 I__1739 (
            .O(N__12860),
            .I(\tok.key_rd_7 ));
    InMux I__1738 (
            .O(N__12857),
            .I(N__12854));
    LocalMux I__1737 (
            .O(N__12854),
            .I(\tok.n22 ));
    InMux I__1736 (
            .O(N__12851),
            .I(bfn_5_8_0_));
    InMux I__1735 (
            .O(N__12848),
            .I(N__12842));
    InMux I__1734 (
            .O(N__12847),
            .I(N__12842));
    LocalMux I__1733 (
            .O(N__12842),
            .I(\tok.A_stk.tail_21 ));
    CascadeMux I__1732 (
            .O(N__12839),
            .I(N__12836));
    InMux I__1731 (
            .O(N__12836),
            .I(N__12830));
    InMux I__1730 (
            .O(N__12835),
            .I(N__12830));
    LocalMux I__1729 (
            .O(N__12830),
            .I(\tok.A_stk.tail_5 ));
    InMux I__1728 (
            .O(N__12827),
            .I(N__12823));
    InMux I__1727 (
            .O(N__12826),
            .I(N__12820));
    LocalMux I__1726 (
            .O(N__12823),
            .I(N__12817));
    LocalMux I__1725 (
            .O(N__12820),
            .I(tail_116));
    Odrv4 I__1724 (
            .O(N__12817),
            .I(tail_116));
    CascadeMux I__1723 (
            .O(N__12812),
            .I(N__12809));
    InMux I__1722 (
            .O(N__12809),
            .I(N__12806));
    LocalMux I__1721 (
            .O(N__12806),
            .I(N__12802));
    InMux I__1720 (
            .O(N__12805),
            .I(N__12799));
    Sp12to4 I__1719 (
            .O(N__12802),
            .I(N__12796));
    LocalMux I__1718 (
            .O(N__12799),
            .I(tail_100));
    Odrv12 I__1717 (
            .O(N__12796),
            .I(tail_100));
    InMux I__1716 (
            .O(N__12791),
            .I(N__12785));
    InMux I__1715 (
            .O(N__12790),
            .I(N__12785));
    LocalMux I__1714 (
            .O(N__12785),
            .I(\tok.A_stk.tail_84 ));
    CascadeMux I__1713 (
            .O(N__12782),
            .I(N__12778));
    CascadeMux I__1712 (
            .O(N__12781),
            .I(N__12775));
    InMux I__1711 (
            .O(N__12778),
            .I(N__12770));
    InMux I__1710 (
            .O(N__12775),
            .I(N__12770));
    LocalMux I__1709 (
            .O(N__12770),
            .I(\tok.A_stk.tail_68 ));
    InMux I__1708 (
            .O(N__12767),
            .I(N__12761));
    InMux I__1707 (
            .O(N__12766),
            .I(N__12761));
    LocalMux I__1706 (
            .O(N__12761),
            .I(\tok.A_stk.tail_52 ));
    InMux I__1705 (
            .O(N__12758),
            .I(N__12752));
    InMux I__1704 (
            .O(N__12757),
            .I(N__12752));
    LocalMux I__1703 (
            .O(N__12752),
            .I(\tok.A_stk.tail_36 ));
    InMux I__1702 (
            .O(N__12749),
            .I(N__12743));
    InMux I__1701 (
            .O(N__12748),
            .I(N__12743));
    LocalMux I__1700 (
            .O(N__12743),
            .I(\tok.A_stk.tail_20 ));
    CascadeMux I__1699 (
            .O(N__12740),
            .I(N__12736));
    InMux I__1698 (
            .O(N__12739),
            .I(N__12733));
    InMux I__1697 (
            .O(N__12736),
            .I(N__12730));
    LocalMux I__1696 (
            .O(N__12733),
            .I(tail_117));
    LocalMux I__1695 (
            .O(N__12730),
            .I(tail_117));
    InMux I__1694 (
            .O(N__12725),
            .I(N__12721));
    InMux I__1693 (
            .O(N__12724),
            .I(N__12718));
    LocalMux I__1692 (
            .O(N__12721),
            .I(tail_101));
    LocalMux I__1691 (
            .O(N__12718),
            .I(tail_101));
    InMux I__1690 (
            .O(N__12713),
            .I(N__12707));
    InMux I__1689 (
            .O(N__12712),
            .I(N__12707));
    LocalMux I__1688 (
            .O(N__12707),
            .I(\tok.A_stk.tail_67 ));
    CascadeMux I__1687 (
            .O(N__12704),
            .I(N__12700));
    InMux I__1686 (
            .O(N__12703),
            .I(N__12697));
    InMux I__1685 (
            .O(N__12700),
            .I(N__12694));
    LocalMux I__1684 (
            .O(N__12697),
            .I(tail_99));
    LocalMux I__1683 (
            .O(N__12694),
            .I(tail_99));
    InMux I__1682 (
            .O(N__12689),
            .I(N__12683));
    InMux I__1681 (
            .O(N__12688),
            .I(N__12683));
    LocalMux I__1680 (
            .O(N__12683),
            .I(\tok.A_stk.tail_83 ));
    InMux I__1679 (
            .O(N__12680),
            .I(N__12676));
    InMux I__1678 (
            .O(N__12679),
            .I(N__12673));
    LocalMux I__1677 (
            .O(N__12676),
            .I(\tok.A_stk.tail_35 ));
    LocalMux I__1676 (
            .O(N__12673),
            .I(\tok.A_stk.tail_35 ));
    CascadeMux I__1675 (
            .O(N__12668),
            .I(N__12664));
    InMux I__1674 (
            .O(N__12667),
            .I(N__12661));
    InMux I__1673 (
            .O(N__12664),
            .I(N__12658));
    LocalMux I__1672 (
            .O(N__12661),
            .I(\tok.A_stk.tail_3 ));
    LocalMux I__1671 (
            .O(N__12658),
            .I(\tok.A_stk.tail_3 ));
    CascadeMux I__1670 (
            .O(N__12653),
            .I(N__12649));
    CascadeMux I__1669 (
            .O(N__12652),
            .I(N__12646));
    InMux I__1668 (
            .O(N__12649),
            .I(N__12643));
    InMux I__1667 (
            .O(N__12646),
            .I(N__12640));
    LocalMux I__1666 (
            .O(N__12643),
            .I(\tok.A_stk.tail_19 ));
    LocalMux I__1665 (
            .O(N__12640),
            .I(\tok.A_stk.tail_19 ));
    InMux I__1664 (
            .O(N__12635),
            .I(N__12631));
    InMux I__1663 (
            .O(N__12634),
            .I(N__12628));
    LocalMux I__1662 (
            .O(N__12631),
            .I(\tok.A_stk.tail_85 ));
    LocalMux I__1661 (
            .O(N__12628),
            .I(\tok.A_stk.tail_85 ));
    CascadeMux I__1660 (
            .O(N__12623),
            .I(N__12619));
    InMux I__1659 (
            .O(N__12622),
            .I(N__12616));
    InMux I__1658 (
            .O(N__12619),
            .I(N__12613));
    LocalMux I__1657 (
            .O(N__12616),
            .I(\tok.A_stk.tail_69 ));
    LocalMux I__1656 (
            .O(N__12613),
            .I(\tok.A_stk.tail_69 ));
    CascadeMux I__1655 (
            .O(N__12608),
            .I(N__12604));
    CascadeMux I__1654 (
            .O(N__12607),
            .I(N__12601));
    InMux I__1653 (
            .O(N__12604),
            .I(N__12596));
    InMux I__1652 (
            .O(N__12601),
            .I(N__12596));
    LocalMux I__1651 (
            .O(N__12596),
            .I(\tok.A_stk.tail_53 ));
    InMux I__1650 (
            .O(N__12593),
            .I(N__12587));
    InMux I__1649 (
            .O(N__12592),
            .I(N__12587));
    LocalMux I__1648 (
            .O(N__12587),
            .I(N__12584));
    Odrv4 I__1647 (
            .O(N__12584),
            .I(\tok.A_stk.tail_37 ));
    CascadeMux I__1646 (
            .O(N__12581),
            .I(N__12577));
    InMux I__1645 (
            .O(N__12580),
            .I(N__12572));
    InMux I__1644 (
            .O(N__12577),
            .I(N__12572));
    LocalMux I__1643 (
            .O(N__12572),
            .I(\tok.A_stk.tail_49 ));
    InMux I__1642 (
            .O(N__12569),
            .I(N__12563));
    InMux I__1641 (
            .O(N__12568),
            .I(N__12563));
    LocalMux I__1640 (
            .O(N__12563),
            .I(\tok.A_stk.tail_65 ));
    InMux I__1639 (
            .O(N__12560),
            .I(N__12554));
    InMux I__1638 (
            .O(N__12559),
            .I(N__12554));
    LocalMux I__1637 (
            .O(N__12554),
            .I(\tok.A_stk.tail_81 ));
    InMux I__1636 (
            .O(N__12551),
            .I(N__12545));
    InMux I__1635 (
            .O(N__12550),
            .I(N__12545));
    LocalMux I__1634 (
            .O(N__12545),
            .I(\tok.A_stk.tail_1 ));
    InMux I__1633 (
            .O(N__12542),
            .I(N__12538));
    InMux I__1632 (
            .O(N__12541),
            .I(N__12535));
    LocalMux I__1631 (
            .O(N__12538),
            .I(tail_115));
    LocalMux I__1630 (
            .O(N__12535),
            .I(tail_115));
    InMux I__1629 (
            .O(N__12530),
            .I(N__12524));
    InMux I__1628 (
            .O(N__12529),
            .I(N__12524));
    LocalMux I__1627 (
            .O(N__12524),
            .I(\tok.A_stk.tail_51 ));
    InMux I__1626 (
            .O(N__12521),
            .I(N__12515));
    InMux I__1625 (
            .O(N__12520),
            .I(N__12515));
    LocalMux I__1624 (
            .O(N__12515),
            .I(\tok.A_stk.tail_92 ));
    InMux I__1623 (
            .O(N__12512),
            .I(N__12506));
    InMux I__1622 (
            .O(N__12511),
            .I(N__12506));
    LocalMux I__1621 (
            .O(N__12506),
            .I(\tok.A_stk.tail_76 ));
    CascadeMux I__1620 (
            .O(N__12503),
            .I(N__12500));
    InMux I__1619 (
            .O(N__12500),
            .I(N__12496));
    InMux I__1618 (
            .O(N__12499),
            .I(N__12493));
    LocalMux I__1617 (
            .O(N__12496),
            .I(N__12490));
    LocalMux I__1616 (
            .O(N__12493),
            .I(\tok.A_stk.tail_60 ));
    Odrv4 I__1615 (
            .O(N__12490),
            .I(\tok.A_stk.tail_60 ));
    CascadeMux I__1614 (
            .O(N__12485),
            .I(N__12481));
    CascadeMux I__1613 (
            .O(N__12484),
            .I(N__12478));
    InMux I__1612 (
            .O(N__12481),
            .I(N__12473));
    InMux I__1611 (
            .O(N__12478),
            .I(N__12473));
    LocalMux I__1610 (
            .O(N__12473),
            .I(\tok.A_stk.tail_44 ));
    CascadeMux I__1609 (
            .O(N__12470),
            .I(N__12466));
    CascadeMux I__1608 (
            .O(N__12469),
            .I(N__12463));
    InMux I__1607 (
            .O(N__12466),
            .I(N__12458));
    InMux I__1606 (
            .O(N__12463),
            .I(N__12458));
    LocalMux I__1605 (
            .O(N__12458),
            .I(\tok.A_stk.tail_28 ));
    InMux I__1604 (
            .O(N__12455),
            .I(N__12451));
    InMux I__1603 (
            .O(N__12454),
            .I(N__12448));
    LocalMux I__1602 (
            .O(N__12451),
            .I(\tok.A_stk.tail_12 ));
    LocalMux I__1601 (
            .O(N__12448),
            .I(\tok.A_stk.tail_12 ));
    CascadeMux I__1600 (
            .O(N__12443),
            .I(N__12439));
    InMux I__1599 (
            .O(N__12442),
            .I(N__12434));
    InMux I__1598 (
            .O(N__12439),
            .I(N__12434));
    LocalMux I__1597 (
            .O(N__12434),
            .I(\tok.A_stk.tail_17 ));
    InMux I__1596 (
            .O(N__12431),
            .I(N__12425));
    InMux I__1595 (
            .O(N__12430),
            .I(N__12425));
    LocalMux I__1594 (
            .O(N__12425),
            .I(\tok.A_stk.tail_33 ));
    CascadeMux I__1593 (
            .O(N__12422),
            .I(N__12419));
    InMux I__1592 (
            .O(N__12419),
            .I(N__12416));
    LocalMux I__1591 (
            .O(N__12416),
            .I(N__12413));
    Odrv4 I__1590 (
            .O(N__12413),
            .I(\tok.n290 ));
    InMux I__1589 (
            .O(N__12410),
            .I(N__12407));
    LocalMux I__1588 (
            .O(N__12407),
            .I(N__12404));
    Odrv4 I__1587 (
            .O(N__12404),
            .I(\tok.n6_adj_701 ));
    InMux I__1586 (
            .O(N__12401),
            .I(\tok.n3921 ));
    InMux I__1585 (
            .O(N__12398),
            .I(\tok.n3922 ));
    CascadeMux I__1584 (
            .O(N__12395),
            .I(N__12392));
    InMux I__1583 (
            .O(N__12392),
            .I(N__12389));
    LocalMux I__1582 (
            .O(N__12389),
            .I(N__12386));
    Odrv12 I__1581 (
            .O(N__12386),
            .I(\tok.n288 ));
    InMux I__1580 (
            .O(N__12383),
            .I(\tok.n3923 ));
    InMux I__1579 (
            .O(N__12380),
            .I(bfn_4_13_0_));
    InMux I__1578 (
            .O(N__12377),
            .I(N__12374));
    LocalMux I__1577 (
            .O(N__12374),
            .I(\tok.n292 ));
    InMux I__1576 (
            .O(N__12371),
            .I(N__12368));
    LocalMux I__1575 (
            .O(N__12368),
            .I(\tok.n287 ));
    CascadeMux I__1574 (
            .O(N__12365),
            .I(N__12361));
    CascadeMux I__1573 (
            .O(N__12364),
            .I(N__12358));
    InMux I__1572 (
            .O(N__12361),
            .I(N__12355));
    InMux I__1571 (
            .O(N__12358),
            .I(N__12352));
    LocalMux I__1570 (
            .O(N__12355),
            .I(tail_124));
    LocalMux I__1569 (
            .O(N__12352),
            .I(tail_124));
    CascadeMux I__1568 (
            .O(N__12347),
            .I(N__12343));
    InMux I__1567 (
            .O(N__12346),
            .I(N__12340));
    InMux I__1566 (
            .O(N__12343),
            .I(N__12337));
    LocalMux I__1565 (
            .O(N__12340),
            .I(tail_108));
    LocalMux I__1564 (
            .O(N__12337),
            .I(tail_108));
    InMux I__1563 (
            .O(N__12332),
            .I(\tok.n3913 ));
    InMux I__1562 (
            .O(N__12329),
            .I(\tok.n3914 ));
    InMux I__1561 (
            .O(N__12326),
            .I(\tok.n3915 ));
    InMux I__1560 (
            .O(N__12323),
            .I(N__12320));
    LocalMux I__1559 (
            .O(N__12320),
            .I(N__12317));
    Odrv4 I__1558 (
            .O(N__12317),
            .I(\tok.n295 ));
    InMux I__1557 (
            .O(N__12314),
            .I(N__12311));
    LocalMux I__1556 (
            .O(N__12311),
            .I(N__12308));
    Span4Mux_h I__1555 (
            .O(N__12308),
            .I(N__12305));
    Odrv4 I__1554 (
            .O(N__12305),
            .I(\tok.n6_adj_768 ));
    InMux I__1553 (
            .O(N__12302),
            .I(\tok.n3916 ));
    InMux I__1552 (
            .O(N__12299),
            .I(bfn_4_12_0_));
    InMux I__1551 (
            .O(N__12296),
            .I(\tok.n3918 ));
    InMux I__1550 (
            .O(N__12293),
            .I(\tok.n3919 ));
    CascadeMux I__1549 (
            .O(N__12290),
            .I(N__12287));
    InMux I__1548 (
            .O(N__12287),
            .I(N__12284));
    LocalMux I__1547 (
            .O(N__12284),
            .I(N__12281));
    Span4Mux_v I__1546 (
            .O(N__12281),
            .I(N__12278));
    Odrv4 I__1545 (
            .O(N__12278),
            .I(\tok.n291 ));
    InMux I__1544 (
            .O(N__12275),
            .I(\tok.n3920 ));
    InMux I__1543 (
            .O(N__12272),
            .I(N__12263));
    InMux I__1542 (
            .O(N__12271),
            .I(N__12263));
    InMux I__1541 (
            .O(N__12270),
            .I(N__12263));
    LocalMux I__1540 (
            .O(N__12263),
            .I(capture_7));
    InMux I__1539 (
            .O(N__12260),
            .I(N__12257));
    LocalMux I__1538 (
            .O(N__12257),
            .I(N__12252));
    InMux I__1537 (
            .O(N__12256),
            .I(N__12247));
    InMux I__1536 (
            .O(N__12255),
            .I(N__12247));
    Odrv12 I__1535 (
            .O(N__12252),
            .I(capture_6));
    LocalMux I__1534 (
            .O(N__12247),
            .I(capture_6));
    SRMux I__1533 (
            .O(N__12242),
            .I(N__12236));
    SRMux I__1532 (
            .O(N__12241),
            .I(N__12233));
    InMux I__1531 (
            .O(N__12240),
            .I(N__12227));
    InMux I__1530 (
            .O(N__12239),
            .I(N__12227));
    LocalMux I__1529 (
            .O(N__12236),
            .I(N__12224));
    LocalMux I__1528 (
            .O(N__12233),
            .I(N__12221));
    InMux I__1527 (
            .O(N__12232),
            .I(N__12218));
    LocalMux I__1526 (
            .O(N__12227),
            .I(N__12215));
    Span4Mux_h I__1525 (
            .O(N__12224),
            .I(N__12210));
    Span4Mux_v I__1524 (
            .O(N__12221),
            .I(N__12210));
    LocalMux I__1523 (
            .O(N__12218),
            .I(N__12207));
    Span4Mux_v I__1522 (
            .O(N__12215),
            .I(N__12203));
    Span4Mux_s1_h I__1521 (
            .O(N__12210),
            .I(N__12198));
    Span4Mux_h I__1520 (
            .O(N__12207),
            .I(N__12198));
    InMux I__1519 (
            .O(N__12206),
            .I(N__12195));
    Span4Mux_h I__1518 (
            .O(N__12203),
            .I(N__12192));
    Odrv4 I__1517 (
            .O(N__12198),
            .I(txtick));
    LocalMux I__1516 (
            .O(N__12195),
            .I(txtick));
    Odrv4 I__1515 (
            .O(N__12192),
            .I(txtick));
    InMux I__1514 (
            .O(N__12185),
            .I(bfn_4_11_0_));
    InMux I__1513 (
            .O(N__12182),
            .I(\tok.n3910 ));
    InMux I__1512 (
            .O(N__12179),
            .I(N__12176));
    LocalMux I__1511 (
            .O(N__12176),
            .I(N__12173));
    Odrv4 I__1510 (
            .O(N__12173),
            .I(\tok.n300 ));
    InMux I__1509 (
            .O(N__12170),
            .I(\tok.n3911 ));
    InMux I__1508 (
            .O(N__12167),
            .I(\tok.n3912 ));
    CascadeMux I__1507 (
            .O(N__12164),
            .I(\tok.uart.n6_cascade_ ));
    CascadeMux I__1506 (
            .O(N__12161),
            .I(n23_cascade_));
    CascadeMux I__1505 (
            .O(N__12158),
            .I(N__12155));
    InMux I__1504 (
            .O(N__12155),
            .I(N__12144));
    InMux I__1503 (
            .O(N__12154),
            .I(N__12144));
    InMux I__1502 (
            .O(N__12153),
            .I(N__12144));
    InMux I__1501 (
            .O(N__12152),
            .I(N__12139));
    InMux I__1500 (
            .O(N__12151),
            .I(N__12139));
    LocalMux I__1499 (
            .O(N__12144),
            .I(N__12136));
    LocalMux I__1498 (
            .O(N__12139),
            .I(\tok.uart.sentbits_0 ));
    Odrv4 I__1497 (
            .O(N__12136),
            .I(\tok.uart.sentbits_0 ));
    InMux I__1496 (
            .O(N__12131),
            .I(N__12121));
    InMux I__1495 (
            .O(N__12130),
            .I(N__12121));
    InMux I__1494 (
            .O(N__12129),
            .I(N__12121));
    InMux I__1493 (
            .O(N__12128),
            .I(N__12118));
    LocalMux I__1492 (
            .O(N__12121),
            .I(N__12115));
    LocalMux I__1491 (
            .O(N__12118),
            .I(\tok.uart.sentbits_1 ));
    Odrv4 I__1490 (
            .O(N__12115),
            .I(\tok.uart.sentbits_1 ));
    CEMux I__1489 (
            .O(N__12110),
            .I(N__12106));
    CEMux I__1488 (
            .O(N__12109),
            .I(N__12103));
    LocalMux I__1487 (
            .O(N__12106),
            .I(N__12100));
    LocalMux I__1486 (
            .O(N__12103),
            .I(N__12097));
    Odrv4 I__1485 (
            .O(N__12100),
            .I(\tok.uart.n978 ));
    Odrv4 I__1484 (
            .O(N__12097),
            .I(\tok.uart.n978 ));
    SRMux I__1483 (
            .O(N__12092),
            .I(N__12089));
    LocalMux I__1482 (
            .O(N__12089),
            .I(N__12085));
    SRMux I__1481 (
            .O(N__12088),
            .I(N__12082));
    Span4Mux_s3_h I__1480 (
            .O(N__12085),
            .I(N__12077));
    LocalMux I__1479 (
            .O(N__12082),
            .I(N__12077));
    Odrv4 I__1478 (
            .O(N__12077),
            .I(\tok.uart.n1083 ));
    InMux I__1477 (
            .O(N__12074),
            .I(N__12070));
    InMux I__1476 (
            .O(N__12073),
            .I(N__12067));
    LocalMux I__1475 (
            .O(N__12070),
            .I(\tok.key_rd_14 ));
    LocalMux I__1474 (
            .O(N__12067),
            .I(\tok.key_rd_14 ));
    InMux I__1473 (
            .O(N__12062),
            .I(N__12058));
    InMux I__1472 (
            .O(N__12061),
            .I(N__12055));
    LocalMux I__1471 (
            .O(N__12058),
            .I(\tok.key_rd_11 ));
    LocalMux I__1470 (
            .O(N__12055),
            .I(\tok.key_rd_11 ));
    InMux I__1469 (
            .O(N__12050),
            .I(N__12047));
    LocalMux I__1468 (
            .O(N__12047),
            .I(N__12044));
    Odrv4 I__1467 (
            .O(N__12044),
            .I(\tok.table_wr_data_11 ));
    CascadeMux I__1466 (
            .O(N__12041),
            .I(N__12038));
    InMux I__1465 (
            .O(N__12038),
            .I(N__12034));
    InMux I__1464 (
            .O(N__12037),
            .I(N__12031));
    LocalMux I__1463 (
            .O(N__12034),
            .I(\tok.key_rd_15 ));
    LocalMux I__1462 (
            .O(N__12031),
            .I(\tok.key_rd_15 ));
    InMux I__1461 (
            .O(N__12026),
            .I(N__12022));
    InMux I__1460 (
            .O(N__12025),
            .I(N__12019));
    LocalMux I__1459 (
            .O(N__12022),
            .I(\tok.key_rd_9 ));
    LocalMux I__1458 (
            .O(N__12019),
            .I(\tok.key_rd_9 ));
    InMux I__1457 (
            .O(N__12014),
            .I(N__12011));
    LocalMux I__1456 (
            .O(N__12011),
            .I(N__12008));
    Odrv4 I__1455 (
            .O(N__12008),
            .I(\tok.table_wr_data_7 ));
    InMux I__1454 (
            .O(N__12005),
            .I(N__12002));
    LocalMux I__1453 (
            .O(N__12002),
            .I(N__11999));
    Span4Mux_h I__1452 (
            .O(N__11999),
            .I(N__11996));
    Odrv4 I__1451 (
            .O(N__11996),
            .I(\tok.table_wr_data_4 ));
    InMux I__1450 (
            .O(N__11993),
            .I(N__11990));
    LocalMux I__1449 (
            .O(N__11990),
            .I(N__11987));
    Span4Mux_v I__1448 (
            .O(N__11987),
            .I(N__11984));
    Odrv4 I__1447 (
            .O(N__11984),
            .I(\tok.table_wr_data_1 ));
    InMux I__1446 (
            .O(N__11981),
            .I(N__11978));
    LocalMux I__1445 (
            .O(N__11978),
            .I(N__11975));
    Span4Mux_v I__1444 (
            .O(N__11975),
            .I(N__11972));
    Odrv4 I__1443 (
            .O(N__11972),
            .I(\tok.n15_adj_771 ));
    CascadeMux I__1442 (
            .O(N__11969),
            .I(N__11965));
    CascadeMux I__1441 (
            .O(N__11968),
            .I(N__11962));
    InMux I__1440 (
            .O(N__11965),
            .I(N__11957));
    InMux I__1439 (
            .O(N__11962),
            .I(N__11957));
    LocalMux I__1438 (
            .O(N__11957),
            .I(\tok.A_stk.tail_38 ));
    CascadeMux I__1437 (
            .O(N__11954),
            .I(N__11950));
    CascadeMux I__1436 (
            .O(N__11953),
            .I(N__11947));
    InMux I__1435 (
            .O(N__11950),
            .I(N__11942));
    InMux I__1434 (
            .O(N__11947),
            .I(N__11942));
    LocalMux I__1433 (
            .O(N__11942),
            .I(\tok.A_stk.tail_22 ));
    InMux I__1432 (
            .O(N__11939),
            .I(N__11933));
    InMux I__1431 (
            .O(N__11938),
            .I(N__11933));
    LocalMux I__1430 (
            .O(N__11933),
            .I(\tok.A_stk.tail_6 ));
    CascadeMux I__1429 (
            .O(N__11930),
            .I(\tok.n20_adj_803_cascade_ ));
    InMux I__1428 (
            .O(N__11927),
            .I(N__11921));
    InMux I__1427 (
            .O(N__11926),
            .I(N__11921));
    LocalMux I__1426 (
            .O(N__11921),
            .I(\tok.key_rd_5 ));
    InMux I__1425 (
            .O(N__11918),
            .I(N__11912));
    InMux I__1424 (
            .O(N__11917),
            .I(N__11912));
    LocalMux I__1423 (
            .O(N__11912),
            .I(\tok.key_rd_3 ));
    CascadeMux I__1422 (
            .O(N__11909),
            .I(N__11905));
    InMux I__1421 (
            .O(N__11908),
            .I(N__11900));
    InMux I__1420 (
            .O(N__11905),
            .I(N__11900));
    LocalMux I__1419 (
            .O(N__11900),
            .I(\tok.key_rd_8 ));
    InMux I__1418 (
            .O(N__11897),
            .I(N__11894));
    LocalMux I__1417 (
            .O(N__11894),
            .I(\tok.n28 ));
    CascadeMux I__1416 (
            .O(N__11891),
            .I(\tok.n25_cascade_ ));
    InMux I__1415 (
            .O(N__11888),
            .I(N__11885));
    LocalMux I__1414 (
            .O(N__11885),
            .I(\tok.n26 ));
    InMux I__1413 (
            .O(N__11882),
            .I(N__11876));
    InMux I__1412 (
            .O(N__11881),
            .I(N__11876));
    LocalMux I__1411 (
            .O(N__11876),
            .I(\tok.A_stk.tail_77 ));
    InMux I__1410 (
            .O(N__11873),
            .I(N__11867));
    InMux I__1409 (
            .O(N__11872),
            .I(N__11867));
    LocalMux I__1408 (
            .O(N__11867),
            .I(\tok.A_stk.tail_61 ));
    InMux I__1407 (
            .O(N__11864),
            .I(N__11858));
    InMux I__1406 (
            .O(N__11863),
            .I(N__11858));
    LocalMux I__1405 (
            .O(N__11858),
            .I(\tok.A_stk.tail_45 ));
    CascadeMux I__1404 (
            .O(N__11855),
            .I(N__11851));
    InMux I__1403 (
            .O(N__11854),
            .I(N__11846));
    InMux I__1402 (
            .O(N__11851),
            .I(N__11846));
    LocalMux I__1401 (
            .O(N__11846),
            .I(\tok.A_stk.tail_29 ));
    InMux I__1400 (
            .O(N__11843),
            .I(N__11839));
    InMux I__1399 (
            .O(N__11842),
            .I(N__11836));
    LocalMux I__1398 (
            .O(N__11839),
            .I(\tok.A_stk.tail_13 ));
    LocalMux I__1397 (
            .O(N__11836),
            .I(\tok.A_stk.tail_13 ));
    CascadeMux I__1396 (
            .O(N__11831),
            .I(N__11828));
    InMux I__1395 (
            .O(N__11828),
            .I(N__11824));
    InMux I__1394 (
            .O(N__11827),
            .I(N__11821));
    LocalMux I__1393 (
            .O(N__11824),
            .I(N__11818));
    LocalMux I__1392 (
            .O(N__11821),
            .I(tail_118));
    Odrv12 I__1391 (
            .O(N__11818),
            .I(tail_118));
    CascadeMux I__1390 (
            .O(N__11813),
            .I(N__11810));
    InMux I__1389 (
            .O(N__11810),
            .I(N__11806));
    CascadeMux I__1388 (
            .O(N__11809),
            .I(N__11803));
    LocalMux I__1387 (
            .O(N__11806),
            .I(N__11800));
    InMux I__1386 (
            .O(N__11803),
            .I(N__11797));
    Span4Mux_h I__1385 (
            .O(N__11800),
            .I(N__11794));
    LocalMux I__1384 (
            .O(N__11797),
            .I(tail_102));
    Odrv4 I__1383 (
            .O(N__11794),
            .I(tail_102));
    InMux I__1382 (
            .O(N__11789),
            .I(N__11783));
    InMux I__1381 (
            .O(N__11788),
            .I(N__11783));
    LocalMux I__1380 (
            .O(N__11783),
            .I(\tok.A_stk.tail_86 ));
    InMux I__1379 (
            .O(N__11780),
            .I(N__11774));
    InMux I__1378 (
            .O(N__11779),
            .I(N__11774));
    LocalMux I__1377 (
            .O(N__11774),
            .I(\tok.A_stk.tail_70 ));
    CascadeMux I__1376 (
            .O(N__11771),
            .I(N__11767));
    InMux I__1375 (
            .O(N__11770),
            .I(N__11762));
    InMux I__1374 (
            .O(N__11767),
            .I(N__11762));
    LocalMux I__1373 (
            .O(N__11762),
            .I(\tok.A_stk.tail_54 ));
    CascadeMux I__1372 (
            .O(N__11759),
            .I(N__11756));
    InMux I__1371 (
            .O(N__11756),
            .I(N__11752));
    InMux I__1370 (
            .O(N__11755),
            .I(N__11749));
    LocalMux I__1369 (
            .O(N__11752),
            .I(tail_98));
    LocalMux I__1368 (
            .O(N__11749),
            .I(tail_98));
    CascadeMux I__1367 (
            .O(N__11744),
            .I(N__11740));
    InMux I__1366 (
            .O(N__11743),
            .I(N__11737));
    InMux I__1365 (
            .O(N__11740),
            .I(N__11734));
    LocalMux I__1364 (
            .O(N__11737),
            .I(tail_114));
    LocalMux I__1363 (
            .O(N__11734),
            .I(tail_114));
    InMux I__1362 (
            .O(N__11729),
            .I(N__11725));
    InMux I__1361 (
            .O(N__11728),
            .I(N__11722));
    LocalMux I__1360 (
            .O(N__11725),
            .I(tail_125));
    LocalMux I__1359 (
            .O(N__11722),
            .I(tail_125));
    InMux I__1358 (
            .O(N__11717),
            .I(N__11713));
    InMux I__1357 (
            .O(N__11716),
            .I(N__11710));
    LocalMux I__1356 (
            .O(N__11713),
            .I(tail_109));
    LocalMux I__1355 (
            .O(N__11710),
            .I(tail_109));
    CascadeMux I__1354 (
            .O(N__11705),
            .I(N__11702));
    InMux I__1353 (
            .O(N__11702),
            .I(N__11696));
    InMux I__1352 (
            .O(N__11701),
            .I(N__11696));
    LocalMux I__1351 (
            .O(N__11696),
            .I(\tok.A_stk.tail_93 ));
    InMux I__1350 (
            .O(N__11693),
            .I(N__11687));
    InMux I__1349 (
            .O(N__11692),
            .I(N__11687));
    LocalMux I__1348 (
            .O(N__11687),
            .I(\tok.A_stk.tail_18 ));
    InMux I__1347 (
            .O(N__11684),
            .I(N__11678));
    InMux I__1346 (
            .O(N__11683),
            .I(N__11678));
    LocalMux I__1345 (
            .O(N__11678),
            .I(\tok.A_stk.tail_34 ));
    CascadeMux I__1344 (
            .O(N__11675),
            .I(N__11671));
    InMux I__1343 (
            .O(N__11674),
            .I(N__11666));
    InMux I__1342 (
            .O(N__11671),
            .I(N__11666));
    LocalMux I__1341 (
            .O(N__11666),
            .I(\tok.A_stk.tail_50 ));
    InMux I__1340 (
            .O(N__11663),
            .I(N__11657));
    InMux I__1339 (
            .O(N__11662),
            .I(N__11657));
    LocalMux I__1338 (
            .O(N__11657),
            .I(\tok.A_stk.tail_66 ));
    InMux I__1337 (
            .O(N__11654),
            .I(N__11648));
    InMux I__1336 (
            .O(N__11653),
            .I(N__11648));
    LocalMux I__1335 (
            .O(N__11648),
            .I(\tok.A_stk.tail_82 ));
    CascadeMux I__1334 (
            .O(N__11645),
            .I(N__11642));
    InMux I__1333 (
            .O(N__11642),
            .I(N__11638));
    InMux I__1332 (
            .O(N__11641),
            .I(N__11635));
    LocalMux I__1331 (
            .O(N__11638),
            .I(\tok.A_stk.tail_2 ));
    LocalMux I__1330 (
            .O(N__11635),
            .I(\tok.A_stk.tail_2 ));
    InMux I__1329 (
            .O(N__11630),
            .I(N__11626));
    CascadeMux I__1328 (
            .O(N__11629),
            .I(N__11623));
    LocalMux I__1327 (
            .O(N__11626),
            .I(N__11620));
    InMux I__1326 (
            .O(N__11623),
            .I(N__11617));
    Span4Mux_h I__1325 (
            .O(N__11620),
            .I(N__11614));
    LocalMux I__1324 (
            .O(N__11617),
            .I(tail_110));
    Odrv4 I__1323 (
            .O(N__11614),
            .I(tail_110));
    CascadeMux I__1322 (
            .O(N__11609),
            .I(N__11605));
    CascadeMux I__1321 (
            .O(N__11608),
            .I(N__11602));
    InMux I__1320 (
            .O(N__11605),
            .I(N__11599));
    InMux I__1319 (
            .O(N__11602),
            .I(N__11596));
    LocalMux I__1318 (
            .O(N__11599),
            .I(N__11593));
    LocalMux I__1317 (
            .O(N__11596),
            .I(N__11590));
    Odrv4 I__1316 (
            .O(N__11593),
            .I(tail_126));
    Odrv4 I__1315 (
            .O(N__11590),
            .I(tail_126));
    InMux I__1314 (
            .O(N__11585),
            .I(N__11582));
    LocalMux I__1313 (
            .O(N__11582),
            .I(\tok.n4 ));
    CascadeMux I__1312 (
            .O(N__11579),
            .I(\tok.n206_cascade_ ));
    CascadeMux I__1311 (
            .O(N__11576),
            .I(\tok.n204_cascade_ ));
    CascadeMux I__1310 (
            .O(N__11573),
            .I(\tok.n16_adj_699_cascade_ ));
    CascadeMux I__1309 (
            .O(N__11570),
            .I(N__11567));
    InMux I__1308 (
            .O(N__11567),
            .I(N__11564));
    LocalMux I__1307 (
            .O(N__11564),
            .I(\tok.n4667 ));
    InMux I__1306 (
            .O(N__11561),
            .I(N__11556));
    InMux I__1305 (
            .O(N__11560),
            .I(N__11553));
    InMux I__1304 (
            .O(N__11559),
            .I(N__11550));
    LocalMux I__1303 (
            .O(N__11556),
            .I(N__11547));
    LocalMux I__1302 (
            .O(N__11553),
            .I(capture_9));
    LocalMux I__1301 (
            .O(N__11550),
            .I(capture_9));
    Odrv4 I__1300 (
            .O(N__11547),
            .I(capture_9));
    CascadeMux I__1299 (
            .O(N__11540),
            .I(\tok.n4508_cascade_ ));
    InMux I__1298 (
            .O(N__11537),
            .I(N__11534));
    LocalMux I__1297 (
            .O(N__11534),
            .I(\tok.n4680 ));
    CascadeMux I__1296 (
            .O(N__11531),
            .I(\tok.n16_adj_660_cascade_ ));
    CascadeMux I__1295 (
            .O(N__11528),
            .I(\tok.uart.n3994_cascade_ ));
    InMux I__1294 (
            .O(N__11525),
            .I(N__11522));
    LocalMux I__1293 (
            .O(N__11522),
            .I(N__11518));
    InMux I__1292 (
            .O(N__11521),
            .I(N__11515));
    Odrv4 I__1291 (
            .O(N__11518),
            .I(n795));
    LocalMux I__1290 (
            .O(N__11515),
            .I(n795));
    CascadeMux I__1289 (
            .O(N__11510),
            .I(\tok.uart.n4506_cascade_ ));
    SRMux I__1288 (
            .O(N__11507),
            .I(N__11504));
    LocalMux I__1287 (
            .O(N__11504),
            .I(N__11501));
    Span4Mux_s2_h I__1286 (
            .O(N__11501),
            .I(N__11498));
    Odrv4 I__1285 (
            .O(N__11498),
            .I(\tok.uart.rxclkcounter_6__N_477 ));
    InMux I__1284 (
            .O(N__11495),
            .I(N__11492));
    LocalMux I__1283 (
            .O(N__11492),
            .I(\tok.uart.n4438 ));
    InMux I__1282 (
            .O(N__11489),
            .I(N__11483));
    InMux I__1281 (
            .O(N__11488),
            .I(N__11483));
    LocalMux I__1280 (
            .O(N__11483),
            .I(\tok.uart.n2 ));
    InMux I__1279 (
            .O(N__11480),
            .I(N__11477));
    LocalMux I__1278 (
            .O(N__11477),
            .I(N__11474));
    Odrv4 I__1277 (
            .O(N__11474),
            .I(\tok.n16_adj_769 ));
    InMux I__1276 (
            .O(N__11471),
            .I(N__11465));
    InMux I__1275 (
            .O(N__11470),
            .I(N__11462));
    InMux I__1274 (
            .O(N__11469),
            .I(N__11457));
    InMux I__1273 (
            .O(N__11468),
            .I(N__11457));
    LocalMux I__1272 (
            .O(N__11465),
            .I(\tok.uart.bytephase_1 ));
    LocalMux I__1271 (
            .O(N__11462),
            .I(\tok.uart.bytephase_1 ));
    LocalMux I__1270 (
            .O(N__11457),
            .I(\tok.uart.bytephase_1 ));
    CascadeMux I__1269 (
            .O(N__11450),
            .I(N__11444));
    CascadeMux I__1268 (
            .O(N__11449),
            .I(N__11441));
    InMux I__1267 (
            .O(N__11448),
            .I(N__11438));
    InMux I__1266 (
            .O(N__11447),
            .I(N__11435));
    InMux I__1265 (
            .O(N__11444),
            .I(N__11430));
    InMux I__1264 (
            .O(N__11441),
            .I(N__11430));
    LocalMux I__1263 (
            .O(N__11438),
            .I(\tok.uart.bytephase_5 ));
    LocalMux I__1262 (
            .O(N__11435),
            .I(\tok.uart.bytephase_5 ));
    LocalMux I__1261 (
            .O(N__11430),
            .I(\tok.uart.bytephase_5 ));
    InMux I__1260 (
            .O(N__11423),
            .I(N__11417));
    InMux I__1259 (
            .O(N__11422),
            .I(N__11414));
    InMux I__1258 (
            .O(N__11421),
            .I(N__11409));
    InMux I__1257 (
            .O(N__11420),
            .I(N__11409));
    LocalMux I__1256 (
            .O(N__11417),
            .I(\tok.uart.bytephase_3 ));
    LocalMux I__1255 (
            .O(N__11414),
            .I(\tok.uart.bytephase_3 ));
    LocalMux I__1254 (
            .O(N__11409),
            .I(\tok.uart.bytephase_3 ));
    InMux I__1253 (
            .O(N__11402),
            .I(N__11396));
    InMux I__1252 (
            .O(N__11401),
            .I(N__11393));
    InMux I__1251 (
            .O(N__11400),
            .I(N__11388));
    InMux I__1250 (
            .O(N__11399),
            .I(N__11388));
    LocalMux I__1249 (
            .O(N__11396),
            .I(\tok.uart.bytephase_0 ));
    LocalMux I__1248 (
            .O(N__11393),
            .I(\tok.uart.bytephase_0 ));
    LocalMux I__1247 (
            .O(N__11388),
            .I(\tok.uart.bytephase_0 ));
    InMux I__1246 (
            .O(N__11381),
            .I(N__11376));
    InMux I__1245 (
            .O(N__11380),
            .I(N__11373));
    InMux I__1244 (
            .O(N__11379),
            .I(N__11370));
    LocalMux I__1243 (
            .O(N__11376),
            .I(\tok.uart.bytephase_2 ));
    LocalMux I__1242 (
            .O(N__11373),
            .I(\tok.uart.bytephase_2 ));
    LocalMux I__1241 (
            .O(N__11370),
            .I(\tok.uart.bytephase_2 ));
    CascadeMux I__1240 (
            .O(N__11363),
            .I(\tok.uart.n13_cascade_ ));
    InMux I__1239 (
            .O(N__11360),
            .I(N__11354));
    InMux I__1238 (
            .O(N__11359),
            .I(N__11351));
    InMux I__1237 (
            .O(N__11358),
            .I(N__11346));
    InMux I__1236 (
            .O(N__11357),
            .I(N__11346));
    LocalMux I__1235 (
            .O(N__11354),
            .I(\tok.uart.bytephase_4 ));
    LocalMux I__1234 (
            .O(N__11351),
            .I(\tok.uart.bytephase_4 ));
    LocalMux I__1233 (
            .O(N__11346),
            .I(\tok.uart.bytephase_4 ));
    SRMux I__1232 (
            .O(N__11339),
            .I(N__11336));
    LocalMux I__1231 (
            .O(N__11336),
            .I(N__11332));
    InMux I__1230 (
            .O(N__11335),
            .I(N__11329));
    Odrv12 I__1229 (
            .O(N__11332),
            .I(bytephase_5__N_510));
    LocalMux I__1228 (
            .O(N__11329),
            .I(bytephase_5__N_510));
    InMux I__1227 (
            .O(N__11324),
            .I(N__11320));
    CascadeMux I__1226 (
            .O(N__11323),
            .I(N__11317));
    LocalMux I__1225 (
            .O(N__11320),
            .I(N__11313));
    InMux I__1224 (
            .O(N__11317),
            .I(N__11308));
    InMux I__1223 (
            .O(N__11316),
            .I(N__11308));
    Span4Mux_s3_h I__1222 (
            .O(N__11313),
            .I(N__11303));
    LocalMux I__1221 (
            .O(N__11308),
            .I(N__11303));
    Span4Mux_v I__1220 (
            .O(N__11303),
            .I(N__11300));
    IoSpan4Mux I__1219 (
            .O(N__11300),
            .I(N__11297));
    Odrv4 I__1218 (
            .O(N__11297),
            .I(rx_c));
    CascadeMux I__1217 (
            .O(N__11294),
            .I(\tok.n18_adj_767_cascade_ ));
    CascadeMux I__1216 (
            .O(N__11291),
            .I(\tok.n20_adj_770_cascade_ ));
    CascadeMux I__1215 (
            .O(N__11288),
            .I(\tok.A_15_N_113_7_cascade_ ));
    InMux I__1214 (
            .O(N__11285),
            .I(N__11282));
    LocalMux I__1213 (
            .O(N__11282),
            .I(\tok.A_15_N_84_7 ));
    InMux I__1212 (
            .O(N__11279),
            .I(N__11276));
    LocalMux I__1211 (
            .O(N__11276),
            .I(\tok.A_15_N_113_7 ));
    InMux I__1210 (
            .O(N__11273),
            .I(N__11267));
    InMux I__1209 (
            .O(N__11272),
            .I(N__11267));
    LocalMux I__1208 (
            .O(N__11267),
            .I(\tok.uart.sentbits_3 ));
    CascadeMux I__1207 (
            .O(N__11264),
            .I(N__11259));
    InMux I__1206 (
            .O(N__11263),
            .I(N__11252));
    InMux I__1205 (
            .O(N__11262),
            .I(N__11252));
    InMux I__1204 (
            .O(N__11259),
            .I(N__11252));
    LocalMux I__1203 (
            .O(N__11252),
            .I(\tok.uart.sentbits_2 ));
    InMux I__1202 (
            .O(N__11249),
            .I(N__11245));
    CascadeMux I__1201 (
            .O(N__11248),
            .I(N__11242));
    LocalMux I__1200 (
            .O(N__11245),
            .I(N__11239));
    InMux I__1199 (
            .O(N__11242),
            .I(N__11236));
    Odrv4 I__1198 (
            .O(N__11239),
            .I(tail_106));
    LocalMux I__1197 (
            .O(N__11236),
            .I(tail_106));
    CascadeMux I__1196 (
            .O(N__11231),
            .I(N__11228));
    InMux I__1195 (
            .O(N__11228),
            .I(N__11222));
    InMux I__1194 (
            .O(N__11227),
            .I(N__11222));
    LocalMux I__1193 (
            .O(N__11222),
            .I(\tok.A_stk.tail_90 ));
    InMux I__1192 (
            .O(N__11219),
            .I(N__11213));
    InMux I__1191 (
            .O(N__11218),
            .I(N__11213));
    LocalMux I__1190 (
            .O(N__11213),
            .I(\tok.A_stk.tail_74 ));
    InMux I__1189 (
            .O(N__11210),
            .I(N__11204));
    InMux I__1188 (
            .O(N__11209),
            .I(N__11204));
    LocalMux I__1187 (
            .O(N__11204),
            .I(\tok.A_stk.tail_58 ));
    CascadeMux I__1186 (
            .O(N__11201),
            .I(N__11197));
    CascadeMux I__1185 (
            .O(N__11200),
            .I(N__11194));
    InMux I__1184 (
            .O(N__11197),
            .I(N__11189));
    InMux I__1183 (
            .O(N__11194),
            .I(N__11189));
    LocalMux I__1182 (
            .O(N__11189),
            .I(\tok.A_stk.tail_42 ));
    CascadeMux I__1181 (
            .O(N__11186),
            .I(N__11182));
    InMux I__1180 (
            .O(N__11185),
            .I(N__11177));
    InMux I__1179 (
            .O(N__11182),
            .I(N__11177));
    LocalMux I__1178 (
            .O(N__11177),
            .I(\tok.A_stk.tail_26 ));
    InMux I__1177 (
            .O(N__11174),
            .I(N__11168));
    InMux I__1176 (
            .O(N__11173),
            .I(N__11168));
    LocalMux I__1175 (
            .O(N__11168),
            .I(\tok.A_stk.tail_10 ));
    InMux I__1174 (
            .O(N__11165),
            .I(N__11162));
    LocalMux I__1173 (
            .O(N__11162),
            .I(\tok.n2_adj_763 ));
    CascadeMux I__1172 (
            .O(N__11159),
            .I(\tok.n13_adj_765_cascade_ ));
    InMux I__1171 (
            .O(N__11156),
            .I(N__11152));
    InMux I__1170 (
            .O(N__11155),
            .I(N__11149));
    LocalMux I__1169 (
            .O(N__11152),
            .I(\tok.A_stk.tail_8 ));
    LocalMux I__1168 (
            .O(N__11149),
            .I(\tok.A_stk.tail_8 ));
    InMux I__1167 (
            .O(N__11144),
            .I(N__11140));
    CascadeMux I__1166 (
            .O(N__11143),
            .I(N__11137));
    LocalMux I__1165 (
            .O(N__11140),
            .I(N__11134));
    InMux I__1164 (
            .O(N__11137),
            .I(N__11131));
    Odrv4 I__1163 (
            .O(N__11134),
            .I(tail_96));
    LocalMux I__1162 (
            .O(N__11131),
            .I(tail_96));
    CascadeMux I__1161 (
            .O(N__11126),
            .I(N__11123));
    InMux I__1160 (
            .O(N__11123),
            .I(N__11119));
    InMux I__1159 (
            .O(N__11122),
            .I(N__11116));
    LocalMux I__1158 (
            .O(N__11119),
            .I(N__11113));
    LocalMux I__1157 (
            .O(N__11116),
            .I(tail_112));
    Odrv4 I__1156 (
            .O(N__11113),
            .I(tail_112));
    InMux I__1155 (
            .O(N__11108),
            .I(N__11105));
    LocalMux I__1154 (
            .O(N__11105),
            .I(N__11101));
    InMux I__1153 (
            .O(N__11104),
            .I(N__11098));
    Odrv4 I__1152 (
            .O(N__11101),
            .I(tail_105));
    LocalMux I__1151 (
            .O(N__11098),
            .I(tail_105));
    CascadeMux I__1150 (
            .O(N__11093),
            .I(N__11090));
    InMux I__1149 (
            .O(N__11090),
            .I(N__11086));
    InMux I__1148 (
            .O(N__11089),
            .I(N__11083));
    LocalMux I__1147 (
            .O(N__11086),
            .I(N__11080));
    LocalMux I__1146 (
            .O(N__11083),
            .I(tail_121));
    Odrv4 I__1145 (
            .O(N__11080),
            .I(tail_121));
    InMux I__1144 (
            .O(N__11075),
            .I(N__11071));
    InMux I__1143 (
            .O(N__11074),
            .I(N__11068));
    LocalMux I__1142 (
            .O(N__11071),
            .I(tail_104));
    LocalMux I__1141 (
            .O(N__11068),
            .I(tail_104));
    CascadeMux I__1140 (
            .O(N__11063),
            .I(N__11060));
    InMux I__1139 (
            .O(N__11060),
            .I(N__11056));
    InMux I__1138 (
            .O(N__11059),
            .I(N__11053));
    LocalMux I__1137 (
            .O(N__11056),
            .I(N__11050));
    LocalMux I__1136 (
            .O(N__11053),
            .I(tail_120));
    Odrv4 I__1135 (
            .O(N__11050),
            .I(tail_120));
    CascadeMux I__1134 (
            .O(N__11045),
            .I(N__11042));
    InMux I__1133 (
            .O(N__11042),
            .I(N__11039));
    LocalMux I__1132 (
            .O(N__11039),
            .I(N__11035));
    CascadeMux I__1131 (
            .O(N__11038),
            .I(N__11032));
    Span4Mux_v I__1130 (
            .O(N__11035),
            .I(N__11029));
    InMux I__1129 (
            .O(N__11032),
            .I(N__11026));
    Odrv4 I__1128 (
            .O(N__11029),
            .I(tail_103));
    LocalMux I__1127 (
            .O(N__11026),
            .I(tail_103));
    CascadeMux I__1126 (
            .O(N__11021),
            .I(N__11018));
    InMux I__1125 (
            .O(N__11018),
            .I(N__11015));
    LocalMux I__1124 (
            .O(N__11015),
            .I(N__11011));
    InMux I__1123 (
            .O(N__11014),
            .I(N__11008));
    Span4Mux_v I__1122 (
            .O(N__11011),
            .I(N__11005));
    LocalMux I__1121 (
            .O(N__11008),
            .I(tail_119));
    Odrv4 I__1120 (
            .O(N__11005),
            .I(tail_119));
    InMux I__1119 (
            .O(N__11000),
            .I(N__10997));
    LocalMux I__1118 (
            .O(N__10997),
            .I(N__10994));
    Span4Mux_h I__1117 (
            .O(N__10994),
            .I(N__10991));
    Odrv4 I__1116 (
            .O(N__10991),
            .I(\tok.table_wr_data_12 ));
    CascadeMux I__1115 (
            .O(N__10988),
            .I(N__10985));
    InMux I__1114 (
            .O(N__10985),
            .I(N__10981));
    InMux I__1113 (
            .O(N__10984),
            .I(N__10978));
    LocalMux I__1112 (
            .O(N__10981),
            .I(N__10975));
    LocalMux I__1111 (
            .O(N__10978),
            .I(tail_122));
    Odrv4 I__1110 (
            .O(N__10975),
            .I(tail_122));
    CascadeMux I__1109 (
            .O(N__10970),
            .I(N__10966));
    CascadeMux I__1108 (
            .O(N__10969),
            .I(N__10963));
    InMux I__1107 (
            .O(N__10966),
            .I(N__10958));
    InMux I__1106 (
            .O(N__10963),
            .I(N__10958));
    LocalMux I__1105 (
            .O(N__10958),
            .I(\tok.A_stk.tail_30 ));
    InMux I__1104 (
            .O(N__10955),
            .I(N__10951));
    InMux I__1103 (
            .O(N__10954),
            .I(N__10948));
    LocalMux I__1102 (
            .O(N__10951),
            .I(\tok.A_stk.tail_14 ));
    LocalMux I__1101 (
            .O(N__10948),
            .I(\tok.A_stk.tail_14 ));
    InMux I__1100 (
            .O(N__10943),
            .I(N__10937));
    InMux I__1099 (
            .O(N__10942),
            .I(N__10937));
    LocalMux I__1098 (
            .O(N__10937),
            .I(\tok.A_stk.tail_88 ));
    InMux I__1097 (
            .O(N__10934),
            .I(N__10928));
    InMux I__1096 (
            .O(N__10933),
            .I(N__10928));
    LocalMux I__1095 (
            .O(N__10928),
            .I(\tok.A_stk.tail_72 ));
    CascadeMux I__1094 (
            .O(N__10925),
            .I(N__10921));
    CascadeMux I__1093 (
            .O(N__10924),
            .I(N__10918));
    InMux I__1092 (
            .O(N__10921),
            .I(N__10913));
    InMux I__1091 (
            .O(N__10918),
            .I(N__10913));
    LocalMux I__1090 (
            .O(N__10913),
            .I(N__10910));
    Odrv4 I__1089 (
            .O(N__10910),
            .I(\tok.A_stk.tail_56 ));
    InMux I__1088 (
            .O(N__10907),
            .I(N__10901));
    InMux I__1087 (
            .O(N__10906),
            .I(N__10901));
    LocalMux I__1086 (
            .O(N__10901),
            .I(\tok.A_stk.tail_40 ));
    InMux I__1085 (
            .O(N__10898),
            .I(N__10892));
    InMux I__1084 (
            .O(N__10897),
            .I(N__10892));
    LocalMux I__1083 (
            .O(N__10892),
            .I(\tok.A_stk.tail_24 ));
    InMux I__1082 (
            .O(N__10889),
            .I(N__10883));
    InMux I__1081 (
            .O(N__10888),
            .I(N__10883));
    LocalMux I__1080 (
            .O(N__10883),
            .I(\tok.A_stk.tail_64 ));
    InMux I__1079 (
            .O(N__10880),
            .I(N__10874));
    InMux I__1078 (
            .O(N__10879),
            .I(N__10874));
    LocalMux I__1077 (
            .O(N__10874),
            .I(\tok.A_stk.tail_80 ));
    CascadeMux I__1076 (
            .O(N__10871),
            .I(N__10868));
    InMux I__1075 (
            .O(N__10868),
            .I(N__10864));
    InMux I__1074 (
            .O(N__10867),
            .I(N__10861));
    LocalMux I__1073 (
            .O(N__10864),
            .I(\tok.A_stk.tail_0 ));
    LocalMux I__1072 (
            .O(N__10861),
            .I(\tok.A_stk.tail_0 ));
    CascadeMux I__1071 (
            .O(N__10856),
            .I(N__10853));
    InMux I__1070 (
            .O(N__10853),
            .I(N__10847));
    InMux I__1069 (
            .O(N__10852),
            .I(N__10847));
    LocalMux I__1068 (
            .O(N__10847),
            .I(N__10844));
    Odrv4 I__1067 (
            .O(N__10844),
            .I(\tok.A_stk.tail_94 ));
    InMux I__1066 (
            .O(N__10841),
            .I(N__10835));
    InMux I__1065 (
            .O(N__10840),
            .I(N__10835));
    LocalMux I__1064 (
            .O(N__10835),
            .I(\tok.A_stk.tail_78 ));
    InMux I__1063 (
            .O(N__10832),
            .I(N__10826));
    InMux I__1062 (
            .O(N__10831),
            .I(N__10826));
    LocalMux I__1061 (
            .O(N__10826),
            .I(\tok.A_stk.tail_62 ));
    CascadeMux I__1060 (
            .O(N__10823),
            .I(N__10819));
    CascadeMux I__1059 (
            .O(N__10822),
            .I(N__10816));
    InMux I__1058 (
            .O(N__10819),
            .I(N__10811));
    InMux I__1057 (
            .O(N__10816),
            .I(N__10811));
    LocalMux I__1056 (
            .O(N__10811),
            .I(\tok.A_stk.tail_46 ));
    InMux I__1055 (
            .O(N__10808),
            .I(\tok.uart.n3963 ));
    InMux I__1054 (
            .O(N__10805),
            .I(\tok.uart.n3964 ));
    InMux I__1053 (
            .O(N__10802),
            .I(\tok.uart.n3965 ));
    InMux I__1052 (
            .O(N__10799),
            .I(\tok.uart.n3966 ));
    InMux I__1051 (
            .O(N__10796),
            .I(\tok.uart.n3967 ));
    CEMux I__1050 (
            .O(N__10793),
            .I(N__10790));
    LocalMux I__1049 (
            .O(N__10790),
            .I(N__10787));
    Span4Mux_v I__1048 (
            .O(N__10787),
            .I(N__10784));
    Odrv4 I__1047 (
            .O(N__10784),
            .I(n940));
    CascadeMux I__1046 (
            .O(N__10781),
            .I(N__10778));
    InMux I__1045 (
            .O(N__10778),
            .I(N__10772));
    InMux I__1044 (
            .O(N__10777),
            .I(N__10772));
    LocalMux I__1043 (
            .O(N__10772),
            .I(\tok.A_stk.tail_16 ));
    CascadeMux I__1042 (
            .O(N__10769),
            .I(N__10765));
    InMux I__1041 (
            .O(N__10768),
            .I(N__10762));
    InMux I__1040 (
            .O(N__10765),
            .I(N__10759));
    LocalMux I__1039 (
            .O(N__10762),
            .I(\tok.A_stk.tail_32 ));
    LocalMux I__1038 (
            .O(N__10759),
            .I(\tok.A_stk.tail_32 ));
    CascadeMux I__1037 (
            .O(N__10754),
            .I(N__10750));
    CascadeMux I__1036 (
            .O(N__10753),
            .I(N__10747));
    InMux I__1035 (
            .O(N__10750),
            .I(N__10742));
    InMux I__1034 (
            .O(N__10747),
            .I(N__10742));
    LocalMux I__1033 (
            .O(N__10742),
            .I(\tok.A_stk.tail_48 ));
    InMux I__1032 (
            .O(N__10739),
            .I(N__10736));
    LocalMux I__1031 (
            .O(N__10736),
            .I(N__10733));
    Odrv4 I__1030 (
            .O(N__10733),
            .I(\tok.table_wr_data_8 ));
    InMux I__1029 (
            .O(N__10730),
            .I(N__10727));
    LocalMux I__1028 (
            .O(N__10727),
            .I(N__10724));
    Span4Mux_v I__1027 (
            .O(N__10724),
            .I(N__10721));
    Odrv4 I__1026 (
            .O(N__10721),
            .I(\tok.table_wr_data_15 ));
    InMux I__1025 (
            .O(N__10718),
            .I(N__10715));
    LocalMux I__1024 (
            .O(N__10715),
            .I(N__10712));
    Span4Mux_h I__1023 (
            .O(N__10712),
            .I(N__10709));
    Span4Mux_s1_h I__1022 (
            .O(N__10709),
            .I(N__10706));
    Odrv4 I__1021 (
            .O(N__10706),
            .I(\tok.table_wr_data_14 ));
    InMux I__1020 (
            .O(N__10703),
            .I(N__10700));
    LocalMux I__1019 (
            .O(N__10700),
            .I(N__10697));
    Odrv4 I__1018 (
            .O(N__10697),
            .I(\tok.table_wr_data_13 ));
    InMux I__1017 (
            .O(N__10694),
            .I(N__10691));
    LocalMux I__1016 (
            .O(N__10691),
            .I(N__10688));
    Odrv4 I__1015 (
            .O(N__10688),
            .I(\tok.uart.n12 ));
    InMux I__1014 (
            .O(N__10685),
            .I(N__10681));
    InMux I__1013 (
            .O(N__10684),
            .I(N__10678));
    LocalMux I__1012 (
            .O(N__10681),
            .I(\tok.uart.rxclkcounter_6 ));
    LocalMux I__1011 (
            .O(N__10678),
            .I(\tok.uart.rxclkcounter_6 ));
    CascadeMux I__1010 (
            .O(N__10673),
            .I(N__10669));
    InMux I__1009 (
            .O(N__10672),
            .I(N__10666));
    InMux I__1008 (
            .O(N__10669),
            .I(N__10663));
    LocalMux I__1007 (
            .O(N__10666),
            .I(\tok.uart.rxclkcounter_5 ));
    LocalMux I__1006 (
            .O(N__10663),
            .I(\tok.uart.rxclkcounter_5 ));
    InMux I__1005 (
            .O(N__10658),
            .I(N__10654));
    InMux I__1004 (
            .O(N__10657),
            .I(N__10651));
    LocalMux I__1003 (
            .O(N__10654),
            .I(\tok.uart.rxclkcounter_2 ));
    LocalMux I__1002 (
            .O(N__10651),
            .I(\tok.uart.rxclkcounter_2 ));
    CascadeMux I__1001 (
            .O(N__10646),
            .I(n795_cascade_));
    InMux I__1000 (
            .O(N__10643),
            .I(N__10640));
    LocalMux I__999 (
            .O(N__10640),
            .I(N__10637));
    Span4Mux_h I__998 (
            .O(N__10637),
            .I(N__10634));
    Odrv4 I__997 (
            .O(N__10634),
            .I(\tok.table_wr_data_9 ));
    InMux I__996 (
            .O(N__10631),
            .I(bfn_1_10_0_));
    SRMux I__995 (
            .O(N__10628),
            .I(N__10625));
    LocalMux I__994 (
            .O(N__10625),
            .I(N__10622));
    Span4Mux_h I__993 (
            .O(N__10622),
            .I(N__10619));
    Span4Mux_s0_h I__992 (
            .O(N__10619),
            .I(N__10616));
    Odrv4 I__991 (
            .O(N__10616),
            .I(\tok.uart.n1081 ));
    InMux I__990 (
            .O(N__10613),
            .I(N__10609));
    InMux I__989 (
            .O(N__10612),
            .I(N__10606));
    LocalMux I__988 (
            .O(N__10609),
            .I(\tok.uart.rxclkcounter_0 ));
    LocalMux I__987 (
            .O(N__10606),
            .I(\tok.uart.rxclkcounter_0 ));
    InMux I__986 (
            .O(N__10601),
            .I(bfn_1_8_0_));
    CascadeMux I__985 (
            .O(N__10598),
            .I(N__10595));
    InMux I__984 (
            .O(N__10595),
            .I(N__10591));
    InMux I__983 (
            .O(N__10594),
            .I(N__10588));
    LocalMux I__982 (
            .O(N__10591),
            .I(N__10585));
    LocalMux I__981 (
            .O(N__10588),
            .I(\tok.uart.rxclkcounter_1 ));
    Odrv4 I__980 (
            .O(N__10585),
            .I(\tok.uart.rxclkcounter_1 ));
    InMux I__979 (
            .O(N__10580),
            .I(\tok.uart.n3968 ));
    InMux I__978 (
            .O(N__10577),
            .I(\tok.uart.n3969 ));
    InMux I__977 (
            .O(N__10574),
            .I(N__10570));
    InMux I__976 (
            .O(N__10573),
            .I(N__10567));
    LocalMux I__975 (
            .O(N__10570),
            .I(\tok.uart.rxclkcounter_3 ));
    LocalMux I__974 (
            .O(N__10567),
            .I(\tok.uart.rxclkcounter_3 ));
    InMux I__973 (
            .O(N__10562),
            .I(\tok.uart.n3970 ));
    InMux I__972 (
            .O(N__10559),
            .I(N__10555));
    InMux I__971 (
            .O(N__10558),
            .I(N__10552));
    LocalMux I__970 (
            .O(N__10555),
            .I(\tok.uart.rxclkcounter_4 ));
    LocalMux I__969 (
            .O(N__10552),
            .I(\tok.uart.rxclkcounter_4 ));
    InMux I__968 (
            .O(N__10547),
            .I(\tok.uart.n3971 ));
    InMux I__967 (
            .O(N__10544),
            .I(\tok.uart.n3972 ));
    InMux I__966 (
            .O(N__10541),
            .I(\tok.uart.n3973 ));
    InMux I__965 (
            .O(N__10538),
            .I(\tok.uart.n3960 ));
    InMux I__964 (
            .O(N__10535),
            .I(\tok.uart.n3961 ));
    InMux I__963 (
            .O(N__10532),
            .I(bfn_1_6_0_));
    InMux I__962 (
            .O(N__10529),
            .I(N__10525));
    InMux I__961 (
            .O(N__10528),
            .I(N__10522));
    LocalMux I__960 (
            .O(N__10525),
            .I(N__10519));
    LocalMux I__959 (
            .O(N__10522),
            .I(\tok.uart.txclkcounter_3 ));
    Odrv4 I__958 (
            .O(N__10519),
            .I(\tok.uart.txclkcounter_3 ));
    InMux I__957 (
            .O(N__10514),
            .I(N__10510));
    InMux I__956 (
            .O(N__10513),
            .I(N__10507));
    LocalMux I__955 (
            .O(N__10510),
            .I(N__10504));
    LocalMux I__954 (
            .O(N__10507),
            .I(\tok.uart.txclkcounter_5 ));
    Odrv4 I__953 (
            .O(N__10504),
            .I(\tok.uart.txclkcounter_5 ));
    CascadeMux I__952 (
            .O(N__10499),
            .I(N__10496));
    InMux I__951 (
            .O(N__10496),
            .I(N__10492));
    InMux I__950 (
            .O(N__10495),
            .I(N__10489));
    LocalMux I__949 (
            .O(N__10492),
            .I(N__10486));
    LocalMux I__948 (
            .O(N__10489),
            .I(\tok.uart.txclkcounter_0 ));
    Odrv12 I__947 (
            .O(N__10486),
            .I(\tok.uart.txclkcounter_0 ));
    InMux I__946 (
            .O(N__10481),
            .I(N__10477));
    InMux I__945 (
            .O(N__10480),
            .I(N__10474));
    LocalMux I__944 (
            .O(N__10477),
            .I(N__10471));
    LocalMux I__943 (
            .O(N__10474),
            .I(\tok.uart.txclkcounter_2 ));
    Odrv4 I__942 (
            .O(N__10471),
            .I(\tok.uart.txclkcounter_2 ));
    InMux I__941 (
            .O(N__10466),
            .I(N__10462));
    InMux I__940 (
            .O(N__10465),
            .I(N__10459));
    LocalMux I__939 (
            .O(N__10462),
            .I(N__10456));
    LocalMux I__938 (
            .O(N__10459),
            .I(\tok.uart.txclkcounter_6 ));
    Odrv4 I__937 (
            .O(N__10456),
            .I(\tok.uart.txclkcounter_6 ));
    InMux I__936 (
            .O(N__10451),
            .I(N__10447));
    InMux I__935 (
            .O(N__10450),
            .I(N__10444));
    LocalMux I__934 (
            .O(N__10447),
            .I(N__10441));
    LocalMux I__933 (
            .O(N__10444),
            .I(\tok.uart.txclkcounter_1 ));
    Odrv12 I__932 (
            .O(N__10441),
            .I(\tok.uart.txclkcounter_1 ));
    InMux I__931 (
            .O(N__10436),
            .I(N__10432));
    InMux I__930 (
            .O(N__10435),
            .I(N__10429));
    LocalMux I__929 (
            .O(N__10432),
            .I(N__10426));
    LocalMux I__928 (
            .O(N__10429),
            .I(\tok.uart.txclkcounter_7 ));
    Odrv4 I__927 (
            .O(N__10426),
            .I(\tok.uart.txclkcounter_7 ));
    InMux I__926 (
            .O(N__10421),
            .I(N__10417));
    InMux I__925 (
            .O(N__10420),
            .I(N__10414));
    LocalMux I__924 (
            .O(N__10417),
            .I(N__10411));
    LocalMux I__923 (
            .O(N__10414),
            .I(\tok.uart.txclkcounter_8 ));
    Odrv4 I__922 (
            .O(N__10411),
            .I(\tok.uart.txclkcounter_8 ));
    InMux I__921 (
            .O(N__10406),
            .I(N__10402));
    InMux I__920 (
            .O(N__10405),
            .I(N__10399));
    LocalMux I__919 (
            .O(N__10402),
            .I(N__10396));
    LocalMux I__918 (
            .O(N__10399),
            .I(\tok.uart.txclkcounter_4 ));
    Odrv4 I__917 (
            .O(N__10396),
            .I(\tok.uart.txclkcounter_4 ));
    CascadeMux I__916 (
            .O(N__10391),
            .I(\tok.uart.n14_cascade_ ));
    InMux I__915 (
            .O(N__10388),
            .I(N__10385));
    LocalMux I__914 (
            .O(N__10385),
            .I(\tok.uart.n15_adj_640 ));
    CascadeMux I__913 (
            .O(N__10382),
            .I(txtick_cascade_));
    InMux I__912 (
            .O(N__10379),
            .I(N__10373));
    InMux I__911 (
            .O(N__10378),
            .I(N__10373));
    LocalMux I__910 (
            .O(N__10373),
            .I(\tok.A_stk.tail_43 ));
    CascadeMux I__909 (
            .O(N__10370),
            .I(N__10366));
    InMux I__908 (
            .O(N__10369),
            .I(N__10361));
    InMux I__907 (
            .O(N__10366),
            .I(N__10361));
    LocalMux I__906 (
            .O(N__10361),
            .I(\tok.A_stk.tail_27 ));
    InMux I__905 (
            .O(N__10358),
            .I(N__10354));
    InMux I__904 (
            .O(N__10357),
            .I(N__10351));
    LocalMux I__903 (
            .O(N__10354),
            .I(\tok.A_stk.tail_11 ));
    LocalMux I__902 (
            .O(N__10351),
            .I(\tok.A_stk.tail_11 ));
    InMux I__901 (
            .O(N__10346),
            .I(bfn_1_5_0_));
    InMux I__900 (
            .O(N__10343),
            .I(\tok.uart.n3955 ));
    InMux I__899 (
            .O(N__10340),
            .I(\tok.uart.n3956 ));
    InMux I__898 (
            .O(N__10337),
            .I(\tok.uart.n3957 ));
    InMux I__897 (
            .O(N__10334),
            .I(\tok.uart.n3958 ));
    InMux I__896 (
            .O(N__10331),
            .I(\tok.uart.n3959 ));
    CascadeMux I__895 (
            .O(N__10328),
            .I(N__10324));
    InMux I__894 (
            .O(N__10327),
            .I(N__10321));
    InMux I__893 (
            .O(N__10324),
            .I(N__10318));
    LocalMux I__892 (
            .O(N__10321),
            .I(\tok.A_stk.tail_39 ));
    LocalMux I__891 (
            .O(N__10318),
            .I(\tok.A_stk.tail_39 ));
    CascadeMux I__890 (
            .O(N__10313),
            .I(N__10309));
    CascadeMux I__889 (
            .O(N__10312),
            .I(N__10306));
    InMux I__888 (
            .O(N__10309),
            .I(N__10301));
    InMux I__887 (
            .O(N__10306),
            .I(N__10301));
    LocalMux I__886 (
            .O(N__10301),
            .I(\tok.A_stk.tail_23 ));
    CascadeMux I__885 (
            .O(N__10298),
            .I(N__10295));
    InMux I__884 (
            .O(N__10295),
            .I(N__10289));
    InMux I__883 (
            .O(N__10294),
            .I(N__10289));
    LocalMux I__882 (
            .O(N__10289),
            .I(\tok.A_stk.tail_7 ));
    CascadeMux I__881 (
            .O(N__10286),
            .I(N__10282));
    CascadeMux I__880 (
            .O(N__10285),
            .I(N__10279));
    InMux I__879 (
            .O(N__10282),
            .I(N__10276));
    InMux I__878 (
            .O(N__10279),
            .I(N__10273));
    LocalMux I__877 (
            .O(N__10276),
            .I(tail_123));
    LocalMux I__876 (
            .O(N__10273),
            .I(tail_123));
    InMux I__875 (
            .O(N__10268),
            .I(N__10264));
    InMux I__874 (
            .O(N__10267),
            .I(N__10261));
    LocalMux I__873 (
            .O(N__10264),
            .I(tail_107));
    LocalMux I__872 (
            .O(N__10261),
            .I(tail_107));
    CascadeMux I__871 (
            .O(N__10256),
            .I(N__10253));
    InMux I__870 (
            .O(N__10253),
            .I(N__10247));
    InMux I__869 (
            .O(N__10252),
            .I(N__10247));
    LocalMux I__868 (
            .O(N__10247),
            .I(\tok.A_stk.tail_91 ));
    InMux I__867 (
            .O(N__10244),
            .I(N__10238));
    InMux I__866 (
            .O(N__10243),
            .I(N__10238));
    LocalMux I__865 (
            .O(N__10238),
            .I(\tok.A_stk.tail_75 ));
    InMux I__864 (
            .O(N__10235),
            .I(N__10229));
    InMux I__863 (
            .O(N__10234),
            .I(N__10229));
    LocalMux I__862 (
            .O(N__10229),
            .I(\tok.A_stk.tail_59 ));
    InMux I__861 (
            .O(N__10226),
            .I(N__10220));
    InMux I__860 (
            .O(N__10225),
            .I(N__10220));
    LocalMux I__859 (
            .O(N__10220),
            .I(\tok.A_stk.tail_73 ));
    CascadeMux I__858 (
            .O(N__10217),
            .I(N__10213));
    CascadeMux I__857 (
            .O(N__10216),
            .I(N__10210));
    InMux I__856 (
            .O(N__10213),
            .I(N__10205));
    InMux I__855 (
            .O(N__10210),
            .I(N__10205));
    LocalMux I__854 (
            .O(N__10205),
            .I(N__10202));
    Odrv4 I__853 (
            .O(N__10202),
            .I(\tok.A_stk.tail_57 ));
    InMux I__852 (
            .O(N__10199),
            .I(N__10193));
    InMux I__851 (
            .O(N__10198),
            .I(N__10193));
    LocalMux I__850 (
            .O(N__10193),
            .I(\tok.A_stk.tail_41 ));
    InMux I__849 (
            .O(N__10190),
            .I(N__10184));
    InMux I__848 (
            .O(N__10189),
            .I(N__10184));
    LocalMux I__847 (
            .O(N__10184),
            .I(\tok.A_stk.tail_25 ));
    InMux I__846 (
            .O(N__10181),
            .I(N__10177));
    InMux I__845 (
            .O(N__10180),
            .I(N__10174));
    LocalMux I__844 (
            .O(N__10177),
            .I(\tok.A_stk.tail_9 ));
    LocalMux I__843 (
            .O(N__10174),
            .I(\tok.A_stk.tail_9 ));
    InMux I__842 (
            .O(N__10169),
            .I(N__10163));
    InMux I__841 (
            .O(N__10168),
            .I(N__10163));
    LocalMux I__840 (
            .O(N__10163),
            .I(\tok.A_stk.tail_87 ));
    InMux I__839 (
            .O(N__10160),
            .I(N__10154));
    InMux I__838 (
            .O(N__10159),
            .I(N__10154));
    LocalMux I__837 (
            .O(N__10154),
            .I(\tok.A_stk.tail_71 ));
    CascadeMux I__836 (
            .O(N__10151),
            .I(N__10148));
    InMux I__835 (
            .O(N__10148),
            .I(N__10144));
    InMux I__834 (
            .O(N__10147),
            .I(N__10141));
    LocalMux I__833 (
            .O(N__10144),
            .I(\tok.A_stk.tail_55 ));
    LocalMux I__832 (
            .O(N__10141),
            .I(\tok.A_stk.tail_55 ));
    InMux I__831 (
            .O(N__10136),
            .I(N__10130));
    InMux I__830 (
            .O(N__10135),
            .I(N__10130));
    LocalMux I__829 (
            .O(N__10130),
            .I(\tok.A_stk.tail_89 ));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(\tok.uart.n3962 ),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(\tok.n3917 ),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(\tok.n3924_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(\tok.n3909 ),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(\tok.n3947 ),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\tok.n3932 ),
            .carryinitout(bfn_9_9_0_));
    GND GND (
            .Y(GNDG0));
    defparam OSCInst0.CLKHF_DIV="0b01";
    SB_HFOSC OSCInst0 (
            .CLKHFPU(N__21701),
            .CLKHFEN(N__21700),
            .CLKHF(clk));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i123_LC_0_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i123_LC_0_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i123_LC_0_4_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \tok.A_stk.tail_i0_i123_LC_0_4_1  (
            .in0(N__10268),
            .in1(N__13908),
            .in2(N__10286),
            .in3(N__14468),
            .lcout(tail_123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26195),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i105_LC_0_6_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i105_LC_0_6_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i105_LC_0_6_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i105_LC_0_6_0  (
            .in0(N__10135),
            .in1(N__13892),
            .in2(N__11093),
            .in3(N__14541),
            .lcout(tail_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26199),
            .ce(N__14736),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i89_LC_0_6_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i89_LC_0_6_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i89_LC_0_6_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i89_LC_0_6_1  (
            .in0(N__14539),
            .in1(N__11104),
            .in2(N__13931),
            .in3(N__10225),
            .lcout(\tok.A_stk.tail_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26199),
            .ce(N__14736),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i73_LC_0_6_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i73_LC_0_6_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i73_LC_0_6_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i73_LC_0_6_2  (
            .in0(N__10136),
            .in1(N__13894),
            .in2(N__10216),
            .in3(N__14543),
            .lcout(\tok.A_stk.tail_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26199),
            .ce(N__14736),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i57_LC_0_6_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i57_LC_0_6_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i57_LC_0_6_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i57_LC_0_6_3  (
            .in0(N__14538),
            .in1(N__10198),
            .in2(N__13930),
            .in3(N__10226),
            .lcout(\tok.A_stk.tail_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26199),
            .ce(N__14736),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i41_LC_0_6_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i41_LC_0_6_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i41_LC_0_6_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i41_LC_0_6_4  (
            .in0(N__10189),
            .in1(N__13893),
            .in2(N__10217),
            .in3(N__14542),
            .lcout(\tok.A_stk.tail_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26199),
            .ce(N__14736),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i25_LC_0_6_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i25_LC_0_6_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i25_LC_0_6_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i25_LC_0_6_5  (
            .in0(N__14537),
            .in1(N__10181),
            .in2(N__13929),
            .in3(N__10199),
            .lcout(\tok.A_stk.tail_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26199),
            .ce(N__14736),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i9_LC_0_6_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i9_LC_0_6_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i9_LC_0_6_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i9_LC_0_6_6  (
            .in0(N__10190),
            .in1(N__14540),
            .in2(N__21145),
            .in3(N__13904),
            .lcout(\tok.A_stk.tail_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26199),
            .ce(N__14736),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i9_LC_0_6_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i9_LC_0_6_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i9_LC_0_6_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i9_LC_0_6_7  (
            .in0(N__10180),
            .in1(N__15746),
            .in2(_gnd_net_),
            .in3(N__22651),
            .lcout(\tok.S_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26199),
            .ce(N__14736),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i103_LC_0_7_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i103_LC_0_7_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i103_LC_0_7_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i103_LC_0_7_0  (
            .in0(N__13878),
            .in1(N__10168),
            .in2(N__11021),
            .in3(N__14534),
            .lcout(tail_103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26203),
            .ce(N__14728),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i87_LC_0_7_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i87_LC_0_7_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i87_LC_0_7_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i87_LC_0_7_1  (
            .in0(N__14532),
            .in1(N__10159),
            .in2(N__11038),
            .in3(N__13883),
            .lcout(\tok.A_stk.tail_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26203),
            .ce(N__14728),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i71_LC_0_7_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i71_LC_0_7_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i71_LC_0_7_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i71_LC_0_7_2  (
            .in0(N__13880),
            .in1(N__10169),
            .in2(N__10151),
            .in3(N__14536),
            .lcout(\tok.A_stk.tail_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26203),
            .ce(N__14728),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i55_LC_0_7_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i55_LC_0_7_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i55_LC_0_7_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i55_LC_0_7_3  (
            .in0(N__14531),
            .in1(N__10160),
            .in2(N__10328),
            .in3(N__13882),
            .lcout(\tok.A_stk.tail_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26203),
            .ce(N__14728),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i39_LC_0_7_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i39_LC_0_7_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i39_LC_0_7_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i39_LC_0_7_4  (
            .in0(N__13879),
            .in1(N__10147),
            .in2(N__10312),
            .in3(N__14535),
            .lcout(\tok.A_stk.tail_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26203),
            .ce(N__14728),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i23_LC_0_7_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i23_LC_0_7_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i23_LC_0_7_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i23_LC_0_7_5  (
            .in0(N__14530),
            .in1(N__10327),
            .in2(N__10298),
            .in3(N__13881),
            .lcout(\tok.A_stk.tail_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26203),
            .ce(N__14728),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i7_LC_0_7_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i7_LC_0_7_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i7_LC_0_7_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tok.A_stk.tail_i0_i7_LC_0_7_6  (
            .in0(N__13877),
            .in1(N__14533),
            .in2(N__10313),
            .in3(N__19636),
            .lcout(\tok.A_stk.tail_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26203),
            .ce(N__14728),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i7_LC_0_7_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i7_LC_0_7_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i7_LC_0_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i7_LC_0_7_7  (
            .in0(N__10294),
            .in1(N__15742),
            .in2(_gnd_net_),
            .in3(N__19811),
            .lcout(\tok.S_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26203),
            .ce(N__14728),
            .sr(_gnd_net_));
    defparam \tok.uart.i2_3_lut_LC_0_10_5 .C_ON=1'b0;
    defparam \tok.uart.i2_3_lut_LC_0_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_3_lut_LC_0_10_5 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \tok.uart.i2_3_lut_LC_0_10_5  (
            .in0(N__11521),
            .in1(N__11471),
            .in2(_gnd_net_),
            .in3(N__11401),
            .lcout(n4005),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i107_LC_1_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i107_LC_1_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i107_LC_1_4_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i107_LC_1_4_0  (
            .in0(N__10252),
            .in1(N__13909),
            .in2(N__10285),
            .in3(N__14465),
            .lcout(tail_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26197),
            .ce(N__14729),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i91_LC_1_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i91_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i91_LC_1_4_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i91_LC_1_4_1  (
            .in0(N__14463),
            .in1(N__10267),
            .in2(N__13934),
            .in3(N__10243),
            .lcout(\tok.A_stk.tail_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26197),
            .ce(N__14729),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i75_LC_1_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i75_LC_1_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i75_LC_1_4_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i75_LC_1_4_2  (
            .in0(N__10234),
            .in1(N__13911),
            .in2(N__10256),
            .in3(N__14467),
            .lcout(\tok.A_stk.tail_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26197),
            .ce(N__14729),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i59_LC_1_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i59_LC_1_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i59_LC_1_4_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i59_LC_1_4_3  (
            .in0(N__14462),
            .in1(N__10378),
            .in2(N__13933),
            .in3(N__10244),
            .lcout(\tok.A_stk.tail_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26197),
            .ce(N__14729),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i43_LC_1_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i43_LC_1_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i43_LC_1_4_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i43_LC_1_4_4  (
            .in0(N__10235),
            .in1(N__13910),
            .in2(N__10370),
            .in3(N__14466),
            .lcout(\tok.A_stk.tail_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26197),
            .ce(N__14729),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i27_LC_1_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i27_LC_1_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i27_LC_1_4_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i27_LC_1_4_5  (
            .in0(N__14461),
            .in1(N__10358),
            .in2(N__13932),
            .in3(N__10379),
            .lcout(\tok.A_stk.tail_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26197),
            .ce(N__14729),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i11_LC_1_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i11_LC_1_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i11_LC_1_4_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i11_LC_1_4_6  (
            .in0(N__10369),
            .in1(N__14464),
            .in2(N__20843),
            .in3(N__13921),
            .lcout(\tok.A_stk.tail_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26197),
            .ce(N__14729),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i11_LC_1_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i11_LC_1_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i11_LC_1_4_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i11_LC_1_4_7  (
            .in0(N__10357),
            .in1(N__15744),
            .in2(_gnd_net_),
            .in3(N__21440),
            .lcout(\tok.S_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26197),
            .ce(N__14729),
            .sr(_gnd_net_));
    defparam \tok.uart.txclkcounter_144__i0_LC_1_5_0 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_144__i0_LC_1_5_0 .SEQ_MODE=4'b1001;
    defparam \tok.uart.txclkcounter_144__i0_LC_1_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_144__i0_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(N__10495),
            .in2(_gnd_net_),
            .in3(N__10346),
            .lcout(\tok.uart.txclkcounter_0 ),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(\tok.uart.n3955 ),
            .clk(N__26200),
            .ce(),
            .sr(N__12241));
    defparam \tok.uart.txclkcounter_144__i1_LC_1_5_1 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_144__i1_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_144__i1_LC_1_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_144__i1_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(N__10450),
            .in2(_gnd_net_),
            .in3(N__10343),
            .lcout(\tok.uart.txclkcounter_1 ),
            .ltout(),
            .carryin(\tok.uart.n3955 ),
            .carryout(\tok.uart.n3956 ),
            .clk(N__26200),
            .ce(),
            .sr(N__12241));
    defparam \tok.uart.txclkcounter_144__i2_LC_1_5_2 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_144__i2_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_144__i2_LC_1_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_144__i2_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(N__10480),
            .in2(_gnd_net_),
            .in3(N__10340),
            .lcout(\tok.uart.txclkcounter_2 ),
            .ltout(),
            .carryin(\tok.uart.n3956 ),
            .carryout(\tok.uart.n3957 ),
            .clk(N__26200),
            .ce(),
            .sr(N__12241));
    defparam \tok.uart.txclkcounter_144__i3_LC_1_5_3 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_144__i3_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_144__i3_LC_1_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_144__i3_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(N__10528),
            .in2(_gnd_net_),
            .in3(N__10337),
            .lcout(\tok.uart.txclkcounter_3 ),
            .ltout(),
            .carryin(\tok.uart.n3957 ),
            .carryout(\tok.uart.n3958 ),
            .clk(N__26200),
            .ce(),
            .sr(N__12241));
    defparam \tok.uart.txclkcounter_144__i4_LC_1_5_4 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_144__i4_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_144__i4_LC_1_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_144__i4_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(N__10405),
            .in2(_gnd_net_),
            .in3(N__10334),
            .lcout(\tok.uart.txclkcounter_4 ),
            .ltout(),
            .carryin(\tok.uart.n3958 ),
            .carryout(\tok.uart.n3959 ),
            .clk(N__26200),
            .ce(),
            .sr(N__12241));
    defparam \tok.uart.txclkcounter_144__i5_LC_1_5_5 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_144__i5_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_144__i5_LC_1_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_144__i5_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(N__10513),
            .in2(_gnd_net_),
            .in3(N__10331),
            .lcout(\tok.uart.txclkcounter_5 ),
            .ltout(),
            .carryin(\tok.uart.n3959 ),
            .carryout(\tok.uart.n3960 ),
            .clk(N__26200),
            .ce(),
            .sr(N__12241));
    defparam \tok.uart.txclkcounter_144__i6_LC_1_5_6 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_144__i6_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_144__i6_LC_1_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_144__i6_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(N__10465),
            .in2(_gnd_net_),
            .in3(N__10538),
            .lcout(\tok.uart.txclkcounter_6 ),
            .ltout(),
            .carryin(\tok.uart.n3960 ),
            .carryout(\tok.uart.n3961 ),
            .clk(N__26200),
            .ce(),
            .sr(N__12241));
    defparam \tok.uart.txclkcounter_144__i7_LC_1_5_7 .C_ON=1'b1;
    defparam \tok.uart.txclkcounter_144__i7_LC_1_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_144__i7_LC_1_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_144__i7_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(N__10435),
            .in2(_gnd_net_),
            .in3(N__10535),
            .lcout(\tok.uart.txclkcounter_7 ),
            .ltout(),
            .carryin(\tok.uart.n3961 ),
            .carryout(\tok.uart.n3962 ),
            .clk(N__26200),
            .ce(),
            .sr(N__12241));
    defparam \tok.uart.txclkcounter_144__i8_LC_1_6_0 .C_ON=1'b0;
    defparam \tok.uart.txclkcounter_144__i8_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.txclkcounter_144__i8_LC_1_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.txclkcounter_144__i8_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__10420),
            .in2(_gnd_net_),
            .in3(N__10532),
            .lcout(\tok.uart.txclkcounter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26204),
            .ce(),
            .sr(N__12242));
    defparam \tok.uart.i6_4_lut_LC_1_7_0 .C_ON=1'b0;
    defparam \tok.uart.i6_4_lut_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i6_4_lut_LC_1_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.uart.i6_4_lut_LC_1_7_0  (
            .in0(N__10529),
            .in1(N__10514),
            .in2(N__10499),
            .in3(N__10481),
            .lcout(\tok.uart.n15_adj_640 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1014_2_lut_LC_1_7_1 .C_ON=1'b0;
    defparam \tok.uart.i1014_2_lut_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1014_2_lut_LC_1_7_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.uart.i1014_2_lut_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__12206),
            .in2(_gnd_net_),
            .in3(N__16447),
            .lcout(\tok.uart.n1081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i5_3_lut_LC_1_7_2 .C_ON=1'b0;
    defparam \tok.uart.i5_3_lut_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5_3_lut_LC_1_7_2 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \tok.uart.i5_3_lut_LC_1_7_2  (
            .in0(N__10466),
            .in1(N__10451),
            .in2(_gnd_net_),
            .in3(N__10436),
            .lcout(),
            .ltout(\tok.uart.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i4705_4_lut_LC_1_7_3 .C_ON=1'b0;
    defparam \tok.uart.i4705_4_lut_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i4705_4_lut_LC_1_7_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \tok.uart.i4705_4_lut_LC_1_7_3  (
            .in0(N__10421),
            .in1(N__10406),
            .in2(N__10391),
            .in3(N__10388),
            .lcout(txtick),
            .ltout(txtick_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i4701_2_lut_LC_1_7_4 .C_ON=1'b0;
    defparam \tok.uart.i4701_2_lut_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i4701_2_lut_LC_1_7_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \tok.uart.i4701_2_lut_LC_1_7_4  (
            .in0(N__16448),
            .in1(_gnd_net_),
            .in2(N__10382),
            .in3(_gnd_net_),
            .lcout(\tok.uart.n964 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i10_LC_1_7_5 .C_ON=1'b0;
    defparam \tok.uart.sender_i10_LC_1_7_5 .SEQ_MODE=4'b1001;
    defparam \tok.uart.sender_i10_LC_1_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.sender_i10_LC_1_7_5  (
            .in0(N__17345),
            .in1(N__19648),
            .in2(_gnd_net_),
            .in3(N__11285),
            .lcout(\tok.uart.sender_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26208),
            .ce(N__16367),
            .sr(N__10628));
    defparam \tok.uart.i5_4_lut_LC_1_7_6 .C_ON=1'b0;
    defparam \tok.uart.i5_4_lut_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i5_4_lut_LC_1_7_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.uart.i5_4_lut_LC_1_7_6  (
            .in0(N__10612),
            .in1(N__10558),
            .in2(N__10598),
            .in3(N__10573),
            .lcout(\tok.uart.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rxclkcounter_147__i0_LC_1_8_0 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_147__i0_LC_1_8_0 .SEQ_MODE=4'b1001;
    defparam \tok.uart.rxclkcounter_147__i0_LC_1_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_147__i0_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__10613),
            .in2(_gnd_net_),
            .in3(N__10601),
            .lcout(\tok.uart.rxclkcounter_0 ),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(\tok.uart.n3968 ),
            .clk(N__26213),
            .ce(),
            .sr(N__11507));
    defparam \tok.uart.rxclkcounter_147__i1_LC_1_8_1 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_147__i1_LC_1_8_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_147__i1_LC_1_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_147__i1_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(N__10594),
            .in2(_gnd_net_),
            .in3(N__10580),
            .lcout(\tok.uart.rxclkcounter_1 ),
            .ltout(),
            .carryin(\tok.uart.n3968 ),
            .carryout(\tok.uart.n3969 ),
            .clk(N__26213),
            .ce(),
            .sr(N__11507));
    defparam \tok.uart.rxclkcounter_147__i2_LC_1_8_2 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_147__i2_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_147__i2_LC_1_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_147__i2_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(N__10658),
            .in2(_gnd_net_),
            .in3(N__10577),
            .lcout(\tok.uart.rxclkcounter_2 ),
            .ltout(),
            .carryin(\tok.uart.n3969 ),
            .carryout(\tok.uart.n3970 ),
            .clk(N__26213),
            .ce(),
            .sr(N__11507));
    defparam \tok.uart.rxclkcounter_147__i3_LC_1_8_3 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_147__i3_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_147__i3_LC_1_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_147__i3_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__10574),
            .in2(_gnd_net_),
            .in3(N__10562),
            .lcout(\tok.uart.rxclkcounter_3 ),
            .ltout(),
            .carryin(\tok.uart.n3970 ),
            .carryout(\tok.uart.n3971 ),
            .clk(N__26213),
            .ce(),
            .sr(N__11507));
    defparam \tok.uart.rxclkcounter_147__i4_LC_1_8_4 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_147__i4_LC_1_8_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_147__i4_LC_1_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_147__i4_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__10559),
            .in2(_gnd_net_),
            .in3(N__10547),
            .lcout(\tok.uart.rxclkcounter_4 ),
            .ltout(),
            .carryin(\tok.uart.n3971 ),
            .carryout(\tok.uart.n3972 ),
            .clk(N__26213),
            .ce(),
            .sr(N__11507));
    defparam \tok.uart.rxclkcounter_147__i5_LC_1_8_5 .C_ON=1'b1;
    defparam \tok.uart.rxclkcounter_147__i5_LC_1_8_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_147__i5_LC_1_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_147__i5_LC_1_8_5  (
            .in0(_gnd_net_),
            .in1(N__10672),
            .in2(_gnd_net_),
            .in3(N__10544),
            .lcout(\tok.uart.rxclkcounter_5 ),
            .ltout(),
            .carryin(\tok.uart.n3972 ),
            .carryout(\tok.uart.n3973 ),
            .clk(N__26213),
            .ce(),
            .sr(N__11507));
    defparam \tok.uart.rxclkcounter_147__i6_LC_1_8_6 .C_ON=1'b0;
    defparam \tok.uart.rxclkcounter_147__i6_LC_1_8_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rxclkcounter_147__i6_LC_1_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.rxclkcounter_147__i6_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(N__10685),
            .in2(_gnd_net_),
            .in3(N__10541),
            .lcout(\tok.uart.rxclkcounter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26213),
            .ce(),
            .sr(N__11507));
    defparam \tok.i2577_2_lut_3_lut_LC_1_9_0 .C_ON=1'b0;
    defparam \tok.i2577_2_lut_3_lut_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2577_2_lut_3_lut_LC_1_9_0 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \tok.i2577_2_lut_3_lut_LC_1_9_0  (
            .in0(N__23899),
            .in1(_gnd_net_),
            .in2(N__29327),
            .in3(N__19553),
            .lcout(\tok.table_wr_data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2570_2_lut_3_lut_LC_1_9_1 .C_ON=1'b0;
    defparam \tok.i2570_2_lut_3_lut_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2570_2_lut_3_lut_LC_1_9_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \tok.i2570_2_lut_3_lut_LC_1_9_1  (
            .in0(N__20402),
            .in1(N__29317),
            .in2(_gnd_net_),
            .in3(N__23895),
            .lcout(\tok.table_wr_data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2571_2_lut_3_lut_LC_1_9_2 .C_ON=1'b0;
    defparam \tok.i2571_2_lut_3_lut_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2571_2_lut_3_lut_LC_1_9_2 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \tok.i2571_2_lut_3_lut_LC_1_9_2  (
            .in0(N__23896),
            .in1(_gnd_net_),
            .in2(N__29326),
            .in3(N__20507),
            .lcout(\tok.table_wr_data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2572_2_lut_3_lut_LC_1_9_3 .C_ON=1'b0;
    defparam \tok.i2572_2_lut_3_lut_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2572_2_lut_3_lut_LC_1_9_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \tok.i2572_2_lut_3_lut_LC_1_9_3  (
            .in0(N__20596),
            .in1(N__29321),
            .in2(_gnd_net_),
            .in3(N__23897),
            .lcout(\tok.table_wr_data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i6_4_lut_adj_28_LC_1_9_4 .C_ON=1'b0;
    defparam \tok.uart.i6_4_lut_adj_28_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i6_4_lut_adj_28_LC_1_9_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \tok.uart.i6_4_lut_adj_28_LC_1_9_4  (
            .in0(N__10694),
            .in1(N__10684),
            .in2(N__10673),
            .in3(N__10657),
            .lcout(n795),
            .ltout(n795_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_1_9_5.C_ON=1'b0;
    defparam i1_2_lut_LC_1_9_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_1_9_5.LUT_INIT=16'b1111111100001111;
    LogicCell40 i1_2_lut_LC_1_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10646),
            .in3(N__11335),
            .lcout(n940),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i8_LC_1_9_6 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i8_LC_1_9_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i8_LC_1_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.uart.capture_i0_i8_LC_1_9_6  (
            .in0(N__14914),
            .in1(N__11560),
            .in2(_gnd_net_),
            .in3(N__16922),
            .lcout(capture_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26219),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2576_2_lut_3_lut_LC_1_9_7 .C_ON=1'b0;
    defparam \tok.i2576_2_lut_3_lut_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2576_2_lut_3_lut_LC_1_9_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \tok.i2576_2_lut_3_lut_LC_1_9_7  (
            .in0(N__21158),
            .in1(N__29322),
            .in2(_gnd_net_),
            .in3(N__23898),
            .lcout(\tok.table_wr_data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.bytephase__i0_LC_1_10_0 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i0_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i0_LC_1_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i0_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__11402),
            .in2(_gnd_net_),
            .in3(N__10631),
            .lcout(\tok.uart.bytephase_0 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\tok.uart.n3963 ),
            .clk(N__26227),
            .ce(N__10793),
            .sr(N__11339));
    defparam \tok.uart.bytephase__i1_LC_1_10_1 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i1_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i1_LC_1_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i1_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__11470),
            .in2(_gnd_net_),
            .in3(N__10808),
            .lcout(\tok.uart.bytephase_1 ),
            .ltout(),
            .carryin(\tok.uart.n3963 ),
            .carryout(\tok.uart.n3964 ),
            .clk(N__26227),
            .ce(N__10793),
            .sr(N__11339));
    defparam \tok.uart.bytephase__i2_LC_1_10_2 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i2_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i2_LC_1_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i2_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__11381),
            .in2(_gnd_net_),
            .in3(N__10805),
            .lcout(\tok.uart.bytephase_2 ),
            .ltout(),
            .carryin(\tok.uart.n3964 ),
            .carryout(\tok.uart.n3965 ),
            .clk(N__26227),
            .ce(N__10793),
            .sr(N__11339));
    defparam \tok.uart.bytephase__i3_LC_1_10_3 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i3_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i3_LC_1_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i3_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__11423),
            .in2(_gnd_net_),
            .in3(N__10802),
            .lcout(\tok.uart.bytephase_3 ),
            .ltout(),
            .carryin(\tok.uart.n3965 ),
            .carryout(\tok.uart.n3966 ),
            .clk(N__26227),
            .ce(N__10793),
            .sr(N__11339));
    defparam \tok.uart.bytephase__i4_LC_1_10_4 .C_ON=1'b1;
    defparam \tok.uart.bytephase__i4_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i4_LC_1_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i4_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__11360),
            .in2(_gnd_net_),
            .in3(N__10799),
            .lcout(\tok.uart.bytephase_4 ),
            .ltout(),
            .carryin(\tok.uart.n3966 ),
            .carryout(\tok.uart.n3967 ),
            .clk(N__26227),
            .ce(N__10793),
            .sr(N__11339));
    defparam \tok.uart.bytephase__i5_LC_1_10_5 .C_ON=1'b0;
    defparam \tok.uart.bytephase__i5_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.bytephase__i5_LC_1_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.uart.bytephase__i5_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__11448),
            .in2(_gnd_net_),
            .in3(N__10796),
            .lcout(\tok.uart.bytephase_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26227),
            .ce(N__10793),
            .sr(N__11339));
    defparam \tok.A_stk.tail_i0_i16_LC_2_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i16_LC_2_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i16_LC_2_2_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i16_LC_2_2_0  (
            .in0(N__10768),
            .in1(N__13816),
            .in2(N__10871),
            .in3(N__14514),
            .lcout(\tok.A_stk.tail_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26196),
            .ce(N__14726),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i0_LC_2_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i0_LC_2_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i0_LC_2_3_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tok.A_stk.tail_i0_i0_LC_2_3_1  (
            .in0(N__13779),
            .in1(N__14525),
            .in2(N__10781),
            .in3(N__29518),
            .lcout(\tok.A_stk.tail_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26198),
            .ce(N__14707),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i32_LC_2_3_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i32_LC_2_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i32_LC_2_3_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i32_LC_2_3_2  (
            .in0(N__14522),
            .in1(N__10777),
            .in2(N__10754),
            .in3(N__13782),
            .lcout(\tok.A_stk.tail_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26198),
            .ce(N__14707),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i48_LC_2_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i48_LC_2_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i48_LC_2_3_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i48_LC_2_3_3  (
            .in0(N__13780),
            .in1(N__10889),
            .in2(N__10769),
            .in3(N__14526),
            .lcout(\tok.A_stk.tail_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26198),
            .ce(N__14707),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i64_LC_2_3_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i64_LC_2_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i64_LC_2_3_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i64_LC_2_3_4  (
            .in0(N__14523),
            .in1(N__10880),
            .in2(N__10753),
            .in3(N__13783),
            .lcout(\tok.A_stk.tail_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26198),
            .ce(N__14707),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i80_LC_2_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i80_LC_2_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i80_LC_2_3_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i80_LC_2_3_5  (
            .in0(N__13781),
            .in1(N__10888),
            .in2(N__11143),
            .in3(N__14527),
            .lcout(\tok.A_stk.tail_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26198),
            .ce(N__14707),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i96_LC_2_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i96_LC_2_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i96_LC_2_3_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i96_LC_2_3_6  (
            .in0(N__14524),
            .in1(N__10879),
            .in2(N__11126),
            .in3(N__13784),
            .lcout(tail_96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26198),
            .ce(N__14707),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i0_LC_2_3_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i0_LC_2_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i0_LC_2_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i0_LC_2_3_7  (
            .in0(N__10867),
            .in1(N__15741),
            .in2(_gnd_net_),
            .in3(N__26942),
            .lcout(\tok.S_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26198),
            .ce(N__14707),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i110_LC_2_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i110_LC_2_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i110_LC_2_4_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i110_LC_2_4_0  (
            .in0(N__10852),
            .in1(N__13840),
            .in2(N__11608),
            .in3(N__14458),
            .lcout(tail_110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__14713),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i94_LC_2_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i94_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i94_LC_2_4_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i94_LC_2_4_1  (
            .in0(N__14456),
            .in1(N__10840),
            .in2(N__11629),
            .in3(N__13839),
            .lcout(\tok.A_stk.tail_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__14713),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i78_LC_2_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i78_LC_2_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i78_LC_2_4_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i78_LC_2_4_2  (
            .in0(N__10831),
            .in1(N__13842),
            .in2(N__10856),
            .in3(N__14460),
            .lcout(\tok.A_stk.tail_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__14713),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i62_LC_2_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i62_LC_2_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i62_LC_2_4_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i62_LC_2_4_3  (
            .in0(N__14455),
            .in1(N__10841),
            .in2(N__10822),
            .in3(N__13838),
            .lcout(\tok.A_stk.tail_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__14713),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i46_LC_2_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i46_LC_2_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i46_LC_2_4_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i46_LC_2_4_4  (
            .in0(N__10832),
            .in1(N__13841),
            .in2(N__10969),
            .in3(N__14459),
            .lcout(\tok.A_stk.tail_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__14713),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i30_LC_2_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i30_LC_2_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i30_LC_2_4_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i30_LC_2_4_5  (
            .in0(N__14454),
            .in1(N__10955),
            .in2(N__10823),
            .in3(N__13837),
            .lcout(\tok.A_stk.tail_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__14713),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i14_LC_2_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i14_LC_2_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i14_LC_2_4_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tok.A_stk.tail_i0_i14_LC_2_4_6  (
            .in0(N__13836),
            .in1(N__14457),
            .in2(N__10970),
            .in3(N__20456),
            .lcout(\tok.A_stk.tail_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__14713),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i14_LC_2_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i14_LC_2_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i14_LC_2_4_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i14_LC_2_4_7  (
            .in0(N__10954),
            .in1(N__15743),
            .in2(_gnd_net_),
            .in3(N__24003),
            .lcout(\tok.S_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__14713),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i104_LC_2_5_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i104_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i104_LC_2_5_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i104_LC_2_5_0  (
            .in0(N__10942),
            .in1(N__13755),
            .in2(N__11063),
            .in3(N__14428),
            .lcout(tail_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(N__14737),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i88_LC_2_5_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i88_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i88_LC_2_5_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i88_LC_2_5_1  (
            .in0(N__14426),
            .in1(N__11074),
            .in2(N__13888),
            .in3(N__10933),
            .lcout(\tok.A_stk.tail_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(N__14737),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i72_LC_2_5_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i72_LC_2_5_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i72_LC_2_5_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i72_LC_2_5_2  (
            .in0(N__10943),
            .in1(N__13757),
            .in2(N__10924),
            .in3(N__14430),
            .lcout(\tok.A_stk.tail_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(N__14737),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i56_LC_2_5_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i56_LC_2_5_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i56_LC_2_5_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i56_LC_2_5_3  (
            .in0(N__14425),
            .in1(N__10906),
            .in2(N__13887),
            .in3(N__10934),
            .lcout(\tok.A_stk.tail_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(N__14737),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i40_LC_2_5_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i40_LC_2_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i40_LC_2_5_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i40_LC_2_5_4  (
            .in0(N__10897),
            .in1(N__13756),
            .in2(N__10925),
            .in3(N__14429),
            .lcout(\tok.A_stk.tail_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(N__14737),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i24_LC_2_5_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i24_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i24_LC_2_5_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i24_LC_2_5_5  (
            .in0(N__14424),
            .in1(N__10907),
            .in2(N__13886),
            .in3(N__11156),
            .lcout(\tok.A_stk.tail_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(N__14737),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i8_LC_2_5_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i8_LC_2_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i8_LC_2_5_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i8_LC_2_5_6  (
            .in0(N__10898),
            .in1(N__14427),
            .in2(N__19554),
            .in3(N__13767),
            .lcout(\tok.A_stk.tail_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(N__14737),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i8_LC_2_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i8_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i8_LC_2_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i8_LC_2_5_7  (
            .in0(N__11155),
            .in1(N__15719),
            .in2(_gnd_net_),
            .in3(N__24854),
            .lcout(\tok.S_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(N__14737),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i112_LC_2_6_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i112_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i112_LC_2_6_1 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \tok.A_stk.tail_i0_i112_LC_2_6_1  (
            .in0(N__11122),
            .in1(N__13745),
            .in2(N__14528),
            .in3(N__11144),
            .lcout(tail_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26209),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i122_LC_2_6_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i122_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i122_LC_2_6_2 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i122_LC_2_6_2  (
            .in0(N__14445),
            .in1(N__11249),
            .in2(N__13885),
            .in3(N__10984),
            .lcout(tail_122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26209),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i121_LC_2_6_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i121_LC_2_6_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i121_LC_2_6_3 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \tok.A_stk.tail_i0_i121_LC_2_6_3  (
            .in0(N__11089),
            .in1(N__13748),
            .in2(N__14529),
            .in3(N__11108),
            .lcout(tail_121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26209),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i120_LC_2_6_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i120_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i120_LC_2_6_4 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i120_LC_2_6_4  (
            .in0(N__14444),
            .in1(N__11075),
            .in2(N__13884),
            .in3(N__11059),
            .lcout(tail_120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26209),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i119_LC_2_6_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i119_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i119_LC_2_6_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.A_stk.tail_i0_i119_LC_2_6_5  (
            .in0(N__11014),
            .in1(N__13747),
            .in2(N__11045),
            .in3(N__14447),
            .lcout(tail_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26209),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2573_2_lut_3_lut_LC_2_6_6 .C_ON=1'b0;
    defparam \tok.i2573_2_lut_3_lut_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2573_2_lut_3_lut_LC_2_6_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \tok.i2573_2_lut_3_lut_LC_2_6_6  (
            .in0(N__20752),
            .in1(N__29304),
            .in2(_gnd_net_),
            .in3(N__23900),
            .lcout(\tok.table_wr_data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i118_LC_2_6_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i118_LC_2_6_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i118_LC_2_6_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.A_stk.tail_i0_i118_LC_2_6_7  (
            .in0(N__11827),
            .in1(N__13746),
            .in2(N__11813),
            .in3(N__14446),
            .lcout(tail_118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26209),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i106_LC_2_7_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i106_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i106_LC_2_7_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i106_LC_2_7_0  (
            .in0(N__11227),
            .in1(N__13768),
            .in2(N__10988),
            .in3(N__14421),
            .lcout(tail_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26214),
            .ce(N__14738),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i90_LC_2_7_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i90_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i90_LC_2_7_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i90_LC_2_7_1  (
            .in0(N__14419),
            .in1(N__11218),
            .in2(N__11248),
            .in3(N__13891),
            .lcout(\tok.A_stk.tail_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26214),
            .ce(N__14738),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i74_LC_2_7_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i74_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i74_LC_2_7_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i74_LC_2_7_2  (
            .in0(N__11209),
            .in1(N__13770),
            .in2(N__11231),
            .in3(N__14423),
            .lcout(\tok.A_stk.tail_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26214),
            .ce(N__14738),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i58_LC_2_7_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i58_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i58_LC_2_7_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i58_LC_2_7_3  (
            .in0(N__14418),
            .in1(N__11219),
            .in2(N__11200),
            .in3(N__13890),
            .lcout(\tok.A_stk.tail_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26214),
            .ce(N__14738),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i42_LC_2_7_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i42_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i42_LC_2_7_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i42_LC_2_7_4  (
            .in0(N__11210),
            .in1(N__13769),
            .in2(N__11186),
            .in3(N__14422),
            .lcout(\tok.A_stk.tail_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26214),
            .ce(N__14738),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i26_LC_2_7_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i26_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i26_LC_2_7_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i26_LC_2_7_5  (
            .in0(N__14417),
            .in1(N__11174),
            .in2(N__11201),
            .in3(N__13889),
            .lcout(\tok.A_stk.tail_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26214),
            .ce(N__14738),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i10_LC_2_7_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i10_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i10_LC_2_7_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i10_LC_2_7_6  (
            .in0(N__11185),
            .in1(N__14420),
            .in2(N__20948),
            .in3(N__13771),
            .lcout(\tok.A_stk.tail_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26214),
            .ce(N__14738),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i10_LC_2_7_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i10_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i10_LC_2_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.A_stk.head_i0_i10_LC_2_7_7  (
            .in0(N__21068),
            .in1(N__11173),
            .in2(_gnd_net_),
            .in3(N__15745),
            .lcout(\tok.S_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26214),
            .ce(N__14738),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_7_i2_2_lut_LC_2_8_0 .C_ON=1'b0;
    defparam \tok.select_73_Select_7_i2_2_lut_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_7_i2_2_lut_LC_2_8_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.select_73_Select_7_i2_2_lut_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__21719),
            .in2(_gnd_net_),
            .in3(N__24495),
            .lcout(\tok.n2_adj_763 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_107_LC_2_8_1 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_107_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_107_LC_2_8_1 .LUT_INIT=16'b1010101111111011;
    LogicCell40 \tok.i2_4_lut_adj_107_LC_2_8_1  (
            .in0(N__13031),
            .in1(N__26615),
            .in2(N__19790),
            .in3(N__17923),
            .lcout(),
            .ltout(\tok.n13_adj_765_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_109_LC_2_8_2 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_109_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_109_LC_2_8_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i7_4_lut_adj_109_LC_2_8_2  (
            .in0(N__19673),
            .in1(N__11165),
            .in2(N__11159),
            .in3(N__29465),
            .lcout(),
            .ltout(\tok.n18_adj_767_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_111_LC_2_8_3 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_111_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_111_LC_2_8_3 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \tok.i9_4_lut_adj_111_LC_2_8_3  (
            .in0(N__24074),
            .in1(N__14783),
            .in2(N__11294),
            .in3(N__20313),
            .lcout(),
            .ltout(\tok.n20_adj_770_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_114_LC_2_8_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_114_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_114_LC_2_8_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.i1_4_lut_adj_114_LC_2_8_4  (
            .in0(N__11480),
            .in1(N__17489),
            .in2(N__11291),
            .in3(N__11981),
            .lcout(\tok.A_15_N_113_7 ),
            .ltout(\tok.A_15_N_113_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A__15__I_16_i8_3_lut_LC_2_8_5 .C_ON=1'b0;
    defparam \tok.A__15__I_16_i8_3_lut_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.A__15__I_16_i8_3_lut_LC_2_8_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \tok.A__15__I_16_i8_3_lut_LC_2_8_5  (
            .in0(N__19761),
            .in1(_gnd_net_),
            .in2(N__11288),
            .in3(N__17750),
            .lcout(\tok.A_15_N_84_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i8_LC_2_8_6 .C_ON=1'b0;
    defparam \tok.A_i8_LC_2_8_6 .SEQ_MODE=4'b1010;
    defparam \tok.A_i8_LC_2_8_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_i8_LC_2_8_6  (
            .in0(N__19674),
            .in1(N__17390),
            .in2(_gnd_net_),
            .in3(N__11279),
            .lcout(\tok.A_low_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26220),
            .ce(N__17279),
            .sr(N__19144));
    defparam \tok.i2_4_lut_adj_94_LC_2_8_7 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_94_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_94_LC_2_8_7 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \tok.i2_4_lut_adj_94_LC_2_8_7  (
            .in0(N__19757),
            .in1(N__20312),
            .in2(N__27074),
            .in3(N__17924),
            .lcout(\tok.n13_adj_748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i2_4_lut_LC_2_9_0 .C_ON=1'b0;
    defparam \tok.uart.i2_4_lut_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_4_lut_LC_2_9_0 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \tok.uart.i2_4_lut_LC_2_9_0  (
            .in0(N__11272),
            .in1(N__12153),
            .in2(N__11264),
            .in3(N__12129),
            .lcout(\tok.uart_tx_busy ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sentbits_146__i3_LC_2_9_1 .C_ON=1'b0;
    defparam \tok.uart.sentbits_146__i3_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_146__i3_LC_2_9_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \tok.uart.sentbits_146__i3_LC_2_9_1  (
            .in0(N__12131),
            .in1(N__11263),
            .in2(N__12158),
            .in3(N__11273),
            .lcout(\tok.uart.sentbits_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26228),
            .ce(N__12110),
            .sr(N__12092));
    defparam \tok.uart.sentbits_146__i2_LC_2_9_2 .C_ON=1'b0;
    defparam \tok.uart.sentbits_146__i2_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_146__i2_LC_2_9_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \tok.uart.sentbits_146__i2_LC_2_9_2  (
            .in0(N__11262),
            .in1(N__12154),
            .in2(_gnd_net_),
            .in3(N__12130),
            .lcout(\tok.uart.sentbits_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26228),
            .ce(N__12110),
            .sr(N__12092));
    defparam \tok.uart.i3_4_lut_LC_2_9_3 .C_ON=1'b0;
    defparam \tok.uart.i3_4_lut_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i3_4_lut_LC_2_9_3 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \tok.uart.i3_4_lut_LC_2_9_3  (
            .in0(N__11357),
            .in1(N__11488),
            .in2(N__11449),
            .in3(N__11420),
            .lcout(),
            .ltout(\tok.uart.n3994_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_3_lut_LC_2_9_4 .C_ON=1'b0;
    defparam \tok.uart.i1_3_lut_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_3_lut_LC_2_9_4 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \tok.uart.i1_3_lut_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__14576),
            .in2(N__11528),
            .in3(N__11561),
            .lcout(rx_data_7__N_511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i4355_2_lut_LC_2_9_5 .C_ON=1'b0;
    defparam \tok.uart.i4355_2_lut_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i4355_2_lut_LC_2_9_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \tok.uart.i4355_2_lut_LC_2_9_5  (
            .in0(N__11358),
            .in1(_gnd_net_),
            .in2(N__11450),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\tok.uart.n4506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rxrst_I_0_4_lut_LC_2_9_6 .C_ON=1'b0;
    defparam \tok.uart.rxrst_I_0_4_lut_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.rxrst_I_0_4_lut_LC_2_9_6 .LUT_INIT=16'b0011011100110011;
    LogicCell40 \tok.uart.rxrst_I_0_4_lut_LC_2_9_6  (
            .in0(N__11489),
            .in1(N__11525),
            .in2(N__11510),
            .in3(N__11495),
            .lcout(\tok.uart.rxclkcounter_6__N_477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_adj_29_LC_2_9_7 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_adj_29_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_adj_29_LC_2_9_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \tok.uart.i1_2_lut_adj_29_LC_2_9_7  (
            .in0(N__11324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11421),
            .lcout(\tok.uart.n4438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i2_2_lut_3_lut_LC_2_10_0 .C_ON=1'b0;
    defparam \tok.uart.i2_2_lut_3_lut_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i2_2_lut_3_lut_LC_2_10_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.uart.i2_2_lut_3_lut_LC_2_10_0  (
            .in0(N__11468),
            .in1(N__11399),
            .in2(_gnd_net_),
            .in3(N__11379),
            .lcout(\tok.uart.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_adj_110_LC_2_10_1 .C_ON=1'b0;
    defparam \tok.i5_3_lut_adj_110_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_adj_110_LC_2_10_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i5_3_lut_adj_110_LC_2_10_1  (
            .in0(N__16597),
            .in1(N__12314),
            .in2(_gnd_net_),
            .in3(N__27232),
            .lcout(\tok.n16_adj_769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i24_4_lut_4_lut_LC_2_10_2 .C_ON=1'b0;
    defparam \tok.uart.i24_4_lut_4_lut_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i24_4_lut_4_lut_LC_2_10_2 .LUT_INIT=16'b0100010000100000;
    LogicCell40 \tok.uart.i24_4_lut_4_lut_LC_2_10_2  (
            .in0(N__11469),
            .in1(N__11447),
            .in2(N__11323),
            .in3(N__11422),
            .lcout(),
            .ltout(\tok.uart.n13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_3_lut_4_lut_LC_2_10_3 .C_ON=1'b0;
    defparam \tok.uart.i1_3_lut_4_lut_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_3_lut_4_lut_LC_2_10_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \tok.uart.i1_3_lut_4_lut_LC_2_10_3  (
            .in0(N__11400),
            .in1(N__11380),
            .in2(N__11363),
            .in3(N__11359),
            .lcout(bytephase_5__N_510),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i9_LC_2_10_4 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i9_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i9_LC_2_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i9_LC_2_10_4  (
            .in0(N__11316),
            .in1(N__11559),
            .in2(_gnd_net_),
            .in3(N__16928),
            .lcout(capture_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26232),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i4_LC_2_10_6 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i4_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i4_LC_2_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i4_LC_2_10_6  (
            .in0(N__22138),
            .in1(N__21207),
            .in2(_gnd_net_),
            .in3(N__16926),
            .lcout(capture_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26232),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i5_LC_2_10_7 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i5_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i5_LC_2_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.capture_i0_i5_LC_2_10_7  (
            .in0(N__16927),
            .in1(N__12260),
            .in2(_gnd_net_),
            .in3(N__22137),
            .lcout(capture_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26232),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4607_4_lut_LC_2_11_0 .C_ON=1'b0;
    defparam \tok.i4607_4_lut_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4607_4_lut_LC_2_11_0 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \tok.i4607_4_lut_LC_2_11_0  (
            .in0(N__14987),
            .in1(N__21173),
            .in2(N__21089),
            .in3(N__29458),
            .lcout(\tok.n4680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_3_lut_LC_2_11_1 .C_ON=1'b0;
    defparam \tok.i50_3_lut_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i50_3_lut_LC_2_11_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.i50_3_lut_LC_2_11_1  (
            .in0(N__22589),
            .in1(N__26617),
            .in2(_gnd_net_),
            .in3(N__17922),
            .lcout(),
            .ltout(\tok.n4508_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_41_LC_2_11_2 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_41_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_41_LC_2_11_2 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \tok.i7_4_lut_adj_41_LC_2_11_2  (
            .in0(N__13193),
            .in1(N__17516),
            .in2(N__11540),
            .in3(N__11585),
            .lcout(),
            .ltout(\tok.n16_adj_660_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i10_LC_2_11_3 .C_ON=1'b0;
    defparam \tok.A_i10_LC_2_11_3 .SEQ_MODE=4'b1010;
    defparam \tok.A_i10_LC_2_11_3 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \tok.A_i10_LC_2_11_3  (
            .in0(N__17380),
            .in1(N__11537),
            .in2(N__11531),
            .in3(N__21181),
            .lcout(\tok.n59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26239),
            .ce(N__17275),
            .sr(N__19135));
    defparam \tok.A_i13_LC_2_11_4 .C_ON=1'b0;
    defparam \tok.A_i13_LC_2_11_4 .SEQ_MODE=4'b1010;
    defparam \tok.A_i13_LC_2_11_4 .LUT_INIT=16'b1111001110101010;
    LogicCell40 \tok.A_i13_LC_2_11_4  (
            .in0(N__20753),
            .in1(N__17518),
            .in2(N__11570),
            .in3(N__17381),
            .lcout(\tok.n56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26239),
            .ce(N__17275),
            .sr(N__19135));
    defparam \tok.A_i15_LC_2_11_5 .C_ON=1'b0;
    defparam \tok.A_i15_LC_2_11_5 .SEQ_MODE=4'b1010;
    defparam \tok.A_i15_LC_2_11_5 .LUT_INIT=16'b1111110001011100;
    LogicCell40 \tok.A_i15_LC_2_11_5  (
            .in0(N__17517),
            .in1(N__20495),
            .in2(N__17389),
            .in3(N__15356),
            .lcout(\tok.n54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26239),
            .ce(N__17275),
            .sr(N__19135));
    defparam \tok.i1_4_lut_adj_77_LC_2_11_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_77_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_77_LC_2_11_6 .LUT_INIT=16'b1100110100000101;
    LogicCell40 \tok.i1_4_lut_adj_77_LC_2_11_6  (
            .in0(N__26616),
            .in1(N__22588),
            .in2(N__23982),
            .in3(N__24736),
            .lcout(\tok.n12_adj_723 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_LC_2_11_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_LC_2_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i1_2_lut_LC_2_11_7  (
            .in0(N__24737),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27445),
            .lcout(\tok.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i15_1_lut_LC_2_12_0 .C_ON=1'b0;
    defparam \tok.inv_106_i15_1_lut_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i15_1_lut_LC_2_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i15_1_lut_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23952),
            .lcout(\tok.n288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_2_12_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_12_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_12_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_101_i11_2_lut_LC_2_12_2 .C_ON=1'b0;
    defparam \tok.or_101_i11_2_lut_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.or_101_i11_2_lut_LC_2_12_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.or_101_i11_2_lut_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__22719),
            .in2(_gnd_net_),
            .in3(N__28271),
            .lcout(),
            .ltout(\tok.n206_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_49_LC_2_12_3 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_49_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_49_LC_2_12_3 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \tok.i5_4_lut_adj_49_LC_2_12_3  (
            .in0(N__24497),
            .in1(N__29459),
            .in2(N__11579),
            .in3(N__20958),
            .lcout(\tok.n16_adj_673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i13_1_lut_LC_2_12_4 .C_ON=1'b0;
    defparam \tok.inv_106_i13_1_lut_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i13_1_lut_LC_2_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i13_1_lut_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22932),
            .lcout(\tok.n290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_101_i13_2_lut_LC_2_12_5 .C_ON=1'b0;
    defparam \tok.or_101_i13_2_lut_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.or_101_i13_2_lut_LC_2_12_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.or_101_i13_2_lut_LC_2_12_5  (
            .in0(N__22718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24846),
            .lcout(),
            .ltout(\tok.n204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_63_LC_2_12_6 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_63_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_63_LC_2_12_6 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \tok.i5_4_lut_adj_63_LC_2_12_6  (
            .in0(N__29460),
            .in1(N__20751),
            .in2(N__11576),
            .in3(N__24496),
            .lcout(),
            .ltout(\tok.n16_adj_699_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4676_4_lut_LC_2_12_7 .C_ON=1'b0;
    defparam \tok.i4676_4_lut_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i4676_4_lut_LC_2_12_7 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \tok.i4676_4_lut_LC_2_12_7  (
            .in0(N__22907),
            .in1(N__12410),
            .in2(N__11573),
            .in3(N__17828),
            .lcout(\tok.n4667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i124_LC_4_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i124_LC_4_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i124_LC_4_2_2 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \tok.A_stk.tail_i0_i124_LC_4_2_2  (
            .in0(N__12346),
            .in1(N__13817),
            .in2(N__12365),
            .in3(N__14513),
            .lcout(tail_124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26202),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i18_LC_4_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i18_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i18_LC_4_3_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i18_LC_4_3_0  (
            .in0(N__11684),
            .in1(N__13703),
            .in2(N__11645),
            .in3(N__14488),
            .lcout(\tok.A_stk.tail_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26206),
            .ce(N__14703),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i34_LC_4_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i34_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i34_LC_4_3_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i34_LC_4_3_1  (
            .in0(N__14484),
            .in1(N__11692),
            .in2(N__13873),
            .in3(N__11674),
            .lcout(\tok.A_stk.tail_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26206),
            .ce(N__14703),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i2_LC_4_3_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i2_LC_4_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i2_LC_4_3_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i2_LC_4_3_2  (
            .in0(N__11693),
            .in1(N__14487),
            .in2(N__20028),
            .in3(N__13715),
            .lcout(\tok.A_stk.tail_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26206),
            .ce(N__14703),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i50_LC_4_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i50_LC_4_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i50_LC_4_3_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i50_LC_4_3_3  (
            .in0(N__14485),
            .in1(N__11683),
            .in2(N__13874),
            .in3(N__11663),
            .lcout(\tok.A_stk.tail_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26206),
            .ce(N__14703),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i66_LC_4_3_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i66_LC_4_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i66_LC_4_3_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i66_LC_4_3_4  (
            .in0(N__11654),
            .in1(N__13704),
            .in2(N__11675),
            .in3(N__14489),
            .lcout(\tok.A_stk.tail_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26206),
            .ce(N__14703),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i82_LC_4_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i82_LC_4_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i82_LC_4_3_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i82_LC_4_3_5  (
            .in0(N__14486),
            .in1(N__11755),
            .in2(N__13875),
            .in3(N__11662),
            .lcout(\tok.A_stk.tail_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26206),
            .ce(N__14703),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i98_LC_4_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i98_LC_4_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i98_LC_4_3_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i98_LC_4_3_6  (
            .in0(N__11653),
            .in1(N__13705),
            .in2(N__11744),
            .in3(N__14490),
            .lcout(tail_98),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26206),
            .ce(N__14703),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i2_LC_4_3_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i2_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i2_LC_4_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i2_LC_4_3_7  (
            .in0(N__11641),
            .in1(N__15720),
            .in2(_gnd_net_),
            .in3(N__21987),
            .lcout(\tok.S_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26206),
            .ce(N__14703),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i126_LC_4_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i126_LC_4_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i126_LC_4_4_0 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \tok.A_stk.tail_i0_i126_LC_4_4_0  (
            .in0(N__11630),
            .in1(N__13860),
            .in2(N__11609),
            .in3(N__14338),
            .lcout(tail_126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26210),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i125_LC_4_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i125_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i125_LC_4_4_1 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i125_LC_4_4_1  (
            .in0(N__14335),
            .in1(N__11717),
            .in2(N__13928),
            .in3(N__11729),
            .lcout(tail_125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26210),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i117_LC_4_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i117_LC_4_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i117_LC_4_4_3 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i117_LC_4_4_3  (
            .in0(N__14334),
            .in1(N__12725),
            .in2(N__13927),
            .in3(N__12739),
            .lcout(tail_117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26210),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i116_LC_4_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i116_LC_4_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i116_LC_4_4_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.A_stk.tail_i0_i116_LC_4_4_4  (
            .in0(N__12826),
            .in1(N__13859),
            .in2(N__12812),
            .in3(N__14337),
            .lcout(tail_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26210),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i2_LC_4_4_5 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i2_LC_4_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i2_LC_4_4_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i2_LC_4_4_5  (
            .in0(N__16708),
            .in1(N__22121),
            .in2(_gnd_net_),
            .in3(N__17200),
            .lcout(uart_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26210),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i114_LC_4_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i114_LC_4_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i114_LC_4_4_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.A_stk.tail_i0_i114_LC_4_4_6  (
            .in0(N__11743),
            .in1(N__13858),
            .in2(N__11759),
            .in3(N__14336),
            .lcout(tail_114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26210),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i115_LC_4_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i115_LC_4_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i115_LC_4_4_7 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \tok.A_stk.tail_i0_i115_LC_4_4_7  (
            .in0(N__14333),
            .in1(N__12703),
            .in2(N__13926),
            .in3(N__12542),
            .lcout(tail_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26210),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i109_LC_4_5_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i109_LC_4_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i109_LC_4_5_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \tok.A_stk.tail_i0_i109_LC_4_5_0  (
            .in0(N__11701),
            .in1(N__11728),
            .in2(N__13922),
            .in3(N__14519),
            .lcout(tail_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26215),
            .ce(N__14727),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i93_LC_4_5_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i93_LC_4_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i93_LC_4_5_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i93_LC_4_5_1  (
            .in0(N__14517),
            .in1(N__11716),
            .in2(N__13925),
            .in3(N__11881),
            .lcout(\tok.A_stk.tail_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26215),
            .ce(N__14727),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i77_LC_4_5_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i77_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i77_LC_4_5_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i77_LC_4_5_2  (
            .in0(N__11872),
            .in1(N__13847),
            .in2(N__11705),
            .in3(N__14521),
            .lcout(\tok.A_stk.tail_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26215),
            .ce(N__14727),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i61_LC_4_5_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i61_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i61_LC_4_5_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i61_LC_4_5_3  (
            .in0(N__14516),
            .in1(N__11863),
            .in2(N__13924),
            .in3(N__11882),
            .lcout(\tok.A_stk.tail_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26215),
            .ce(N__14727),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i45_LC_4_5_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i45_LC_4_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i45_LC_4_5_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i45_LC_4_5_4  (
            .in0(N__11873),
            .in1(N__13846),
            .in2(N__11855),
            .in3(N__14520),
            .lcout(\tok.A_stk.tail_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26215),
            .ce(N__14727),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i29_LC_4_5_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i29_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i29_LC_4_5_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i29_LC_4_5_5  (
            .in0(N__14515),
            .in1(N__11843),
            .in2(N__13923),
            .in3(N__11864),
            .lcout(\tok.A_stk.tail_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26215),
            .ce(N__14727),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i13_LC_4_5_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i13_LC_4_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i13_LC_4_5_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i13_LC_4_5_6  (
            .in0(N__11854),
            .in1(N__14518),
            .in2(N__20564),
            .in3(N__13857),
            .lcout(\tok.A_stk.tail_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26215),
            .ce(N__14727),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i13_LC_4_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i13_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i13_LC_4_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i13_LC_4_5_7  (
            .in0(N__11842),
            .in1(N__15682),
            .in2(_gnd_net_),
            .in3(N__20680),
            .lcout(\tok.S_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26215),
            .ce(N__14727),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i102_LC_4_6_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i102_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i102_LC_4_6_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i102_LC_4_6_0  (
            .in0(N__11788),
            .in1(N__13801),
            .in2(N__11831),
            .in3(N__14510),
            .lcout(tail_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26223),
            .ce(N__14708),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i86_LC_4_6_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i86_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i86_LC_4_6_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i86_LC_4_6_1  (
            .in0(N__14508),
            .in1(N__11779),
            .in2(N__11809),
            .in3(N__13872),
            .lcout(\tok.A_stk.tail_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26223),
            .ce(N__14708),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i70_LC_4_6_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i70_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i70_LC_4_6_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i70_LC_4_6_2  (
            .in0(N__11789),
            .in1(N__13803),
            .in2(N__11771),
            .in3(N__14512),
            .lcout(\tok.A_stk.tail_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26223),
            .ce(N__14708),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i54_LC_4_6_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i54_LC_4_6_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i54_LC_4_6_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i54_LC_4_6_3  (
            .in0(N__14507),
            .in1(N__11780),
            .in2(N__11968),
            .in3(N__13871),
            .lcout(\tok.A_stk.tail_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26223),
            .ce(N__14708),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i38_LC_4_6_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i38_LC_4_6_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i38_LC_4_6_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i38_LC_4_6_4  (
            .in0(N__11770),
            .in1(N__13802),
            .in2(N__11953),
            .in3(N__14511),
            .lcout(\tok.A_stk.tail_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26223),
            .ce(N__14708),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i22_LC_4_6_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i22_LC_4_6_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i22_LC_4_6_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i22_LC_4_6_5  (
            .in0(N__14506),
            .in1(N__11939),
            .in2(N__11969),
            .in3(N__13870),
            .lcout(\tok.A_stk.tail_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26223),
            .ce(N__14708),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i6_LC_4_6_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i6_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i6_LC_4_6_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i6_LC_4_6_6  (
            .in0(N__21269),
            .in1(N__14509),
            .in2(N__11954),
            .in3(N__13800),
            .lcout(\tok.A_stk.tail_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26223),
            .ce(N__14708),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i6_LC_4_6_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i6_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i6_LC_4_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_stk.head_i0_i6_LC_4_6_7  (
            .in0(N__15732),
            .in1(N__11938),
            .in2(_gnd_net_),
            .in3(N__28255),
            .lcout(\tok.S_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26223),
            .ce(N__14708),
            .sr(_gnd_net_));
    defparam \tok.i12_4_lut_LC_4_7_0 .C_ON=1'b0;
    defparam \tok.i12_4_lut_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i12_4_lut_LC_4_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i12_4_lut_LC_4_7_0  (
            .in0(N__12026),
            .in1(N__12074),
            .in2(N__12041),
            .in3(N__12062),
            .lcout(\tok.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_198_LC_4_7_1 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_198_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_198_LC_4_7_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i4_4_lut_adj_198_LC_4_7_1  (
            .in0(N__11926),
            .in1(N__11917),
            .in2(N__22403),
            .in3(N__21840),
            .lcout(),
            .ltout(\tok.n20_adj_803_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_136_LC_4_7_2 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_136_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_136_LC_4_7_2 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \tok.i10_4_lut_adj_136_LC_4_7_2  (
            .in0(N__24835),
            .in1(N__11908),
            .in2(N__11930),
            .in3(N__12953),
            .lcout(\tok.n26_adj_805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_80_LC_4_7_3 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_80_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_80_LC_4_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i10_4_lut_adj_80_LC_4_7_3  (
            .in0(N__11927),
            .in1(N__11918),
            .in2(N__11909),
            .in3(N__12967),
            .lcout(\tok.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_86_LC_4_7_4 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_86_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_86_LC_4_7_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_86_LC_4_7_4  (
            .in0(N__15094),
            .in1(N__15043),
            .in2(N__15121),
            .in3(N__15067),
            .lcout(),
            .ltout(\tok.n25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i15_4_lut_adj_178_LC_4_7_5 .C_ON=1'b0;
    defparam \tok.i15_4_lut_adj_178_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i15_4_lut_adj_178_LC_4_7_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i15_4_lut_adj_178_LC_4_7_5  (
            .in0(N__12947),
            .in1(N__11897),
            .in2(N__11891),
            .in3(N__11888),
            .lcout(\tok.found_slot_N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_51_LC_4_8_0 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_51_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_51_LC_4_8_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i7_4_lut_adj_51_LC_4_8_0  (
            .in0(N__12073),
            .in1(N__12061),
            .in2(N__24009),
            .in3(N__21429),
            .lcout(\tok.n23_adj_677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i12_1_lut_LC_4_8_1 .C_ON=1'b0;
    defparam \tok.inv_106_i12_1_lut_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i12_1_lut_LC_4_8_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \tok.inv_106_i12_1_lut_LC_4_8_1  (
            .in0(N__21430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2574_2_lut_3_lut_LC_4_8_2 .C_ON=1'b0;
    defparam \tok.i2574_2_lut_3_lut_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2574_2_lut_3_lut_LC_4_8_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \tok.i2574_2_lut_3_lut_LC_4_8_2  (
            .in0(N__20842),
            .in1(N__29265),
            .in2(_gnd_net_),
            .in3(N__23878),
            .lcout(\tok.table_wr_data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_4_lut_LC_4_8_3 .C_ON=1'b0;
    defparam \tok.i8_4_lut_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i8_4_lut_LC_4_8_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i8_4_lut_LC_4_8_3  (
            .in0(N__12037),
            .in1(N__12025),
            .in2(N__20311),
            .in3(N__22636),
            .lcout(\tok.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1512_3_lut_4_lut_LC_4_8_4 .C_ON=1'b0;
    defparam \tok.i1512_3_lut_4_lut_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1512_3_lut_4_lut_LC_4_8_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \tok.i1512_3_lut_4_lut_LC_4_8_4  (
            .in0(N__18890),
            .in1(N__29260),
            .in2(N__19691),
            .in3(N__23875),
            .lcout(\tok.table_wr_data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i8_1_lut_LC_4_8_5 .C_ON=1'b0;
    defparam \tok.inv_106_i8_1_lut_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i8_1_lut_LC_4_8_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \tok.inv_106_i8_1_lut_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(N__19774),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1623_3_lut_4_lut_LC_4_8_6 .C_ON=1'b0;
    defparam \tok.i1623_3_lut_4_lut_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1623_3_lut_4_lut_LC_4_8_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \tok.i1623_3_lut_4_lut_LC_4_8_6  (
            .in0(N__24375),
            .in1(N__29261),
            .in2(N__25307),
            .in3(N__23876),
            .lcout(\tok.table_wr_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1734_3_lut_4_lut_LC_4_8_7 .C_ON=1'b0;
    defparam \tok.i1734_3_lut_4_lut_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1734_3_lut_4_lut_LC_4_8_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \tok.i1734_3_lut_4_lut_LC_4_8_7  (
            .in0(N__23877),
            .in1(N__18650),
            .in2(N__29291),
            .in3(N__20154),
            .lcout(\tok.table_wr_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_112_LC_4_9_0 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_112_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_112_LC_4_9_0 .LUT_INIT=16'b1111010011111000;
    LogicCell40 \tok.i4_4_lut_adj_112_LC_4_9_0  (
            .in0(N__21977),
            .in1(N__24726),
            .in2(N__19592),
            .in3(N__28834),
            .lcout(\tok.n15_adj_771 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i3_1_lut_LC_4_9_1 .C_ON=1'b0;
    defparam \tok.inv_106_i3_1_lut_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i3_1_lut_LC_4_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i3_1_lut_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21976),
            .lcout(\tok.n300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i4707_2_lut_3_lut_LC_4_9_2 .C_ON=1'b0;
    defparam \tok.uart.i4707_2_lut_3_lut_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i4707_2_lut_3_lut_LC_4_9_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \tok.uart.i4707_2_lut_3_lut_LC_4_9_2  (
            .in0(N__19344),
            .in1(N__12239),
            .in2(_gnd_net_),
            .in3(N__16423),
            .lcout(\tok.uart.n1083 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_LC_4_9_3 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_LC_4_9_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.uart.i1_2_lut_LC_4_9_3  (
            .in0(N__28835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16079),
            .lcout(),
            .ltout(\tok.uart.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i4698_4_lut_LC_4_9_4 .C_ON=1'b0;
    defparam \tok.uart.i4698_4_lut_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i4698_4_lut_LC_4_9_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \tok.uart.i4698_4_lut_LC_4_9_4  (
            .in0(N__19343),
            .in1(N__28014),
            .in2(N__12164),
            .in3(N__30441),
            .lcout(n23),
            .ltout(n23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_3_lut_LC_4_9_5 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_3_lut_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_3_lut_LC_4_9_5 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \tok.uart.i1_2_lut_3_lut_LC_4_9_5  (
            .in0(N__12240),
            .in1(_gnd_net_),
            .in2(N__12161),
            .in3(N__19345),
            .lcout(\tok.uart.n978 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sentbits_146__i0_LC_4_9_6 .C_ON=1'b0;
    defparam \tok.uart.sentbits_146__i0_LC_4_9_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_146__i0_LC_4_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.uart.sentbits_146__i0_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12151),
            .lcout(\tok.uart.sentbits_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26240),
            .ce(N__12109),
            .sr(N__12088));
    defparam \tok.uart.sentbits_146__i1_LC_4_9_7 .C_ON=1'b0;
    defparam \tok.uart.sentbits_146__i1_LC_4_9_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sentbits_146__i1_LC_4_9_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \tok.uart.sentbits_146__i1_LC_4_9_7  (
            .in0(N__12152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12128),
            .lcout(\tok.uart.sentbits_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26240),
            .ce(N__12109),
            .sr(N__12088));
    defparam \tok.i5_4_lut_adj_203_LC_4_10_0 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_203_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_203_LC_4_10_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i5_4_lut_adj_203_LC_4_10_0  (
            .in0(N__20953),
            .in1(N__22969),
            .in2(N__20761),
            .in3(N__21047),
            .lcout(\tok.n21_adj_857 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i5_LC_4_10_1 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i5_LC_4_10_1 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i5_LC_4_10_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i5_LC_4_10_1  (
            .in0(N__12256),
            .in1(N__22101),
            .in2(_gnd_net_),
            .in3(N__15322),
            .lcout(uart_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26244),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i3_LC_4_10_2 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i3_LC_4_10_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i3_LC_4_10_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.capture_i0_i3_LC_4_10_2  (
            .in0(N__16701),
            .in1(N__16942),
            .in2(_gnd_net_),
            .in3(N__21214),
            .lcout(capture_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26244),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_4_lut_adj_200_LC_4_10_3 .C_ON=1'b0;
    defparam \tok.i8_4_lut_adj_200_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i8_4_lut_adj_200_LC_4_10_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i8_4_lut_adj_200_LC_4_10_3  (
            .in0(N__21169),
            .in1(N__20280),
            .in2(N__20400),
            .in3(N__22631),
            .lcout(\tok.n24_adj_854 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i7_LC_4_10_4 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i7_LC_4_10_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i7_LC_4_10_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.capture_i0_i7_LC_4_10_4  (
            .in0(N__12270),
            .in1(N__16944),
            .in2(_gnd_net_),
            .in3(N__14929),
            .lcout(capture_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26244),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i6_LC_4_10_5 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i6_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i6_LC_4_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.rx_data_i0_i6_LC_4_10_5  (
            .in0(N__21340),
            .in1(N__12272),
            .in2(_gnd_net_),
            .in3(N__22102),
            .lcout(uart_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26244),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i6_LC_4_10_6 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i6_LC_4_10_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i6_LC_4_10_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.capture_i0_i6_LC_4_10_6  (
            .in0(N__12271),
            .in1(N__16943),
            .in2(_gnd_net_),
            .in3(N__12255),
            .lcout(capture_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26244),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i2_LC_4_10_7 .C_ON=1'b0;
    defparam \tok.uart.sender_i2_LC_4_10_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i2_LC_4_10_7 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \tok.uart.sender_i2_LC_4_10_7  (
            .in0(N__12232),
            .in1(N__13300),
            .in2(N__16268),
            .in3(N__16427),
            .lcout(sender_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26244),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_2_lut_LC_4_11_0 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_2_lut_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_2_lut_LC_4_11_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_2_lut_LC_4_11_0  (
            .in0(N__17088),
            .in1(N__13139),
            .in2(N__29571),
            .in3(N__12185),
            .lcout(\tok.n6_adj_684 ),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\tok.n3910 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_3_lut_LC_4_11_1 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_3_lut_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_3_lut_LC_4_11_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_3_lut_LC_4_11_1  (
            .in0(N__17643),
            .in1(N__14963),
            .in2(N__20170),
            .in3(N__12182),
            .lcout(\tok.n10_adj_786 ),
            .ltout(),
            .carryin(\tok.n3910 ),
            .carryout(\tok.n3911 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_4_lut_LC_4_11_2 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_4_lut_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_4_lut_LC_4_11_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_4_lut_LC_4_11_2  (
            .in0(N__17086),
            .in1(N__12179),
            .in2(N__20064),
            .in3(N__12170),
            .lcout(\tok.n6_adj_667 ),
            .ltout(),
            .carryin(\tok.n3911 ),
            .carryout(\tok.n3912 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_5_lut_LC_4_11_3 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_5_lut_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_5_lut_LC_4_11_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_5_lut_LC_4_11_3  (
            .in0(N__17642),
            .in1(N__15419),
            .in2(N__21550),
            .in3(N__12167),
            .lcout(\tok.n9_adj_836 ),
            .ltout(),
            .carryin(\tok.n3912 ),
            .carryout(\tok.n3913 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_6_lut_LC_4_11_4 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_6_lut_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_6_lut_LC_4_11_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_6_lut_LC_4_11_4  (
            .in0(N__17644),
            .in1(N__24367),
            .in2(N__13220),
            .in3(N__12332),
            .lcout(\tok.n3_adj_826 ),
            .ltout(),
            .carryin(\tok.n3913 ),
            .carryout(\tok.n3914 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_7_lut_LC_4_11_5 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_7_lut_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_7_lut_LC_4_11_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_7_lut_LC_4_11_5  (
            .in0(N__17090),
            .in1(N__15452),
            .in2(N__19946),
            .in3(N__12329),
            .lcout(\tok.n6_adj_814 ),
            .ltout(),
            .carryin(\tok.n3914 ),
            .carryout(\tok.n3915 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_8_lut_LC_4_11_6 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_8_lut_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_8_lut_LC_4_11_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_8_lut_LC_4_11_6  (
            .in0(N__17087),
            .in1(N__21299),
            .in2(N__22739),
            .in3(N__12326),
            .lcout(\tok.n6_adj_780 ),
            .ltout(),
            .carryin(\tok.n3915 ),
            .carryout(\tok.n3916 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_9_lut_LC_4_11_7 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_9_lut_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_9_lut_LC_4_11_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_9_lut_LC_4_11_7  (
            .in0(N__17089),
            .in1(N__12323),
            .in2(N__19689),
            .in3(N__12302),
            .lcout(\tok.n6_adj_768 ),
            .ltout(),
            .carryin(\tok.n3916 ),
            .carryout(\tok.n3917 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_10_lut_LC_4_12_0 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_10_lut_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_10_lut_LC_4_12_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_10_lut_LC_4_12_0  (
            .in0(N__17109),
            .in1(N__19563),
            .in2(N__13247),
            .in3(N__12299),
            .lcout(\tok.n6_adj_653 ),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\tok.n3918 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_11_lut_LC_4_12_1 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_11_lut_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_11_lut_LC_4_12_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_11_lut_LC_4_12_1  (
            .in0(N__17645),
            .in1(N__21180),
            .in2(N__14873),
            .in3(N__12296),
            .lcout(\tok.n13_adj_657 ),
            .ltout(),
            .carryin(\tok.n3918 ),
            .carryout(\tok.n3919 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_12_lut_LC_4_12_2 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_12_lut_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_12_lut_LC_4_12_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_12_lut_LC_4_12_2  (
            .in0(N__17111),
            .in1(N__12377),
            .in2(N__20966),
            .in3(N__12293),
            .lcout(\tok.n6_adj_676 ),
            .ltout(),
            .carryin(\tok.n3919 ),
            .carryout(\tok.n3920 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_13_lut_LC_4_12_3 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_13_lut_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_13_lut_LC_4_12_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_13_lut_LC_4_12_3  (
            .in0(N__17113),
            .in1(N__20867),
            .in2(N__12290),
            .in3(N__12275),
            .lcout(\tok.n6_adj_692 ),
            .ltout(),
            .carryin(\tok.n3920 ),
            .carryout(\tok.n3921 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_14_lut_LC_4_12_4 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_14_lut_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_14_lut_LC_4_12_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_14_lut_LC_4_12_4  (
            .in0(N__17110),
            .in1(N__20762),
            .in2(N__12422),
            .in3(N__12401),
            .lcout(\tok.n6_adj_701 ),
            .ltout(),
            .carryin(\tok.n3921 ),
            .carryout(\tok.n3922 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_15_lut_LC_4_12_5 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_15_lut_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_15_lut_LC_4_12_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_15_lut_LC_4_12_5  (
            .in0(N__17112),
            .in1(N__20563),
            .in2(N__13211),
            .in3(N__12398),
            .lcout(\tok.n6_adj_711 ),
            .ltout(),
            .carryin(\tok.n3922 ),
            .carryout(\tok.n3923 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_16_lut_LC_4_12_6 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_16_lut_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_16_lut_LC_4_12_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_105_add_2_16_lut_LC_4_12_6  (
            .in0(N__17108),
            .in1(N__20505),
            .in2(N__12395),
            .in3(N__12383),
            .lcout(\tok.n6_adj_731 ),
            .ltout(),
            .carryin(\tok.n3923 ),
            .carryout(\tok.n3924 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_16_THRU_CRY_0_LC_4_12_7 .C_ON=1'b1;
    defparam \tok.sub_105_add_2_16_THRU_CRY_0_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_16_THRU_CRY_0_LC_4_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \tok.sub_105_add_2_16_THRU_CRY_0_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(N__21610),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\tok.n3924 ),
            .carryout(\tok.n3924_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_add_2_17_lut_LC_4_13_0 .C_ON=1'b0;
    defparam \tok.sub_105_add_2_17_lut_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_add_2_17_lut_LC_4_13_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \tok.sub_105_add_2_17_lut_LC_4_13_0  (
            .in0(N__12371),
            .in1(N__20401),
            .in2(N__17117),
            .in3(N__12380),
            .lcout(\tok.n6_adj_753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i11_1_lut_LC_4_13_1 .C_ON=1'b0;
    defparam \tok.inv_106_i11_1_lut_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i11_1_lut_LC_4_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i11_1_lut_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21059),
            .lcout(\tok.n292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i16_1_lut_LC_4_13_3 .C_ON=1'b0;
    defparam \tok.inv_106_i16_1_lut_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i16_1_lut_LC_4_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i16_1_lut_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20305),
            .lcout(\tok.n287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i108_LC_5_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i108_LC_5_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i108_LC_5_2_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i108_LC_5_2_0  (
            .in0(N__14410),
            .in1(N__12520),
            .in2(N__12364),
            .in3(N__13504),
            .lcout(tail_108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26207),
            .ce(N__14681),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i92_LC_5_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i92_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i92_LC_5_2_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i92_LC_5_2_1  (
            .in0(N__13502),
            .in1(N__12511),
            .in2(N__12347),
            .in3(N__14416),
            .lcout(\tok.A_stk.tail_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26207),
            .ce(N__14681),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i76_LC_5_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i76_LC_5_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i76_LC_5_2_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i76_LC_5_2_2  (
            .in0(N__14413),
            .in1(N__12521),
            .in2(N__12503),
            .in3(N__13506),
            .lcout(\tok.A_stk.tail_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26207),
            .ce(N__14681),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i60_LC_5_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i60_LC_5_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i60_LC_5_2_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i60_LC_5_2_3  (
            .in0(N__13501),
            .in1(N__12512),
            .in2(N__12484),
            .in3(N__14415),
            .lcout(\tok.A_stk.tail_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26207),
            .ce(N__14681),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i44_LC_5_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i44_LC_5_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i44_LC_5_2_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i44_LC_5_2_4  (
            .in0(N__14412),
            .in1(N__12499),
            .in2(N__12469),
            .in3(N__13505),
            .lcout(\tok.A_stk.tail_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26207),
            .ce(N__14681),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i28_LC_5_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i28_LC_5_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i28_LC_5_2_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i28_LC_5_2_5  (
            .in0(N__13500),
            .in1(N__12455),
            .in2(N__12485),
            .in3(N__14414),
            .lcout(\tok.A_stk.tail_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26207),
            .ce(N__14681),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i12_LC_5_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i12_LC_5_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i12_LC_5_2_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tok.A_stk.tail_i0_i12_LC_5_2_6  (
            .in0(N__14411),
            .in1(N__13503),
            .in2(N__12470),
            .in3(N__20723),
            .lcout(\tok.A_stk.tail_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26207),
            .ce(N__14681),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i12_LC_5_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i12_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i12_LC_5_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i12_LC_5_2_7  (
            .in0(N__12454),
            .in1(N__15739),
            .in2(_gnd_net_),
            .in3(N__23006),
            .lcout(\tok.S_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26207),
            .ce(N__14681),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i17_LC_5_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i17_LC_5_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i17_LC_5_3_0 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \tok.A_stk.tail_i0_i17_LC_5_3_0  (
            .in0(N__12431),
            .in1(N__12551),
            .in2(N__13876),
            .in3(N__14242),
            .lcout(\tok.A_stk.tail_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26211),
            .ce(N__14664),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i1_LC_5_3_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i1_LC_5_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i1_LC_5_3_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i1_LC_5_3_1  (
            .in0(N__14239),
            .in1(N__12442),
            .in2(N__13723),
            .in3(N__20113),
            .lcout(\tok.A_stk.tail_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26211),
            .ce(N__14664),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i33_LC_5_3_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i33_LC_5_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i33_LC_5_3_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i33_LC_5_3_2  (
            .in0(N__12580),
            .in1(N__13524),
            .in2(N__12443),
            .in3(N__14243),
            .lcout(\tok.A_stk.tail_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26211),
            .ce(N__14664),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i49_LC_5_3_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i49_LC_5_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i49_LC_5_3_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i49_LC_5_3_3  (
            .in0(N__14240),
            .in1(N__12430),
            .in2(N__13724),
            .in3(N__12569),
            .lcout(\tok.A_stk.tail_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26211),
            .ce(N__14664),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i65_LC_5_3_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i65_LC_5_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i65_LC_5_3_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i65_LC_5_3_4  (
            .in0(N__12560),
            .in1(N__13525),
            .in2(N__12581),
            .in3(N__14244),
            .lcout(\tok.A_stk.tail_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26211),
            .ce(N__14664),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i81_LC_5_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i81_LC_5_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i81_LC_5_3_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i81_LC_5_3_5  (
            .in0(N__14241),
            .in1(N__13960),
            .in2(N__13725),
            .in3(N__12568),
            .lcout(\tok.A_stk.tail_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26211),
            .ce(N__14664),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i97_LC_5_3_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i97_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i97_LC_5_3_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i97_LC_5_3_6  (
            .in0(N__12559),
            .in1(N__13526),
            .in2(N__13949),
            .in3(N__14245),
            .lcout(tail_97),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26211),
            .ce(N__14664),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i1_LC_5_3_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i1_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i1_LC_5_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i1_LC_5_3_7  (
            .in0(N__12550),
            .in1(N__15740),
            .in2(_gnd_net_),
            .in3(N__24188),
            .lcout(\tok.S_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26211),
            .ce(N__14664),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i99_LC_5_4_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i99_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i99_LC_5_4_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i99_LC_5_4_0  (
            .in0(N__14235),
            .in1(N__12541),
            .in2(N__13729),
            .in3(N__12688),
            .lcout(tail_99),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26216),
            .ce(N__14682),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i35_LC_5_4_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i35_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i35_LC_5_4_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i35_LC_5_4_1  (
            .in0(N__12530),
            .in1(N__13537),
            .in2(N__12653),
            .in3(N__14237),
            .lcout(\tok.A_stk.tail_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26216),
            .ce(N__14682),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i67_LC_5_4_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i67_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i67_LC_5_4_2 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i67_LC_5_4_2  (
            .in0(N__14233),
            .in1(N__12529),
            .in2(N__13727),
            .in3(N__12689),
            .lcout(\tok.A_stk.tail_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26216),
            .ce(N__14682),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i3_LC_5_4_3 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i3_LC_5_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i3_LC_5_4_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i3_LC_5_4_3  (
            .in0(N__12667),
            .in1(N__15724),
            .in2(_gnd_net_),
            .in3(N__21851),
            .lcout(\tok.S_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26216),
            .ce(N__14682),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i51_LC_5_4_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i51_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i51_LC_5_4_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i51_LC_5_4_4  (
            .in0(N__14232),
            .in1(N__12679),
            .in2(N__13726),
            .in3(N__12713),
            .lcout(\tok.A_stk.tail_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26216),
            .ce(N__14682),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i101_LC_5_4_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i101_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i101_LC_5_4_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i101_LC_5_4_5  (
            .in0(N__12634),
            .in1(N__13536),
            .in2(N__12740),
            .in3(N__14236),
            .lcout(tail_101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26216),
            .ce(N__14682),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i85_LC_5_4_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i85_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i85_LC_5_4_6 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i85_LC_5_4_6  (
            .in0(N__14234),
            .in1(N__12724),
            .in2(N__13728),
            .in3(N__12622),
            .lcout(\tok.A_stk.tail_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26216),
            .ce(N__14682),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i83_LC_5_4_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i83_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i83_LC_5_4_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i83_LC_5_4_7  (
            .in0(N__12712),
            .in1(N__13538),
            .in2(N__12704),
            .in3(N__14238),
            .lcout(\tok.A_stk.tail_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26216),
            .ce(N__14682),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i3_LC_5_5_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i3_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i3_LC_5_5_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tok.A_stk.tail_i0_i3_LC_5_5_0  (
            .in0(N__14247),
            .in1(N__13641),
            .in2(N__12652),
            .in3(N__21491),
            .lcout(\tok.A_stk.tail_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26224),
            .ce(N__14712),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i19_LC_5_5_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i19_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i19_LC_5_5_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i19_LC_5_5_1  (
            .in0(N__13638),
            .in1(N__12680),
            .in2(N__12668),
            .in3(N__14250),
            .lcout(\tok.A_stk.tail_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26224),
            .ce(N__14712),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i69_LC_5_5_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i69_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i69_LC_5_5_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i69_LC_5_5_2  (
            .in0(N__14249),
            .in1(N__12635),
            .in2(N__12607),
            .in3(N__13644),
            .lcout(\tok.A_stk.tail_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26224),
            .ce(N__14712),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i53_LC_5_5_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i53_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i53_LC_5_5_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i53_LC_5_5_3  (
            .in0(N__13640),
            .in1(N__12593),
            .in2(N__12623),
            .in3(N__14252),
            .lcout(\tok.A_stk.tail_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26224),
            .ce(N__14712),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i37_LC_5_5_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i37_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i37_LC_5_5_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i37_LC_5_5_4  (
            .in0(N__14246),
            .in1(N__12847),
            .in2(N__12608),
            .in3(N__13643),
            .lcout(\tok.A_stk.tail_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26224),
            .ce(N__14712),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i21_LC_5_5_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i21_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i21_LC_5_5_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i21_LC_5_5_5  (
            .in0(N__13639),
            .in1(N__12592),
            .in2(N__12839),
            .in3(N__14251),
            .lcout(\tok.A_stk.tail_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26224),
            .ce(N__14712),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i5_LC_5_5_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i5_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i5_LC_5_5_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tok.A_stk.tail_i0_i5_LC_5_5_6  (
            .in0(N__14248),
            .in1(N__13642),
            .in2(N__19919),
            .in3(N__12848),
            .lcout(\tok.A_stk.tail_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26224),
            .ce(N__14712),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i5_LC_5_5_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i5_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i5_LC_5_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i5_LC_5_5_7  (
            .in0(N__12835),
            .in1(N__15681),
            .in2(_gnd_net_),
            .in3(N__22402),
            .lcout(\tok.S_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26224),
            .ce(N__14712),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i100_LC_5_6_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i100_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i100_LC_5_6_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \tok.A_stk.tail_i0_i100_LC_5_6_0  (
            .in0(N__12790),
            .in1(N__12827),
            .in2(N__13905),
            .in3(N__14385),
            .lcout(tail_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26229),
            .ce(N__14722),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i84_LC_5_6_1 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i84_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i84_LC_5_6_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i84_LC_5_6_1  (
            .in0(N__14383),
            .in1(N__12805),
            .in2(N__12781),
            .in3(N__13815),
            .lcout(\tok.A_stk.tail_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26229),
            .ce(N__14722),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i68_LC_5_6_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i68_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i68_LC_5_6_2 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i68_LC_5_6_2  (
            .in0(N__12791),
            .in1(N__14387),
            .in2(N__13907),
            .in3(N__12766),
            .lcout(\tok.A_stk.tail_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26229),
            .ce(N__14722),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i52_LC_5_6_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i52_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i52_LC_5_6_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \tok.A_stk.tail_i0_i52_LC_5_6_3  (
            .in0(N__14382),
            .in1(N__12757),
            .in2(N__12782),
            .in3(N__13814),
            .lcout(\tok.A_stk.tail_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26229),
            .ce(N__14722),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i36_LC_5_6_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i36_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i36_LC_5_6_4 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \tok.A_stk.tail_i0_i36_LC_5_6_4  (
            .in0(N__12748),
            .in1(N__14386),
            .in2(N__13906),
            .in3(N__12767),
            .lcout(\tok.A_stk.tail_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26229),
            .ce(N__14722),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i20_LC_5_6_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i20_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i20_LC_5_6_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i20_LC_5_6_5  (
            .in0(N__14381),
            .in1(N__12758),
            .in2(N__13013),
            .in3(N__13813),
            .lcout(\tok.A_stk.tail_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26229),
            .ce(N__14722),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i4_LC_5_6_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i4_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i4_LC_5_6_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i4_LC_5_6_6  (
            .in0(N__12749),
            .in1(N__14384),
            .in2(N__24376),
            .in3(N__13645),
            .lcout(\tok.A_stk.tail_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26229),
            .ce(N__14722),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i4_LC_5_6_7 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i4_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i4_LC_5_6_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_stk.head_i0_i4_LC_5_6_7  (
            .in0(N__13009),
            .in1(N__15731),
            .in2(_gnd_net_),
            .in3(N__27434),
            .lcout(\tok.S_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26229),
            .ce(N__14722),
            .sr(_gnd_net_));
    defparam \tok.i14_4_lut_LC_5_7_0 .C_ON=1'b0;
    defparam \tok.i14_4_lut_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i14_4_lut_LC_5_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i14_4_lut_LC_5_7_0  (
            .in0(N__12857),
            .in1(N__12902),
            .in2(N__13001),
            .in3(N__12992),
            .lcout(),
            .ltout(\tok.n30_adj_824_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4597_4_lut_LC_5_7_1 .C_ON=1'b0;
    defparam \tok.i4597_4_lut_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i4597_4_lut_LC_5_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i4597_4_lut_LC_5_7_1  (
            .in0(N__12986),
            .in1(N__15080),
            .in2(N__12980),
            .in3(N__15029),
            .lcout(),
            .ltout(\tok.n4642_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_190_LC_5_7_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_190_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_190_LC_5_7_2 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \tok.i1_4_lut_adj_190_LC_5_7_2  (
            .in0(N__12977),
            .in1(N__14855),
            .in2(N__12971),
            .in3(N__22519),
            .lcout(\tok.found_slot ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.key_rd_15__I_0_241_i14_2_lut_LC_5_7_3 .C_ON=1'b0;
    defparam \tok.key_rd_15__I_0_241_i14_2_lut_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.key_rd_15__I_0_241_i14_2_lut_LC_5_7_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.key_rd_15__I_0_241_i14_2_lut_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(N__12968),
            .in2(_gnd_net_),
            .in3(N__20677),
            .lcout(\tok.n14_adj_804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i11_4_lut_adj_85_LC_5_7_4 .C_ON=1'b0;
    defparam \tok.i11_4_lut_adj_85_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i11_4_lut_adj_85_LC_5_7_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i11_4_lut_adj_85_LC_5_7_4  (
            .in0(N__12919),
            .in1(N__12877),
            .in2(N__12941),
            .in3(N__12895),
            .lcout(\tok.n27_adj_734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_70_LC_5_7_5 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_70_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_70_LC_5_7_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i5_4_lut_adj_70_LC_5_7_5  (
            .in0(N__12940),
            .in1(N__21034),
            .in2(N__12923),
            .in3(N__22979),
            .lcout(\tok.n21_adj_714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_44_LC_5_7_7 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_44_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_44_LC_5_7_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i6_4_lut_adj_44_LC_5_7_7  (
            .in0(N__12896),
            .in1(N__12881),
            .in2(N__19812),
            .in3(N__21967),
            .lcout(\tok.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_2_lut_LC_5_8_0 .C_ON=1'b1;
    defparam \tok.add_109_2_lut_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_2_lut_LC_5_8_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_2_lut_LC_5_8_0  (
            .in0(N__29078),
            .in1(N__29548),
            .in2(_gnd_net_),
            .in3(N__12851),
            .lcout(\tok.n10_adj_679 ),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\tok.n3940 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_3_lut_LC_5_8_1 .C_ON=1'b1;
    defparam \tok.add_109_3_lut_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_3_lut_LC_5_8_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_3_lut_LC_5_8_1  (
            .in0(N__23746),
            .in1(N__20150),
            .in2(_gnd_net_),
            .in3(N__13049),
            .lcout(\tok.n28_adj_821 ),
            .ltout(),
            .carryin(\tok.n3940 ),
            .carryout(\tok.n3941 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_4_lut_LC_5_8_2 .C_ON=1'b1;
    defparam \tok.add_109_4_lut_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_4_lut_LC_5_8_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_4_lut_LC_5_8_2  (
            .in0(N__29077),
            .in1(N__20035),
            .in2(_gnd_net_),
            .in3(N__13046),
            .lcout(\tok.n10_adj_818 ),
            .ltout(),
            .carryin(\tok.n3941 ),
            .carryout(\tok.n3942 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_5_lut_LC_5_8_3 .C_ON=1'b1;
    defparam \tok.add_109_5_lut_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_5_lut_LC_5_8_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_5_lut_LC_5_8_3  (
            .in0(N__23745),
            .in1(_gnd_net_),
            .in2(N__21540),
            .in3(N__13043),
            .lcout(\tok.n6_adj_812 ),
            .ltout(),
            .carryin(\tok.n3942 ),
            .carryout(\tok.n3943 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_6_lut_LC_5_8_4 .C_ON=1'b1;
    defparam \tok.add_109_6_lut_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_6_lut_LC_5_8_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_6_lut_LC_5_8_4  (
            .in0(N__23744),
            .in1(N__24366),
            .in2(_gnd_net_),
            .in3(N__13040),
            .lcout(\tok.n9_adj_807 ),
            .ltout(),
            .carryin(\tok.n3943 ),
            .carryout(\tok.n3944 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_7_lut_LC_5_8_5 .C_ON=1'b1;
    defparam \tok.add_109_7_lut_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_7_lut_LC_5_8_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_7_lut_LC_5_8_5  (
            .in0(N__29080),
            .in1(N__19906),
            .in2(_gnd_net_),
            .in3(N__13037),
            .lcout(\tok.n10_adj_806 ),
            .ltout(),
            .carryin(\tok.n3944 ),
            .carryout(\tok.n3945 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_8_lut_LC_5_8_6 .C_ON=1'b1;
    defparam \tok.add_109_8_lut_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_8_lut_LC_5_8_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_8_lut_LC_5_8_6  (
            .in0(N__29079),
            .in1(N__21298),
            .in2(_gnd_net_),
            .in3(N__13034),
            .lcout(\tok.n10_adj_783 ),
            .ltout(),
            .carryin(\tok.n3945 ),
            .carryout(\tok.n3946 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_9_lut_LC_5_8_7 .C_ON=1'b1;
    defparam \tok.add_109_9_lut_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_9_lut_LC_5_8_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_9_lut_LC_5_8_7  (
            .in0(N__29081),
            .in1(N__19679),
            .in2(_gnd_net_),
            .in3(N__13022),
            .lcout(\tok.n10_adj_764 ),
            .ltout(),
            .carryin(\tok.n3946 ),
            .carryout(\tok.n3947 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_10_lut_LC_5_9_0 .C_ON=1'b1;
    defparam \tok.add_109_10_lut_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_10_lut_LC_5_9_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_10_lut_LC_5_9_0  (
            .in0(N__29103),
            .in1(N__19549),
            .in2(_gnd_net_),
            .in3(N__13019),
            .lcout(\tok.n10_adj_652 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\tok.n3948 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_11_lut_LC_5_9_1 .C_ON=1'b1;
    defparam \tok.add_109_11_lut_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_11_lut_LC_5_9_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_11_lut_LC_5_9_1  (
            .in0(N__23750),
            .in1(N__21168),
            .in2(_gnd_net_),
            .in3(N__13016),
            .lcout(\tok.n10_adj_656 ),
            .ltout(),
            .carryin(\tok.n3948 ),
            .carryout(\tok.n3949 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_12_lut_LC_5_9_2 .C_ON=1'b1;
    defparam \tok.add_109_12_lut_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_12_lut_LC_5_9_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_12_lut_LC_5_9_2  (
            .in0(N__29105),
            .in1(N__20952),
            .in2(_gnd_net_),
            .in3(N__13097),
            .lcout(\tok.n10_adj_671 ),
            .ltout(),
            .carryin(\tok.n3949 ),
            .carryout(\tok.n3950 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_13_lut_LC_5_9_3 .C_ON=1'b1;
    defparam \tok.add_109_13_lut_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_13_lut_LC_5_9_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_13_lut_LC_5_9_3  (
            .in0(N__29108),
            .in1(N__20853),
            .in2(_gnd_net_),
            .in3(N__13094),
            .lcout(\tok.n4674 ),
            .ltout(),
            .carryin(\tok.n3950 ),
            .carryout(\tok.n3951 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_14_lut_LC_5_9_4 .C_ON=1'b1;
    defparam \tok.add_109_14_lut_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_14_lut_LC_5_9_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_14_lut_LC_5_9_4  (
            .in0(N__29102),
            .in1(N__20732),
            .in2(_gnd_net_),
            .in3(N__13091),
            .lcout(\tok.n10_adj_697 ),
            .ltout(),
            .carryin(\tok.n3951 ),
            .carryout(\tok.n3952 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_15_lut_LC_5_9_5 .C_ON=1'b1;
    defparam \tok.add_109_15_lut_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_15_lut_LC_5_9_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_15_lut_LC_5_9_5  (
            .in0(N__29107),
            .in1(N__20587),
            .in2(_gnd_net_),
            .in3(N__13088),
            .lcout(\tok.n10_adj_705 ),
            .ltout(),
            .carryin(\tok.n3952 ),
            .carryout(\tok.n3953 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_16_lut_LC_5_9_6 .C_ON=1'b1;
    defparam \tok.add_109_16_lut_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_16_lut_LC_5_9_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_109_16_lut_LC_5_9_6  (
            .in0(N__29104),
            .in1(N__20506),
            .in2(_gnd_net_),
            .in3(N__13085),
            .lcout(\tok.n4661 ),
            .ltout(),
            .carryin(\tok.n3953 ),
            .carryout(\tok.n3954 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_109_17_lut_LC_5_9_7 .C_ON=1'b0;
    defparam \tok.add_109_17_lut_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_109_17_lut_LC_5_9_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \tok.add_109_17_lut_LC_5_9_7  (
            .in0(N__20395),
            .in1(N__29106),
            .in2(_gnd_net_),
            .in3(N__13082),
            .lcout(\tok.n4656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_15_i2_3_lut_LC_5_10_0 .C_ON=1'b0;
    defparam \tok.select_73_Select_15_i2_3_lut_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_15_i2_3_lut_LC_5_10_0 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \tok.select_73_Select_15_i2_3_lut_LC_5_10_0  (
            .in0(N__22717),
            .in1(N__21402),
            .in2(_gnd_net_),
            .in3(N__24494),
            .lcout(),
            .ltout(\tok.n2_adj_739_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_89_LC_5_10_1 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_89_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_89_LC_5_10_1 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \tok.i3_4_lut_adj_89_LC_5_10_1  (
            .in0(N__21403),
            .in1(N__28348),
            .in2(N__13079),
            .in3(N__26810),
            .lcout(),
            .ltout(\tok.n14_adj_741_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_96_LC_5_10_2 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_96_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_96_LC_5_10_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_96_LC_5_10_2  (
            .in0(N__13076),
            .in1(N__15254),
            .in2(N__13064),
            .in3(N__13061),
            .lcout(),
            .ltout(\tok.n20_adj_754_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4673_4_lut_LC_5_10_3 .C_ON=1'b0;
    defparam \tok.i4673_4_lut_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4673_4_lut_LC_5_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i4673_4_lut_LC_5_10_3  (
            .in0(N__13181),
            .in1(N__13145),
            .in2(N__13175),
            .in3(N__13172),
            .lcout(\tok.n4653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_15_i9_2_lut_LC_5_10_4 .C_ON=1'b0;
    defparam \tok.select_73_Select_15_i9_2_lut_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_15_i9_2_lut_LC_5_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.select_73_Select_15_i9_2_lut_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__20394),
            .in2(_gnd_net_),
            .in3(N__29461),
            .lcout(\tok.n9_adj_749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_adj_95_LC_5_10_5 .C_ON=1'b0;
    defparam \tok.i5_3_lut_adj_95_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_adj_95_LC_5_10_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i5_3_lut_adj_95_LC_5_10_5  (
            .in0(N__13163),
            .in1(N__20213),
            .in2(_gnd_net_),
            .in3(N__27245),
            .lcout(\tok.n16_adj_751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_105_inv_0_i1_1_lut_LC_5_10_6 .C_ON=1'b0;
    defparam \tok.sub_105_inv_0_i1_1_lut_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_105_inv_0_i1_1_lut_LC_5_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.sub_105_inv_0_i1_1_lut_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26899),
            .lcout(\tok.n17_adj_774 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_65_LC_5_10_7 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_65_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_65_LC_5_10_7 .LUT_INIT=16'b1010101011101111;
    LogicCell40 \tok.i4_4_lut_adj_65_LC_5_10_7  (
            .in0(N__13133),
            .in1(N__22632),
            .in2(N__28349),
            .in3(N__26811),
            .lcout(\tok.n16_adj_706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_57_LC_5_11_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_57_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_57_LC_5_11_0 .LUT_INIT=16'b1111000100010001;
    LogicCell40 \tok.i1_4_lut_adj_57_LC_5_11_0  (
            .in0(N__21400),
            .in1(N__26598),
            .in2(N__28270),
            .in3(N__24727),
            .lcout(\tok.n12_adj_687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_58_LC_5_11_1 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_58_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_58_LC_5_11_1 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \tok.i2_4_lut_adj_58_LC_5_11_1  (
            .in0(N__21841),
            .in1(N__21401),
            .in2(N__27072),
            .in3(N__17921),
            .lcout(),
            .ltout(\tok.n13_adj_688_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_59_LC_5_11_2 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_59_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_59_LC_5_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_59_LC_5_11_2  (
            .in0(N__13124),
            .in1(N__13310),
            .in2(N__13118),
            .in3(N__13115),
            .lcout(),
            .ltout(\tok.n20_adj_693_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4672_4_lut_LC_5_11_3 .C_ON=1'b0;
    defparam \tok.i4672_4_lut_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4672_4_lut_LC_5_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i4672_4_lut_LC_5_11_3  (
            .in0(N__17978),
            .in1(N__13109),
            .in2(N__13100),
            .in3(N__15134),
            .lcout(\tok.n4671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_adj_177_LC_5_11_5 .C_ON=1'b0;
    defparam \tok.i5_3_lut_adj_177_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_adj_177_LC_5_11_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i5_3_lut_adj_177_LC_5_11_5  (
            .in0(N__25792),
            .in1(N__13256),
            .in2(_gnd_net_),
            .in3(N__27242),
            .lcout(\tok.n16_adj_845 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i9_1_lut_LC_5_11_6 .C_ON=1'b0;
    defparam \tok.inv_106_i9_1_lut_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i9_1_lut_LC_5_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \tok.inv_106_i9_1_lut_LC_5_11_6  (
            .in0(N__24785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1660_3_lut_4_lut_LC_5_12_0 .C_ON=1'b0;
    defparam \tok.i1660_3_lut_4_lut_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1660_3_lut_4_lut_LC_5_12_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \tok.i1660_3_lut_4_lut_LC_5_12_0  (
            .in0(N__23893),
            .in1(N__21539),
            .in2(N__23627),
            .in3(N__29305),
            .lcout(\tok.table_wr_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i5_1_lut_LC_5_12_1 .C_ON=1'b0;
    defparam \tok.inv_106_i5_1_lut_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i5_1_lut_LC_5_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i5_1_lut_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27427),
            .lcout(\tok.n298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i14_1_lut_LC_5_12_2 .C_ON=1'b0;
    defparam \tok.inv_106_i14_1_lut_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i14_1_lut_LC_5_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i14_1_lut_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20652),
            .lcout(\tok.n289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_adj_145_LC_5_12_3 .C_ON=1'b0;
    defparam \tok.i5_3_lut_adj_145_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_adj_145_LC_5_12_3 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \tok.i5_3_lut_adj_145_LC_5_12_3  (
            .in0(N__13202),
            .in1(N__23428),
            .in2(_gnd_net_),
            .in3(N__27243),
            .lcout(\tok.n16_adj_820 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_LC_5_12_4 .C_ON=1'b0;
    defparam \tok.i1_3_lut_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_LC_5_12_4 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \tok.i1_3_lut_LC_5_12_4  (
            .in0(N__22701),
            .in1(N__22375),
            .in2(_gnd_net_),
            .in3(N__24493),
            .lcout(),
            .ltout(\tok.n34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_LC_5_12_5 .C_ON=1'b0;
    defparam \tok.i4_4_lut_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_LC_5_12_5 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \tok.i4_4_lut_LC_5_12_5  (
            .in0(N__22376),
            .in1(N__28344),
            .in2(N__13196),
            .in3(N__26816),
            .lcout(\tok.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_11_i2_3_lut_LC_5_12_6 .C_ON=1'b0;
    defparam \tok.select_73_Select_11_i2_3_lut_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_11_i2_3_lut_LC_5_12_6 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \tok.select_73_Select_11_i2_3_lut_LC_5_12_6  (
            .in0(N__19806),
            .in1(_gnd_net_),
            .in2(N__22716),
            .in3(N__24492),
            .lcout(),
            .ltout(\tok.n2_adj_685_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_56_LC_5_12_7 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_56_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_56_LC_5_12_7 .LUT_INIT=16'b1111000011111101;
    LogicCell40 \tok.i3_4_lut_adj_56_LC_5_12_7  (
            .in0(N__28337),
            .in1(N__19807),
            .in2(N__13313),
            .in3(N__26815),
            .lcout(\tok.n14_adj_686 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i1_LC_5_13_4 .C_ON=1'b0;
    defparam \tok.uart.sender_i1_LC_5_13_4 .SEQ_MODE=4'b1001;
    defparam \tok.uart.sender_i1_LC_5_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tok.uart.sender_i1_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13304),
            .lcout(tx_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26263),
            .ce(N__16386),
            .sr(N__16465));
    defparam \tok.reset_I_0_1_lut_LC_5_14_1 .C_ON=1'b0;
    defparam \tok.reset_I_0_1_lut_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \tok.reset_I_0_1_lut_LC_5_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.reset_I_0_1_lut_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13280),
            .lcout(\tok.reset_N_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i111_LC_6_2_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i111_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i111_LC_6_2_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i111_LC_6_2_0  (
            .in0(N__14005),
            .in1(N__13511),
            .in2(N__13985),
            .in3(N__14407),
            .lcout(tail_111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26212),
            .ce(N__14680),
            .sr(_gnd_net_));
    defparam \tok.A_stk.head_i0_i15_LC_6_2_1 .C_ON=1'b0;
    defparam \tok.A_stk.head_i0_i15_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.head_i0_i15_LC_6_2_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A_stk.head_i0_i15_LC_6_2_1  (
            .in0(N__20310),
            .in1(N__15712),
            .in2(_gnd_net_),
            .in3(N__14026),
            .lcout(\tok.S_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26212),
            .ce(N__14680),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i79_LC_6_2_2 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i79_LC_6_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i79_LC_6_2_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tok.A_stk.tail_i0_i79_LC_6_2_2  (
            .in0(N__13273),
            .in1(N__13513),
            .in2(N__14009),
            .in3(N__14409),
            .lcout(\tok.A_stk.tail_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26212),
            .ce(N__14680),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i63_LC_6_2_3 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i63_LC_6_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i63_LC_6_2_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i63_LC_6_2_3  (
            .in0(N__14404),
            .in1(N__13264),
            .in2(N__13721),
            .in3(N__14018),
            .lcout(\tok.A_stk.tail_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26212),
            .ce(N__14680),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i47_LC_6_2_4 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i47_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i47_LC_6_2_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i47_LC_6_2_4  (
            .in0(N__13274),
            .in1(N__13512),
            .in2(N__14039),
            .in3(N__14408),
            .lcout(\tok.A_stk.tail_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26212),
            .ce(N__14680),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i31_LC_6_2_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i31_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i31_LC_6_2_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tok.A_stk.tail_i0_i31_LC_6_2_5  (
            .in0(N__14403),
            .in1(N__14027),
            .in2(N__13720),
            .in3(N__13265),
            .lcout(\tok.A_stk.tail_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26212),
            .ce(N__14680),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i15_LC_6_2_6 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i15_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i15_LC_6_2_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tok.A_stk.tail_i0_i15_LC_6_2_6  (
            .in0(N__14038),
            .in1(N__14406),
            .in2(N__20369),
            .in3(N__13523),
            .lcout(\tok.A_stk.tail_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26212),
            .ce(N__14680),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i95_LC_6_2_7 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i95_LC_6_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i95_LC_6_2_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \tok.A_stk.tail_i0_i95_LC_6_2_7  (
            .in0(N__14405),
            .in1(N__13996),
            .in2(N__13722),
            .in3(N__14017),
            .lcout(\tok.A_stk.tail_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26212),
            .ce(N__14680),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i127_LC_6_3_0 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i127_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i127_LC_6_3_0 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \tok.A_stk.tail_i0_i127_LC_6_3_0  (
            .in0(N__14135),
            .in1(N__13981),
            .in2(N__13719),
            .in3(N__13997),
            .lcout(tail_127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26217),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_189_LC_6_3_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_189_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_189_LC_6_3_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_189_LC_6_3_1  (
            .in0(N__22520),
            .in1(N__15941),
            .in2(_gnd_net_),
            .in3(N__28832),
            .lcout(\tok.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i58_LC_6_3_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i58_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i58_LC_6_3_2 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i58_LC_6_3_2  (
            .in0(N__15478),
            .in1(N__25598),
            .in2(N__16580),
            .in3(N__25422),
            .lcout(\tok.tail_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26217),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i57_LC_6_3_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i57_LC_6_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i57_LC_6_3_3 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \tok.C_stk.tail_i0_i57_LC_6_3_3  (
            .in0(N__25420),
            .in1(N__15491),
            .in2(N__25660),
            .in3(N__15512),
            .lcout(\tok.tail_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26217),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i56_LC_6_3_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i56_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i56_LC_6_3_4 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i56_LC_6_3_4  (
            .in0(N__18493),
            .in1(N__25597),
            .in2(N__18470),
            .in3(N__25421),
            .lcout(\tok.tail_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26217),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.tail_i0_i113_LC_6_3_5 .C_ON=1'b0;
    defparam \tok.A_stk.tail_i0_i113_LC_6_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.A_stk.tail_i0_i113_LC_6_3_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \tok.A_stk.tail_i0_i113_LC_6_3_5  (
            .in0(N__13945),
            .in1(N__13507),
            .in2(N__13964),
            .in3(N__14136),
            .lcout(tail_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26217),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_4_lut_LC_6_3_6 .C_ON=1'b0;
    defparam \tok.i2_3_lut_4_lut_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_4_lut_LC_6_3_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \tok.i2_3_lut_4_lut_LC_6_3_6  (
            .in0(N__28833),
            .in1(N__15597),
            .in2(N__16631),
            .in3(N__28691),
            .lcout(n29),
            .ltout(n29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_stk.i567_2_lut_LC_6_3_7 .C_ON=1'b0;
    defparam \tok.A_stk.i567_2_lut_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \tok.A_stk.i567_2_lut_LC_6_3_7 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \tok.A_stk.i567_2_lut_LC_6_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14741),
            .in3(N__14134),
            .lcout(\tok.A_stk.rd_15__N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_103_LC_6_4_0 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_103_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_103_LC_6_4_0 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_103_LC_6_4_0  (
            .in0(N__23110),
            .in1(N__30448),
            .in2(N__15224),
            .in3(N__30163),
            .lcout(),
            .ltout(\tok.n83_adj_735_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4602_2_lut_3_lut_LC_6_4_1 .C_ON=1'b0;
    defparam \tok.i4602_2_lut_3_lut_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.i4602_2_lut_3_lut_LC_6_4_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i4602_2_lut_3_lut_LC_6_4_1  (
            .in0(_gnd_net_),
            .in1(N__29029),
            .in2(N__14588),
            .in3(N__29869),
            .lcout(\tok.n4649 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_155_LC_6_4_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_155_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_155_LC_6_4_2 .LUT_INIT=16'b1011111101111111;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_155_LC_6_4_2  (
            .in0(N__29868),
            .in1(N__30447),
            .in2(N__28544),
            .in3(N__30162),
            .lcout(),
            .ltout(\tok.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_69_LC_6_4_3 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_69_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_69_LC_6_4_3 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \tok.i5_4_lut_adj_69_LC_6_4_3  (
            .in0(N__14582),
            .in1(N__14557),
            .in2(N__14585),
            .in3(N__29028),
            .lcout(\tok.n2503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4364_2_lut_LC_6_4_4 .C_ON=1'b0;
    defparam \tok.i4364_2_lut_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4364_2_lut_LC_6_4_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \tok.i4364_2_lut_LC_6_4_4  (
            .in0(N__28015),
            .in1(N__28689),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n4516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i0_LC_6_4_5 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i0_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i0_LC_6_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.capture_i0_i0_LC_6_4_5  (
            .in0(N__17180),
            .in1(N__14572),
            .in2(_gnd_net_),
            .in3(N__16960),
            .lcout(capture_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26225),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_LC_6_4_6 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_LC_6_4_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.i1_3_lut_4_lut_LC_6_4_6  (
            .in0(N__28517),
            .in1(N__28690),
            .in2(N__30452),
            .in3(N__30164),
            .lcout(),
            .ltout(\tok.n4_adj_654_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_173_LC_6_4_7 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_173_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_173_LC_6_4_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i2_4_lut_adj_173_LC_6_4_7  (
            .in0(N__14558),
            .in1(N__28016),
            .in2(N__14546),
            .in3(N__29030),
            .lcout(n786),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_72_LC_6_5_0 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_72_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_72_LC_6_5_0 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \tok.i125_4_lut_adj_72_LC_6_5_0  (
            .in0(N__16801),
            .in1(N__30146),
            .in2(N__17563),
            .in3(N__30417),
            .lcout(),
            .ltout(\tok.n83_adj_716_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4631_2_lut_3_lut_LC_6_5_1 .C_ON=1'b0;
    defparam \tok.i4631_2_lut_3_lut_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i4631_2_lut_3_lut_LC_6_5_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \tok.i4631_2_lut_3_lut_LC_6_5_1  (
            .in0(N__29854),
            .in1(_gnd_net_),
            .in2(N__14804),
            .in3(N__28999),
            .lcout(\tok.n4690 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_2_lut_LC_6_5_2 .C_ON=1'b0;
    defparam \tok.i26_2_lut_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i26_2_lut_LC_6_5_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.i26_2_lut_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(N__30145),
            .in2(_gnd_net_),
            .in3(N__29853),
            .lcout(),
            .ltout(\tok.n12_adj_740_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_134_LC_6_5_3 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_134_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_134_LC_6_5_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \tok.i5_4_lut_adj_134_LC_6_5_3  (
            .in0(N__30416),
            .in1(N__14795),
            .in2(N__14801),
            .in3(N__15599),
            .lcout(),
            .ltout(\tok.n12_adj_801_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_153_LC_6_5_4 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_153_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_153_LC_6_5_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \tok.i6_4_lut_adj_153_LC_6_5_4  (
            .in0(N__28523),
            .in1(N__28822),
            .in2(N__14798),
            .in3(N__27999),
            .lcout(\tok.n240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i226_2_lut_LC_6_5_5 .C_ON=1'b0;
    defparam \tok.i226_2_lut_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i226_2_lut_LC_6_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i226_2_lut_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(N__28678),
            .in2(_gnd_net_),
            .in3(N__28998),
            .lcout(\tok.n284 ),
            .ltout(\tok.n284_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_99_i8_3_lut_4_lut_LC_6_5_6 .C_ON=1'b0;
    defparam \tok.or_99_i8_3_lut_4_lut_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i8_3_lut_4_lut_LC_6_5_6 .LUT_INIT=16'b1111111011001101;
    LogicCell40 \tok.or_99_i8_3_lut_4_lut_LC_6_5_6  (
            .in0(N__28524),
            .in1(N__21846),
            .in2(N__14789),
            .in3(N__28821),
            .lcout(),
            .ltout(\tok.n182_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_108_LC_6_5_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_108_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_108_LC_6_5_7 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \tok.i1_4_lut_adj_108_LC_6_5_7  (
            .in0(N__14899),
            .in1(N__27067),
            .in2(N__14786),
            .in3(N__26812),
            .lcout(\tok.n12_adj_766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i14_4_lut_adj_208_LC_6_6_0 .C_ON=1'b0;
    defparam \tok.i14_4_lut_adj_208_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i14_4_lut_adj_208_LC_6_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i14_4_lut_adj_208_LC_6_6_0  (
            .in0(N__16088),
            .in1(N__16058),
            .in2(N__14771),
            .in3(N__14756),
            .lcout(),
            .ltout(\tok.n30_adj_862_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_210_LC_6_6_1 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_210_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_210_LC_6_6_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \tok.i1_3_lut_adj_210_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__14942),
            .in2(N__14744),
            .in3(N__26486),
            .lcout(\tok.n4051 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_207_LC_6_6_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_207_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_207_LC_6_6_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i1_4_lut_adj_207_LC_6_6_2  (
            .in0(N__28253),
            .in1(N__29549),
            .in2(N__21303),
            .in3(N__26928),
            .lcout(\tok.n17_adj_861 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_206_LC_6_6_3 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_206_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_206_LC_6_6_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i3_4_lut_adj_206_LC_6_6_3  (
            .in0(N__20679),
            .in1(N__19555),
            .in2(N__20583),
            .in3(N__24794),
            .lcout(),
            .ltout(\tok.n19_adj_860_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i13_4_lut_LC_6_6_4 .C_ON=1'b0;
    defparam \tok.i13_4_lut_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i13_4_lut_LC_6_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i13_4_lut_LC_6_6_4  (
            .in0(N__15431),
            .in1(N__16094),
            .in2(N__14951),
            .in3(N__14948),
            .lcout(\tok.n29_adj_864 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i7_LC_6_6_6 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i7_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i7_LC_6_6_6 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \tok.uart.rx_data_i0_i7_LC_6_6_6  (
            .in0(N__14936),
            .in1(N__22114),
            .in2(N__14903),
            .in3(_gnd_net_),
            .lcout(uart_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26235),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2575_2_lut_3_lut_LC_6_7_0 .C_ON=1'b0;
    defparam \tok.i2575_2_lut_3_lut_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2575_2_lut_3_lut_LC_6_7_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \tok.i2575_2_lut_3_lut_LC_6_7_0  (
            .in0(N__29281),
            .in1(N__20947),
            .in2(_gnd_net_),
            .in3(N__23871),
            .lcout(\tok.table_wr_data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i10_1_lut_LC_6_7_1 .C_ON=1'b0;
    defparam \tok.inv_106_i10_1_lut_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i10_1_lut_LC_6_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i10_1_lut_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22650),
            .lcout(\tok.n293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2580_3_lut_LC_6_7_2 .C_ON=1'b0;
    defparam \tok.i2580_3_lut_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2580_3_lut_LC_6_7_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \tok.i2580_3_lut_LC_6_7_2  (
            .in0(N__29279),
            .in1(N__23869),
            .in2(_gnd_net_),
            .in3(N__26416),
            .lcout(\tok.n2634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_4_lut_LC_6_7_3 .C_ON=1'b0;
    defparam \tok.i2_2_lut_4_lut_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_4_lut_LC_6_7_3 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \tok.i2_2_lut_4_lut_LC_6_7_3  (
            .in0(N__26417),
            .in1(N__19371),
            .in2(N__23894),
            .in3(N__29282),
            .lcout(\tok.write_slot ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1586_3_lut_4_lut_LC_6_7_4 .C_ON=1'b0;
    defparam \tok.i1586_3_lut_4_lut_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1586_3_lut_4_lut_LC_6_7_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \tok.i1586_3_lut_4_lut_LC_6_7_4  (
            .in0(N__29280),
            .in1(N__23383),
            .in2(N__19950),
            .in3(N__23870),
            .lcout(\tok.table_wr_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_97_LC_6_7_5 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_97_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_97_LC_6_7_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \tok.i2_4_lut_adj_97_LC_6_7_5  (
            .in0(N__24131),
            .in1(N__15122),
            .in2(N__15101),
            .in3(N__27435),
            .lcout(\tok.n18_adj_756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i1_2_lut_3_lut_4_lut_LC_6_7_6 .C_ON=1'b0;
    defparam \tok.uart.i1_2_lut_3_lut_4_lut_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i1_2_lut_3_lut_4_lut_LC_6_7_6 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \tok.uart.i1_2_lut_3_lut_4_lut_LC_6_7_6  (
            .in0(N__29283),
            .in1(N__22112),
            .in2(N__19313),
            .in3(N__27806),
            .lcout(\tok.uart.n922 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4599_4_lut_LC_6_7_7 .C_ON=1'b0;
    defparam \tok.i4599_4_lut_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i4599_4_lut_LC_6_7_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i4599_4_lut_LC_6_7_7  (
            .in0(N__15074),
            .in1(N__28259),
            .in2(N__15053),
            .in3(N__26929),
            .lcout(\tok.n4645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_39_LC_6_8_0 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_39_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_39_LC_6_8_0 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \tok.i2_4_lut_adj_39_LC_6_8_0  (
            .in0(N__15020),
            .in1(N__15008),
            .in2(N__24149),
            .in3(N__27804),
            .lcout(),
            .ltout(\tok.n30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_40_LC_6_8_1 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_40_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_40_LC_6_8_1 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \tok.i3_4_lut_adj_40_LC_6_8_1  (
            .in0(N__15002),
            .in1(N__29258),
            .in2(N__14990),
            .in3(N__27244),
            .lcout(\tok.n12_adj_659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.valid_54_LC_6_8_2 .C_ON=1'b0;
    defparam \tok.uart.valid_54_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \tok.uart.valid_54_LC_6_8_2 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \tok.uart.valid_54_LC_6_8_2  (
            .in0(N__29259),
            .in1(N__19299),
            .in2(_gnd_net_),
            .in3(N__27805),
            .lcout(\tok.uart_rx_valid ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26245),
            .ce(N__14972),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i2_1_lut_LC_6_8_3 .C_ON=1'b0;
    defparam \tok.inv_106_i2_1_lut_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i2_1_lut_LC_6_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i2_1_lut_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24118),
            .lcout(\tok.n301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_99_i6_3_lut_LC_6_8_4 .C_ON=1'b0;
    defparam \tok.or_99_i6_3_lut_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i6_3_lut_LC_6_8_4 .LUT_INIT=16'b1111111101011010;
    LogicCell40 \tok.or_99_i6_3_lut_LC_6_8_4  (
            .in0(N__29027),
            .in1(_gnd_net_),
            .in2(N__28700),
            .in3(N__24140),
            .lcout(\tok.n184 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_142_i15_2_lut_LC_6_8_5 .C_ON=1'b0;
    defparam \tok.equal_142_i15_2_lut_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.equal_142_i15_2_lut_LC_6_8_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \tok.equal_142_i15_2_lut_LC_6_8_5  (
            .in0(_gnd_net_),
            .in1(N__28692),
            .in2(_gnd_net_),
            .in3(N__29025),
            .lcout(),
            .ltout(\tok.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.i3_4_lut_adj_27_LC_6_8_6 .C_ON=1'b0;
    defparam \tok.uart.i3_4_lut_adj_27_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.uart.i3_4_lut_adj_27_LC_6_8_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.uart.i3_4_lut_adj_27_LC_6_8_6  (
            .in0(N__30135),
            .in1(N__29848),
            .in2(N__15236),
            .in3(N__28528),
            .lcout(\tok.n880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_99_i7_3_lut_4_lut_LC_6_8_7 .C_ON=1'b0;
    defparam \tok.or_99_i7_3_lut_4_lut_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i7_3_lut_4_lut_LC_6_8_7 .LUT_INIT=16'b1111100111110101;
    LogicCell40 \tok.or_99_i7_3_lut_4_lut_LC_6_8_7  (
            .in0(N__28529),
            .in1(N__28693),
            .in2(N__21971),
            .in3(N__29026),
            .lcout(\tok.n183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_117_LC_6_9_0 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_117_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_117_LC_6_9_0 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \tok.i4_4_lut_adj_117_LC_6_9_0  (
            .in0(N__21866),
            .in1(N__24473),
            .in2(N__15233),
            .in3(N__26790),
            .lcout(),
            .ltout(\tok.n16_adj_778_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_4_lut_adj_119_LC_6_9_1 .C_ON=1'b0;
    defparam \tok.i8_4_lut_adj_119_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i8_4_lut_adj_119_LC_6_9_1 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \tok.i8_4_lut_adj_119_LC_6_9_1  (
            .in0(N__15220),
            .in1(N__27209),
            .in2(N__15194),
            .in3(N__15191),
            .lcout(\tok.n20_adj_781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_0_i1_2_lut_LC_6_9_2 .C_ON=1'b0;
    defparam \tok.select_73_Select_0_i1_2_lut_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_0_i1_2_lut_LC_6_9_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \tok.select_73_Select_0_i1_2_lut_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__26789),
            .in2(_gnd_net_),
            .in3(N__30148),
            .lcout(\tok.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4624_4_lut_LC_6_9_3 .C_ON=1'b0;
    defparam \tok.i4624_4_lut_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4624_4_lut_LC_6_9_3 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \tok.i4624_4_lut_LC_6_9_3  (
            .in0(N__20588),
            .in1(N__27211),
            .in2(N__15179),
            .in3(N__29411),
            .lcout(\tok.n4664 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_adj_46_LC_6_9_4 .C_ON=1'b0;
    defparam \tok.i3_3_lut_adj_46_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_adj_46_LC_6_9_4 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \tok.i3_3_lut_adj_46_LC_6_9_4  (
            .in0(N__27208),
            .in1(N__20882),
            .in2(_gnd_net_),
            .in3(N__15167),
            .lcout(),
            .ltout(\tok.n14_adj_669_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_48_LC_6_9_5 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_48_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_48_LC_6_9_5 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \tok.i7_4_lut_adj_48_LC_6_9_5  (
            .in0(N__27063),
            .in1(N__15155),
            .in2(N__15149),
            .in3(N__21957),
            .lcout(\tok.n18_adj_672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_LC_6_9_7 .C_ON=1'b0;
    defparam \tok.i5_3_lut_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_LC_6_9_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \tok.i5_3_lut_LC_6_9_7  (
            .in0(N__15146),
            .in1(N__27210),
            .in2(_gnd_net_),
            .in3(N__20774),
            .lcout(\tok.n16_adj_691 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i9_LC_6_10_0 .C_ON=1'b0;
    defparam \tok.A_i9_LC_6_10_0 .SEQ_MODE=4'b1010;
    defparam \tok.A_i9_LC_6_10_0 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \tok.A_i9_LC_6_10_0  (
            .in0(N__17499),
            .in1(N__17370),
            .in2(N__19571),
            .in3(N__17936),
            .lcout(\tok.n60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26255),
            .ce(N__17252),
            .sr(N__19118));
    defparam \tok.A_i16_LC_6_10_1 .C_ON=1'b0;
    defparam \tok.A_i16_LC_6_10_1 .SEQ_MODE=4'b1010;
    defparam \tok.A_i16_LC_6_10_1 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \tok.A_i16_LC_6_10_1  (
            .in0(N__20368),
            .in1(N__17500),
            .in2(N__17385),
            .in3(N__15305),
            .lcout(\tok.n53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26255),
            .ce(N__17252),
            .sr(N__19118));
    defparam \tok.A_i12_LC_6_10_2 .C_ON=1'b0;
    defparam \tok.A_i12_LC_6_10_2 .SEQ_MODE=4'b1010;
    defparam \tok.A_i12_LC_6_10_2 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \tok.A_i12_LC_6_10_2  (
            .in0(N__17498),
            .in1(N__17369),
            .in2(N__20868),
            .in3(N__15299),
            .lcout(\tok.n57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26255),
            .ce(N__17252),
            .sr(N__19118));
    defparam \tok.i9_4_lut_adj_50_LC_6_10_3 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_50_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_50_LC_6_10_3 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i9_4_lut_adj_50_LC_6_10_3  (
            .in0(N__24729),
            .in1(N__15242),
            .in2(N__15293),
            .in3(N__22373),
            .lcout(),
            .ltout(\tok.n20_adj_674_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4674_4_lut_LC_6_10_4 .C_ON=1'b0;
    defparam \tok.i4674_4_lut_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4674_4_lut_LC_6_10_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \tok.i4674_4_lut_LC_6_10_4  (
            .in0(N__15248),
            .in1(N__15284),
            .in2(N__15272),
            .in3(N__15269),
            .lcout(),
            .ltout(\tok.n4676_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i11_LC_6_10_5 .C_ON=1'b0;
    defparam \tok.A_i11_LC_6_10_5 .SEQ_MODE=4'b1010;
    defparam \tok.A_i11_LC_6_10_5 .LUT_INIT=16'b1110010011101110;
    LogicCell40 \tok.A_i11_LC_6_10_5  (
            .in0(N__17368),
            .in1(N__20954),
            .in2(N__15257),
            .in3(N__17501),
            .lcout(\tok.n58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26255),
            .ce(N__17252),
            .sr(N__19118));
    defparam \tok.i1_4_lut_adj_91_LC_6_10_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_91_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_91_LC_6_10_6 .LUT_INIT=16'b1010101100000011;
    LogicCell40 \tok.i1_4_lut_adj_91_LC_6_10_6  (
            .in0(N__21032),
            .in1(N__26622),
            .in2(N__20287),
            .in3(N__24728),
            .lcout(\tok.n12_adj_744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4371_2_lut_LC_6_10_7 .C_ON=1'b0;
    defparam \tok.i4371_2_lut_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i4371_2_lut_LC_6_10_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i4371_2_lut_LC_6_10_7  (
            .in0(N__26623),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21033),
            .lcout(\tok.n4524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_47_LC_6_11_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_47_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_47_LC_6_11_0 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i1_4_lut_adj_47_LC_6_11_0  (
            .in0(N__26804),
            .in1(N__21031),
            .in2(N__28148),
            .in3(N__17908),
            .lcout(\tok.n12_adj_670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_14_i2_3_lut_LC_6_11_1 .C_ON=1'b0;
    defparam \tok.select_73_Select_14_i2_3_lut_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_14_i2_3_lut_LC_6_11_1 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \tok.select_73_Select_14_i2_3_lut_LC_6_11_1  (
            .in0(N__21029),
            .in1(N__22720),
            .in2(_gnd_net_),
            .in3(N__24485),
            .lcout(),
            .ltout(\tok.n2_adj_720_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_76_LC_6_11_2 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_76_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_76_LC_6_11_2 .LUT_INIT=16'b1111010111110001;
    LogicCell40 \tok.i3_4_lut_adj_76_LC_6_11_2  (
            .in0(N__26803),
            .in1(N__28325),
            .in2(N__15404),
            .in3(N__21030),
            .lcout(\tok.n14_adj_722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_79_LC_6_11_4 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_79_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_79_LC_6_11_4 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \tok.i2_4_lut_adj_79_LC_6_11_4  (
            .in0(N__23984),
            .in1(N__28264),
            .in2(N__27071),
            .in3(N__17909),
            .lcout(),
            .ltout(\tok.n13_adj_726_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_83_LC_6_11_5 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_83_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_83_LC_6_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_83_LC_6_11_5  (
            .in0(N__15401),
            .in1(N__15395),
            .in2(N__15383),
            .in3(N__15380),
            .lcout(),
            .ltout(\tok.n20_adj_732_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4671_4_lut_LC_6_11_6 .C_ON=1'b0;
    defparam \tok.i4671_4_lut_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i4671_4_lut_LC_6_11_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i4671_4_lut_LC_6_11_6  (
            .in0(N__15371),
            .in1(N__17132),
            .in2(N__15359),
            .in3(N__15347),
            .lcout(\tok.n4658 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_14_i9_2_lut_LC_6_11_7 .C_ON=1'b0;
    defparam \tok.select_73_Select_14_i9_2_lut_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_14_i9_2_lut_LC_6_11_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \tok.select_73_Select_14_i9_2_lut_LC_6_11_7  (
            .in0(N__20509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29440),
            .lcout(\tok.n9_adj_728 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_142_LC_6_12_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_142_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_142_LC_6_12_1 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \tok.i1_4_lut_adj_142_LC_6_12_1  (
            .in0(N__15341),
            .in1(N__27057),
            .in2(N__15329),
            .in3(N__26813),
            .lcout(),
            .ltout(\tok.n12_adj_815_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_146_LC_6_12_2 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_146_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_146_LC_6_12_2 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \tok.i9_4_lut_adj_146_LC_6_12_2  (
            .in0(N__24073),
            .in1(N__20641),
            .in2(N__15308),
            .in3(N__16292),
            .lcout(),
            .ltout(\tok.n20_adj_822_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_151_LC_6_12_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_151_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_151_LC_6_12_3 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.i1_4_lut_adj_151_LC_6_12_3  (
            .in0(N__15467),
            .in1(N__17497),
            .in2(N__15458),
            .in3(N__16286),
            .lcout(\tok.A_15_N_113_5 ),
            .ltout(\tok.A_15_N_113_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A__15__I_16_i6_3_lut_LC_6_12_4 .C_ON=1'b0;
    defparam \tok.A__15__I_16_i6_3_lut_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.A__15__I_16_i6_3_lut_LC_6_12_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \tok.A__15__I_16_i6_3_lut_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(N__22334),
            .in2(N__15455),
            .in3(N__17749),
            .lcout(\tok.A_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_LC_6_12_5 .C_ON=1'b0;
    defparam \tok.i5_4_lut_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_LC_6_12_5 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i5_4_lut_LC_6_12_5  (
            .in0(N__24491),
            .in1(N__19570),
            .in2(N__15440),
            .in3(N__29445),
            .lcout(\tok.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i6_1_lut_LC_6_12_6 .C_ON=1'b0;
    defparam \tok.inv_106_i6_1_lut_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i6_1_lut_LC_6_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i6_1_lut_LC_6_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22333),
            .lcout(\tok.n297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_101_i9_2_lut_LC_6_12_7 .C_ON=1'b0;
    defparam \tok.or_101_i9_2_lut_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.or_101_i9_2_lut_LC_6_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.or_101_i9_2_lut_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(N__22721),
            .in2(_gnd_net_),
            .in3(N__27428),
            .lcout(\tok.n208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_204_LC_6_13_0 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_204_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_204_LC_6_13_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \tok.i4_4_lut_adj_204_LC_6_13_0  (
            .in0(N__21832),
            .in1(N__21538),
            .in2(N__19949),
            .in3(N__22332),
            .lcout(\tok.n20_adj_858 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i4_1_lut_LC_6_13_1 .C_ON=1'b0;
    defparam \tok.inv_106_i4_1_lut_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i4_1_lut_LC_6_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i4_1_lut_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21831),
            .lcout(\tok.n299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_30_LC_6_13_4 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_30_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_30_LC_6_13_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \tok.i50_4_lut_adj_30_LC_6_13_4  (
            .in0(N__22528),
            .in1(N__19817),
            .in2(N__22277),
            .in3(N__17999),
            .lcout(),
            .ltout(\tok.n27_adj_644_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i7_LC_6_13_5 .C_ON=1'b0;
    defparam \tok.idx_i7_LC_6_13_5 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i7_LC_6_13_5 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.idx_i7_LC_6_13_5  (
            .in0(N__19280),
            .in1(N__18037),
            .in2(N__15407),
            .in3(N__18974),
            .lcout(\tok.n39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26266),
            .ce(),
            .sr(N__19096));
    defparam \tok.idx_i5_LC_6_13_6 .C_ON=1'b0;
    defparam \tok.idx_i5_LC_6_13_6 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i5_LC_6_13_6 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \tok.idx_i5_LC_6_13_6  (
            .in0(N__18973),
            .in1(N__19279),
            .in2(N__18114),
            .in3(N__22190),
            .lcout(\tok.n44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26266),
            .ce(),
            .sr(N__19096));
    defparam \tok.C_stk.tail_i0_i9_LC_7_2_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i9_LC_7_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i9_LC_7_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i9_LC_7_2_0  (
            .in0(N__15545),
            .in1(N__16822),
            .in2(_gnd_net_),
            .in3(N__25588),
            .lcout(\tok.tail_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26218),
            .ce(N__25426),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i1_LC_7_2_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i1_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i1_LC_7_2_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i1_LC_7_2_1  (
            .in0(N__25581),
            .in1(N__15554),
            .in2(_gnd_net_),
            .in3(N__16805),
            .lcout(\tok.C_stk.tail_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26218),
            .ce(N__25426),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i17_LC_7_2_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i17_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i17_LC_7_2_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i17_LC_7_2_2  (
            .in0(N__15553),
            .in1(_gnd_net_),
            .in2(N__15536),
            .in3(N__25585),
            .lcout(\tok.C_stk.tail_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26218),
            .ce(N__25426),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i25_LC_7_2_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i25_LC_7_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i25_LC_7_2_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.C_stk.tail_i0_i25_LC_7_2_3  (
            .in0(N__25582),
            .in1(N__15544),
            .in2(_gnd_net_),
            .in3(N__15521),
            .lcout(\tok.tail_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26218),
            .ce(N__25426),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i33_LC_7_2_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i33_LC_7_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i33_LC_7_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i33_LC_7_2_4  (
            .in0(N__15532),
            .in1(N__15500),
            .in2(_gnd_net_),
            .in3(N__25586),
            .lcout(\tok.C_stk.tail_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26218),
            .ce(N__25426),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i41_LC_7_2_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i41_LC_7_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i41_LC_7_2_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i41_LC_7_2_5  (
            .in0(N__25583),
            .in1(N__15490),
            .in2(_gnd_net_),
            .in3(N__15520),
            .lcout(\tok.tail_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26218),
            .ce(N__25426),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i49_LC_7_2_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i49_LC_7_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i49_LC_7_2_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i49_LC_7_2_6  (
            .in0(N__15511),
            .in1(N__15499),
            .in2(_gnd_net_),
            .in3(N__25587),
            .lcout(\tok.tail_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26218),
            .ce(N__25426),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i50_LC_7_2_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i50_LC_7_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i50_LC_7_2_7 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \tok.C_stk.tail_i0_i50_LC_7_2_7  (
            .in0(N__25584),
            .in1(N__15479),
            .in2(N__16550),
            .in3(_gnd_net_),
            .lcout(\tok.tail_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26218),
            .ce(N__25426),
            .sr(_gnd_net_));
    defparam \tok.i2559_2_lut_4_lut_LC_7_3_0 .C_ON=1'b0;
    defparam \tok.i2559_2_lut_4_lut_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2559_2_lut_4_lut_LC_7_3_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \tok.i2559_2_lut_4_lut_LC_7_3_0  (
            .in0(N__16616),
            .in1(N__15598),
            .in2(N__16685),
            .in3(N__15578),
            .lcout(\tok.C_stk_delta_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_135_LC_7_3_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_135_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_135_LC_7_3_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_135_LC_7_3_1  (
            .in0(_gnd_net_),
            .in1(N__16049),
            .in2(_gnd_net_),
            .in3(N__15817),
            .lcout(\tok.n875 ),
            .ltout(\tok.n875_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2510_2_lut_3_lut_4_lut_LC_7_3_2 .C_ON=1'b0;
    defparam \tok.i2510_2_lut_3_lut_4_lut_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2510_2_lut_3_lut_4_lut_LC_7_3_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i2510_2_lut_3_lut_4_lut_LC_7_3_2  (
            .in0(N__22521),
            .in1(N__15784),
            .in2(N__15602),
            .in3(N__15895),
            .lcout(\tok.n2562 ),
            .ltout(\tok.n2562_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i568_2_lut_4_lut_LC_7_3_3 .C_ON=1'b0;
    defparam \tok.i568_2_lut_4_lut_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \tok.i568_2_lut_4_lut_LC_7_3_3 .LUT_INIT=16'b0101110101010101;
    LogicCell40 \tok.i568_2_lut_4_lut_LC_7_3_3  (
            .in0(N__15577),
            .in1(N__16680),
            .in2(N__15569),
            .in3(N__16615),
            .lcout(\tok.rd_7__N_374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4325_2_lut_LC_7_3_4 .C_ON=1'b0;
    defparam \tok.i4325_2_lut_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4325_2_lut_LC_7_3_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i4325_2_lut_LC_7_3_4  (
            .in0(N__15818),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15897),
            .lcout(),
            .ltout(\tok.n4474_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_115_LC_7_3_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_115_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_115_LC_7_3_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \tok.i1_4_lut_adj_115_LC_7_3_5  (
            .in0(N__15786),
            .in1(N__16681),
            .in2(N__15566),
            .in3(N__16050),
            .lcout(\tok.n802 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_142_i20_2_lut_LC_7_3_6 .C_ON=1'b0;
    defparam \tok.equal_142_i20_2_lut_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.equal_142_i20_2_lut_LC_7_3_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.equal_142_i20_2_lut_LC_7_3_6  (
            .in0(_gnd_net_),
            .in1(N__15785),
            .in2(_gnd_net_),
            .in3(N__15896),
            .lcout(),
            .ltout(\tok.n20_adj_772_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_113_LC_7_3_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_113_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_113_LC_7_3_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i1_4_lut_adj_113_LC_7_3_7  (
            .in0(N__15563),
            .in1(N__28829),
            .in2(N__15557),
            .in3(N__28017),
            .lcout(\tok.n4446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_i3_LC_7_4_0 .C_ON=1'b0;
    defparam \tok.depth_i3_LC_7_4_0 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i3_LC_7_4_0 .LUT_INIT=16'b1011110101000010;
    LogicCell40 \tok.depth_i3_LC_7_4_0  (
            .in0(N__15911),
            .in1(N__15860),
            .in2(N__15899),
            .in3(N__15788),
            .lcout(\tok.n61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26230),
            .ce(),
            .sr(N__19131));
    defparam \tok.depth_i1_LC_7_4_1 .C_ON=1'b0;
    defparam \tok.depth_i1_LC_7_4_1 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i1_LC_7_4_1 .LUT_INIT=16'b1001011011110000;
    LogicCell40 \tok.depth_i1_LC_7_4_1  (
            .in0(N__16048),
            .in1(N__15943),
            .in2(N__15823),
            .in3(N__16008),
            .lcout(\tok.n63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26230),
            .ce(),
            .sr(N__19131));
    defparam \tok.i2_4_lut_4_lut_LC_7_4_2 .C_ON=1'b0;
    defparam \tok.i2_4_lut_4_lut_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_4_lut_LC_7_4_2 .LUT_INIT=16'b1001011011110000;
    LogicCell40 \tok.i2_4_lut_4_lut_LC_7_4_2  (
            .in0(N__15942),
            .in1(N__16047),
            .in2(N__15824),
            .in3(N__16002),
            .lcout(\tok.depth_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_4_lut_LC_7_4_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_4_lut_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_4_lut_LC_7_4_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i1_2_lut_4_lut_LC_7_4_3  (
            .in0(N__15813),
            .in1(N__15783),
            .in2(N__16052),
            .in3(N__15889),
            .lcout(\tok.A_stk_delta_1__N_4 ),
            .ltout(\tok.A_stk_delta_1__N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_LC_7_4_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_LC_7_4_4 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \tok.i1_4_lut_4_lut_LC_7_4_4  (
            .in0(N__15819),
            .in1(N__16046),
            .in2(N__15791),
            .in3(N__16001),
            .lcout(\tok.n4_adj_809 ),
            .ltout(\tok.n4_adj_809_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_196_LC_7_4_5 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_196_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_196_LC_7_4_5 .LUT_INIT=16'b1010100101101010;
    LogicCell40 \tok.i2_4_lut_adj_196_LC_7_4_5  (
            .in0(N__15787),
            .in1(N__15890),
            .in2(N__15761),
            .in3(N__15909),
            .lcout(),
            .ltout(\tok.depth_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_197_LC_7_4_6 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_197_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_197_LC_7_4_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \tok.i1_2_lut_adj_197_LC_7_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15758),
            .in3(N__15755),
            .lcout(\tok.n6_adj_853 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_i2_LC_7_4_7 .C_ON=1'b0;
    defparam \tok.depth_i2_LC_7_4_7 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i2_LC_7_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \tok.depth_i2_LC_7_4_7  (
            .in0(N__15859),
            .in1(N__15894),
            .in2(_gnd_net_),
            .in3(N__15910),
            .lcout(\tok.n62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26230),
            .ce(),
            .sr(N__19131));
    defparam \tok.i4353_2_lut_3_lut_LC_7_5_0 .C_ON=1'b0;
    defparam \tok.i4353_2_lut_3_lut_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4353_2_lut_3_lut_LC_7_5_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i4353_2_lut_3_lut_LC_7_5_0  (
            .in0(N__22492),
            .in1(N__28812),
            .in2(_gnd_net_),
            .in3(N__28512),
            .lcout(\tok.n4504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4400_2_lut_4_lut_LC_7_5_1 .C_ON=1'b0;
    defparam \tok.i4400_2_lut_4_lut_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.i4400_2_lut_4_lut_LC_7_5_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i4400_2_lut_4_lut_LC_7_5_1  (
            .in0(N__28513),
            .in1(N__22493),
            .in2(N__28831),
            .in3(N__15940),
            .lcout(),
            .ltout(\tok.n4554_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_164_LC_7_5_2 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_164_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_164_LC_7_5_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \tok.i5_4_lut_adj_164_LC_7_5_2  (
            .in0(N__27993),
            .in1(N__27311),
            .in2(N__15749),
            .in3(N__15962),
            .lcout(\tok.n237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_161_LC_7_5_3 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_161_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_161_LC_7_5_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.i1_2_lut_adj_161_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(N__28662),
            .in2(_gnd_net_),
            .in3(N__28972),
            .lcout(\tok.n6_adj_832 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_194_LC_7_5_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_194_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_194_LC_7_5_4 .LUT_INIT=16'b0010000000000010;
    LogicCell40 \tok.i1_4_lut_adj_194_LC_7_5_4  (
            .in0(N__27992),
            .in1(N__30394),
            .in2(N__15944),
            .in3(N__30137),
            .lcout(),
            .ltout(\tok.n4432_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_195_LC_7_5_5 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_195_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_195_LC_7_5_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \tok.i4_4_lut_adj_195_LC_7_5_5  (
            .in0(N__15961),
            .in1(N__15953),
            .in2(N__15947),
            .in3(N__29852),
            .lcout(\tok.n1_adj_802 ),
            .ltout(\tok.n1_adj_802_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2578_2_lut_LC_7_5_6 .C_ON=1'b0;
    defparam \tok.i2578_2_lut_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i2578_2_lut_LC_7_5_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \tok.i2578_2_lut_LC_7_5_6  (
            .in0(N__15939),
            .in1(_gnd_net_),
            .in2(N__15914),
            .in3(_gnd_net_),
            .lcout(\tok.n189 ),
            .ltout(\tok.n189_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_192_LC_7_5_7 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_192_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_192_LC_7_5_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \tok.i2_3_lut_adj_192_LC_7_5_7  (
            .in0(N__15898),
            .in1(_gnd_net_),
            .in2(N__15863),
            .in3(N__15858),
            .lcout(\tok.depth_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i11_4_lut_adj_128_LC_7_6_0 .C_ON=1'b0;
    defparam \tok.i11_4_lut_adj_128_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.i11_4_lut_adj_128_LC_7_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i11_4_lut_adj_128_LC_7_6_0  (
            .in0(N__22996),
            .in1(N__21937),
            .in2(N__19825),
            .in3(N__21054),
            .lcout(),
            .ltout(\tok.n27_adj_793_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i15_4_lut_LC_7_6_1 .C_ON=1'b0;
    defparam \tok.i15_4_lut_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i15_4_lut_LC_7_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i15_4_lut_LC_7_6_1  (
            .in0(N__15836),
            .in1(N__15830),
            .in2(N__15845),
            .in3(N__15842),
            .lcout(\tok.tc__7__N_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_129_LC_7_6_2 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_129_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_129_LC_7_6_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i9_4_lut_adj_129_LC_7_6_2  (
            .in0(N__24129),
            .in1(N__28254),
            .in2(N__27446),
            .in3(N__26927),
            .lcout(\tok.n25_adj_794 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_127_LC_7_6_3 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_127_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_127_LC_7_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i10_4_lut_adj_127_LC_7_6_3  (
            .in0(N__22366),
            .in1(N__21839),
            .in2(N__24847),
            .in3(N__20678),
            .lcout(\tok.n26_adj_792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i12_4_lut_adj_126_LC_7_6_4 .C_ON=1'b0;
    defparam \tok.i12_4_lut_adj_126_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i12_4_lut_adj_126_LC_7_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i12_4_lut_adj_126_LC_7_6_4  (
            .in0(N__24013),
            .in1(N__22655),
            .in2(N__20309),
            .in3(N__21428),
            .lcout(\tok.n28_adj_791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_205_LC_7_6_5 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_205_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_205_LC_7_6_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i2_4_lut_adj_205_LC_7_6_5  (
            .in0(N__20143),
            .in1(N__27433),
            .in2(N__24368),
            .in3(N__24130),
            .lcout(\tok.n18_adj_859 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_201_LC_7_7_0 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_201_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_201_LC_7_7_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i6_4_lut_adj_201_LC_7_7_0  (
            .in0(N__20042),
            .in1(N__19813),
            .in2(N__19660),
            .in3(N__21938),
            .lcout(\tok.n22_adj_855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i3_LC_7_7_1 .C_ON=1'b0;
    defparam \tok.A_i3_LC_7_7_1 .SEQ_MODE=4'b1010;
    defparam \tok.A_i3_LC_7_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_i3_LC_7_7_1  (
            .in0(N__17344),
            .in1(N__20043),
            .in2(_gnd_net_),
            .in3(N__16856),
            .lcout(\tok.A_low_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26246),
            .ce(N__17268),
            .sr(N__19142));
    defparam \tok.i2_3_lut_LC_7_7_2 .C_ON=1'b0;
    defparam \tok.i2_3_lut_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_LC_7_7_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i2_3_lut_LC_7_7_2  (
            .in0(N__16075),
            .in1(N__16520),
            .in2(_gnd_net_),
            .in3(N__30411),
            .lcout(\tok.n23 ),
            .ltout(\tok.n23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i2_LC_7_7_3 .C_ON=1'b0;
    defparam \tok.A_i2_LC_7_7_3 .SEQ_MODE=4'b1010;
    defparam \tok.A_i2_LC_7_7_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \tok.A_i2_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__20155),
            .in2(N__16061),
            .in3(N__16127),
            .lcout(\tok.A_low_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26246),
            .ce(N__17268),
            .sr(N__19142));
    defparam \tok.i7_4_lut_adj_202_LC_7_7_7 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_202_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_202_LC_7_7_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \tok.i7_4_lut_adj_202_LC_7_7_7  (
            .in0(N__20857),
            .in1(N__24008),
            .in2(N__20508),
            .in3(N__21410),
            .lcout(\tok.n23_adj_856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.depth_i0_LC_7_8_0 .C_ON=1'b0;
    defparam \tok.depth_i0_LC_7_8_0 .SEQ_MODE=4'b1010;
    defparam \tok.depth_i0_LC_7_8_0 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \tok.depth_i0_LC_7_8_0  (
            .in0(N__16010),
            .in1(_gnd_net_),
            .in2(N__16051),
            .in3(_gnd_net_),
            .lcout(\tok.n64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26250),
            .ce(),
            .sr(N__19114));
    defparam \tok.i1_2_lut_adj_193_LC_7_8_1 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_193_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_193_LC_7_8_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.i1_2_lut_adj_193_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__16039),
            .in2(_gnd_net_),
            .in3(N__16009),
            .lcout(),
            .ltout(\tok.depth_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_199_LC_7_8_2 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_199_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_199_LC_7_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i4_4_lut_adj_199_LC_7_8_2  (
            .in0(N__22503),
            .in1(N__15983),
            .in2(N__15974),
            .in3(N__15971),
            .lcout(\tok.A__15__N_129 ),
            .ltout(\tok.A__15__N_129_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A__15__I_16_i3_3_lut_LC_7_8_3 .C_ON=1'b0;
    defparam \tok.A__15__I_16_i3_3_lut_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.A__15__I_16_i3_3_lut_LC_7_8_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \tok.A__15__I_16_i3_3_lut_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__21942),
            .in2(N__16112),
            .in3(N__16855),
            .lcout(\tok.A_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_214_LC_7_8_4 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_214_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_214_LC_7_8_4 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \tok.i50_4_lut_adj_214_LC_7_8_4  (
            .in0(N__21823),
            .in1(N__22237),
            .in2(N__22522),
            .in3(N__18236),
            .lcout(\tok.n27_adj_866 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.search_clk_198_LC_7_8_5 .C_ON=1'b0;
    defparam \tok.search_clk_198_LC_7_8_5 .SEQ_MODE=4'b1010;
    defparam \tok.search_clk_198_LC_7_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \tok.search_clk_198_LC_7_8_5  (
            .in0(N__22239),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.search_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26250),
            .ce(),
            .sr(N__19114));
    defparam \tok.i50_4_lut_adj_216_LC_7_8_6 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_216_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_216_LC_7_8_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \tok.i50_4_lut_adj_216_LC_7_8_6  (
            .in0(N__22507),
            .in1(N__22238),
            .in2(N__18155),
            .in3(N__27429),
            .lcout(),
            .ltout(\tok.n27_adj_867_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i4_LC_7_8_7 .C_ON=1'b0;
    defparam \tok.idx_i4_LC_7_8_7 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i4_LC_7_8_7 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.idx_i4_LC_7_8_7  (
            .in0(N__19260),
            .in1(N__18174),
            .in2(N__16109),
            .in3(N__18954),
            .lcout(\tok.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26250),
            .ce(),
            .sr(N__19114));
    defparam \tok.i4390_2_lut_LC_7_9_0 .C_ON=1'b0;
    defparam \tok.i4390_2_lut_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4390_2_lut_LC_7_9_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \tok.i4390_2_lut_LC_7_9_0  (
            .in0(N__30150),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24705),
            .lcout(\tok.n4544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_2_lut_LC_7_9_1 .C_ON=1'b0;
    defparam \tok.sub_100_add_2_2_lut_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_2_lut_LC_7_9_1 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \tok.sub_100_add_2_2_lut_LC_7_9_1  (
            .in0(N__21685),
            .in1(N__22181),
            .in2(_gnd_net_),
            .in3(N__30149),
            .lcout(\tok.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_52_LC_7_9_2 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_52_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_52_LC_7_9_2 .LUT_INIT=16'b1111000111111011;
    LogicCell40 \tok.i2_4_lut_adj_52_LC_7_9_2  (
            .in0(N__26925),
            .in1(N__26604),
            .in2(N__16106),
            .in3(N__17904),
            .lcout(),
            .ltout(\tok.n14_adj_678_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_54_LC_7_9_3 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_54_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_54_LC_7_9_3 .LUT_INIT=16'b1111001011111111;
    LogicCell40 \tok.i7_4_lut_adj_54_LC_7_9_3  (
            .in0(N__17155),
            .in1(N__27062),
            .in2(N__16097),
            .in3(N__17509),
            .lcout(),
            .ltout(\tok.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_LC_7_9_4 .C_ON=1'b0;
    defparam \tok.i10_4_lut_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_LC_7_9_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i10_4_lut_LC_7_9_4  (
            .in0(N__18929),
            .in1(N__16169),
            .in2(N__16163),
            .in3(N__29342),
            .lcout(),
            .ltout(\tok.n22_adj_683_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i11_4_lut_LC_7_9_5 .C_ON=1'b0;
    defparam \tok.i11_4_lut_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i11_4_lut_LC_7_9_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i11_4_lut_LC_7_9_5  (
            .in0(N__16160),
            .in1(N__24200),
            .in2(N__16148),
            .in3(N__16145),
            .lcout(\tok.A_15_N_113_0 ),
            .ltout(\tok.A_15_N_113_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A__15__I_16_i1_3_lut_LC_7_9_6 .C_ON=1'b0;
    defparam \tok.A__15__I_16_i1_3_lut_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.A__15__I_16_i1_3_lut_LC_7_9_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \tok.A__15__I_16_i1_3_lut_LC_7_9_6  (
            .in0(N__26926),
            .in1(_gnd_net_),
            .in2(N__16139),
            .in3(N__17715),
            .lcout(\tok.A_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_171_LC_7_10_0 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_171_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_171_LC_7_10_0 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \tok.i1_4_lut_adj_171_LC_7_10_0  (
            .in0(N__21449),
            .in1(N__24242),
            .in2(N__17520),
            .in3(N__16136),
            .lcout(\tok.A_15_N_113_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i44_3_lut_LC_7_10_1 .C_ON=1'b0;
    defparam \tok.i44_3_lut_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i44_3_lut_LC_7_10_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.i44_3_lut_LC_7_10_1  (
            .in0(N__21795),
            .in1(N__26618),
            .in2(_gnd_net_),
            .in3(N__17890),
            .lcout(\tok.n4520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_3_lut_adj_187_LC_7_10_2 .C_ON=1'b0;
    defparam \tok.i50_3_lut_adj_187_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i50_3_lut_adj_187_LC_7_10_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \tok.i50_3_lut_adj_187_LC_7_10_2  (
            .in0(N__17891),
            .in1(_gnd_net_),
            .in2(N__26624),
            .in3(N__24168),
            .lcout(),
            .ltout(\tok.n46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_188_LC_7_10_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_188_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_188_LC_7_10_3 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \tok.i1_4_lut_adj_188_LC_7_10_3  (
            .in0(N__17534),
            .in1(N__17508),
            .in2(N__16130),
            .in3(N__17573),
            .lcout(\tok.A_15_N_113_1 ),
            .ltout(\tok.A_15_N_113_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A__15__I_16_i2_3_lut_LC_7_10_4 .C_ON=1'b0;
    defparam \tok.A__15__I_16_i2_3_lut_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.A__15__I_16_i2_3_lut_LC_7_10_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \tok.A__15__I_16_i2_3_lut_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__17738),
            .in2(N__16118),
            .in3(N__24169),
            .lcout(),
            .ltout(\tok.A_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i4_LC_7_10_5 .C_ON=1'b0;
    defparam \tok.uart.sender_i4_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i4_LC_7_10_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.uart.sender_i4_LC_7_10_5  (
            .in0(N__16467),
            .in1(_gnd_net_),
            .in2(N__16115),
            .in3(N__16247),
            .lcout(\tok.uart.sender_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26261),
            .ce(N__16388),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i3_LC_7_10_6 .C_ON=1'b0;
    defparam \tok.uart.sender_i3_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i3_LC_7_10_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i3_LC_7_10_6  (
            .in0(N__16280),
            .in1(N__16466),
            .in2(_gnd_net_),
            .in3(N__16274),
            .lcout(sender_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26261),
            .ce(N__16388),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i5_LC_7_10_7 .C_ON=1'b0;
    defparam \tok.uart.sender_i5_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i5_LC_7_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.sender_i5_LC_7_10_7  (
            .in0(N__16468),
            .in1(N__16397),
            .in2(_gnd_net_),
            .in3(N__16256),
            .lcout(\tok.uart.sender_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26261),
            .ce(N__16388),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_118_LC_7_11_0 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_118_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_118_LC_7_11_0 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \tok.i2_3_lut_adj_118_LC_7_11_0  (
            .in0(N__26603),
            .in1(N__28218),
            .in2(_gnd_net_),
            .in3(N__17889),
            .lcout(),
            .ltout(\tok.n14_adj_779_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_121_LC_7_11_1 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_121_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_121_LC_7_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \tok.i10_4_lut_adj_121_LC_7_11_1  (
            .in0(N__16241),
            .in1(N__19841),
            .in2(N__16229),
            .in3(N__16226),
            .lcout(),
            .ltout(\tok.n22_adj_784_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_123_LC_7_11_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_123_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_123_LC_7_11_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.i1_4_lut_adj_123_LC_7_11_2  (
            .in0(N__21233),
            .in1(N__17521),
            .in2(N__16214),
            .in3(N__23909),
            .lcout(\tok.A_15_N_113_6 ),
            .ltout(\tok.A_15_N_113_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A__15__I_16_i7_3_lut_LC_7_11_3 .C_ON=1'b0;
    defparam \tok.A__15__I_16_i7_3_lut_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.A__15__I_16_i7_3_lut_LC_7_11_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \tok.A__15__I_16_i7_3_lut_LC_7_11_3  (
            .in0(N__28219),
            .in1(_gnd_net_),
            .in2(N__16211),
            .in3(N__17748),
            .lcout(),
            .ltout(\tok.A_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i9_LC_7_11_4 .C_ON=1'b0;
    defparam \tok.uart.sender_i9_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i9_LC_7_11_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.uart.sender_i9_LC_7_11_4  (
            .in0(N__16472),
            .in1(_gnd_net_),
            .in2(N__16208),
            .in3(N__16205),
            .lcout(\tok.uart.sender_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26264),
            .ce(N__16387),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i8_LC_7_11_5 .C_ON=1'b0;
    defparam \tok.uart.sender_i8_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i8_LC_7_11_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i8_LC_7_11_5  (
            .in0(N__16187),
            .in1(N__16471),
            .in2(_gnd_net_),
            .in3(N__16181),
            .lcout(\tok.uart.sender_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26264),
            .ce(N__16387),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i7_LC_7_11_6 .C_ON=1'b0;
    defparam \tok.uart.sender_i7_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i7_LC_7_11_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.uart.sender_i7_LC_7_11_6  (
            .in0(N__16470),
            .in1(N__16175),
            .in2(_gnd_net_),
            .in3(N__17528),
            .lcout(\tok.uart.sender_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26264),
            .ce(N__16387),
            .sr(_gnd_net_));
    defparam \tok.uart.sender_i6_LC_7_11_7 .C_ON=1'b0;
    defparam \tok.uart.sender_i6_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.sender_i6_LC_7_11_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.uart.sender_i6_LC_7_11_7  (
            .in0(N__16478),
            .in1(N__16469),
            .in2(_gnd_net_),
            .in3(N__17684),
            .lcout(\tok.uart.sender_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26264),
            .ce(N__16387),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_66_LC_7_12_0 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_66_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_66_LC_7_12_0 .LUT_INIT=16'b0000110001011101;
    LogicCell40 \tok.i2_4_lut_adj_66_LC_7_12_0  (
            .in0(N__26602),
            .in1(N__22349),
            .in2(N__27073),
            .in3(N__20642),
            .lcout(\tok.n14_adj_707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_4_lut_adj_67_LC_7_12_1 .C_ON=1'b0;
    defparam \tok.i8_4_lut_adj_67_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i8_4_lut_adj_67_LC_7_12_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i8_4_lut_adj_67_LC_7_12_1  (
            .in0(N__20643),
            .in1(N__16337),
            .in2(N__22541),
            .in3(N__17881),
            .lcout(),
            .ltout(\tok.n20_adj_708_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i10_4_lut_adj_68_LC_7_12_2 .C_ON=1'b0;
    defparam \tok.i10_4_lut_adj_68_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i10_4_lut_adj_68_LC_7_12_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \tok.i10_4_lut_adj_68_LC_7_12_2  (
            .in0(N__17522),
            .in1(N__16325),
            .in2(N__16319),
            .in3(N__24635),
            .lcout(),
            .ltout(\tok.n22_adj_709_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i14_LC_7_12_3 .C_ON=1'b0;
    defparam \tok.A_i14_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \tok.A_i14_LC_7_12_3 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \tok.A_i14_LC_7_12_3  (
            .in0(N__17378),
            .in1(N__22763),
            .in2(N__16316),
            .in3(N__20597),
            .lcout(\tok.n55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26267),
            .ce(N__17267),
            .sr(N__19066));
    defparam \tok.A_i6_LC_7_12_4 .C_ON=1'b0;
    defparam \tok.A_i6_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \tok.A_i6_LC_7_12_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_i6_LC_7_12_4  (
            .in0(N__19948),
            .in1(N__17379),
            .in2(_gnd_net_),
            .in3(N__16313),
            .lcout(\tok.A_low_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26267),
            .ce(N__17267),
            .sr(N__19066));
    defparam \tok.i2_4_lut_adj_140_LC_7_12_5 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_140_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_140_LC_7_12_5 .LUT_INIT=16'b1010101111111011;
    LogicCell40 \tok.i2_4_lut_adj_140_LC_7_12_5  (
            .in0(N__16307),
            .in1(N__26601),
            .in2(N__22374),
            .in3(N__17880),
            .lcout(),
            .ltout(\tok.n13_adj_813_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_144_LC_7_12_6 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_144_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_144_LC_7_12_6 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i7_4_lut_adj_144_LC_7_12_6  (
            .in0(N__19947),
            .in1(N__22805),
            .in2(N__16295),
            .in3(N__29444),
            .lcout(\tok.n18_adj_819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_149_LC_7_13_0 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_149_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_149_LC_7_13_0 .LUT_INIT=16'b1111010011111000;
    LogicCell40 \tok.i4_4_lut_adj_149_LC_7_13_0  (
            .in0(N__26920),
            .in1(N__24735),
            .in2(N__19862),
            .in3(N__28698),
            .lcout(\tok.n15_adj_823 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_43_LC_7_13_1 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_43_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_43_LC_7_13_1 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \tok.i50_4_lut_adj_43_LC_7_13_1  (
            .in0(N__17759),
            .in1(N__26921),
            .in2(N__22529),
            .in3(N__22272),
            .lcout(\tok.n27_adj_664 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_209_LC_7_13_2 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_209_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_209_LC_7_13_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \tok.i50_4_lut_adj_209_LC_7_13_2  (
            .in0(N__22527),
            .in1(N__18374),
            .in2(N__22282),
            .in3(N__24185),
            .lcout(),
            .ltout(\tok.n27_adj_863_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i1_LC_7_13_3 .C_ON=1'b0;
    defparam \tok.idx_i1_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i1_LC_7_13_3 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.idx_i1_LC_7_13_3  (
            .in0(N__19276),
            .in1(N__18408),
            .in2(N__16502),
            .in3(N__18970),
            .lcout(\tok.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26269),
            .ce(),
            .sr(N__19086));
    defparam \tok.i50_4_lut_adj_212_LC_7_13_4 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_212_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_212_LC_7_13_4 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \tok.i50_4_lut_adj_212_LC_7_13_4  (
            .in0(N__22273),
            .in1(N__22526),
            .in2(N__18308),
            .in3(N__21972),
            .lcout(),
            .ltout(\tok.n27_adj_865_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i2_LC_7_13_5 .C_ON=1'b0;
    defparam \tok.idx_i2_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i2_LC_7_13_5 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.idx_i2_LC_7_13_5  (
            .in0(N__19277),
            .in1(N__18334),
            .in2(N__16499),
            .in3(N__18971),
            .lcout(\tok.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26269),
            .ce(),
            .sr(N__19086));
    defparam \tok.idx_i0_LC_7_13_6 .C_ON=1'b0;
    defparam \tok.idx_i0_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i0_LC_7_13_6 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.idx_i0_LC_7_13_6  (
            .in0(N__18969),
            .in1(N__16496),
            .in2(N__17796),
            .in3(N__19275),
            .lcout(\tok.n52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26269),
            .ce(),
            .sr(N__19086));
    defparam \tok.idx_i3_LC_7_13_7 .C_ON=1'b0;
    defparam \tok.idx_i3_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i3_LC_7_13_7 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \tok.idx_i3_LC_7_13_7  (
            .in0(N__19278),
            .in1(N__18972),
            .in2(N__18273),
            .in3(N__16490),
            .lcout(\tok.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26269),
            .ce(),
            .sr(N__19086));
    defparam \tok.C_stk.tail_i0_i26_LC_8_2_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i26_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i26_LC_8_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i26_LC_8_2_0  (
            .in0(N__16559),
            .in1(N__23323),
            .in2(_gnd_net_),
            .in3(N__25594),
            .lcout(\tok.tail_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26226),
            .ce(N__25427),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i34_LC_8_2_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i34_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i34_LC_8_2_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \tok.C_stk.tail_i0_i34_LC_8_2_1  (
            .in0(N__25590),
            .in1(N__18535),
            .in2(N__16549),
            .in3(_gnd_net_),
            .lcout(\tok.C_stk.tail_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26226),
            .ce(N__25427),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i36_LC_8_2_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i36_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i36_LC_8_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i36_LC_8_2_2  (
            .in0(N__23344),
            .in1(N__16531),
            .in2(_gnd_net_),
            .in3(N__25596),
            .lcout(\tok.C_stk.tail_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26226),
            .ce(N__25427),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i42_LC_8_2_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i42_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i42_LC_8_2_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.C_stk.tail_i0_i42_LC_8_2_3  (
            .in0(N__25592),
            .in1(_gnd_net_),
            .in2(N__16576),
            .in3(N__16558),
            .lcout(\tok.tail_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26226),
            .ce(N__25427),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i20_LC_8_2_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i20_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i20_LC_8_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i20_LC_8_2_4  (
            .in0(N__18523),
            .in1(N__16532),
            .in2(_gnd_net_),
            .in3(N__25593),
            .lcout(\tok.C_stk.tail_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26226),
            .ce(N__25427),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i32_LC_8_2_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i32_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i32_LC_8_2_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i32_LC_8_2_5  (
            .in0(N__25589),
            .in1(N__18482),
            .in2(_gnd_net_),
            .in3(N__23156),
            .lcout(\tok.C_stk.tail_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26226),
            .ce(N__25427),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i28_LC_8_2_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i28_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i28_LC_8_2_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i28_LC_8_2_6  (
            .in0(N__17989),
            .in1(N__18512),
            .in2(_gnd_net_),
            .in3(N__25595),
            .lcout(\tok.tail_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26226),
            .ce(N__25427),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i40_LC_8_2_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i40_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i40_LC_8_2_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i40_LC_8_2_7  (
            .in0(N__25591),
            .in1(N__18460),
            .in2(_gnd_net_),
            .in3(N__23167),
            .lcout(\tok.tail_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26226),
            .ce(N__25427),
            .sr(_gnd_net_));
    defparam \tok.i127_4_lut_4_lut_LC_8_3_0 .C_ON=1'b0;
    defparam \tok.i127_4_lut_4_lut_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.i127_4_lut_4_lut_LC_8_3_0 .LUT_INIT=16'b1011010000111111;
    LogicCell40 \tok.i127_4_lut_4_lut_LC_8_3_0  (
            .in0(N__30445),
            .in1(N__29870),
            .in2(N__28555),
            .in3(N__30157),
            .lcout(),
            .ltout(\tok.n127_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_116_LC_8_3_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_116_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_116_LC_8_3_1 .LUT_INIT=16'b1111010011111110;
    LogicCell40 \tok.i1_4_lut_adj_116_LC_8_3_1  (
            .in0(N__29871),
            .in1(N__25872),
            .in2(N__16523),
            .in3(N__29032),
            .lcout(),
            .ltout(\tok.n4394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_124_LC_8_3_2 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_124_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_124_LC_8_3_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \tok.i3_4_lut_adj_124_LC_8_3_2  (
            .in0(N__16516),
            .in1(N__27310),
            .in2(N__16505),
            .in3(N__28697),
            .lcout(\tok.n86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_2_lut_LC_8_3_3 .C_ON=1'b0;
    defparam \tok.i2_2_lut_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_2_lut_LC_8_3_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i2_2_lut_LC_8_3_3  (
            .in0(N__29872),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30446),
            .lcout(),
            .ltout(\tok.n28_adj_834_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4564_4_lut_LC_8_3_4 .C_ON=1'b0;
    defparam \tok.i4564_4_lut_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4564_4_lut_LC_8_3_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \tok.i4564_4_lut_LC_8_3_4  (
            .in0(N__29033),
            .in1(N__28019),
            .in2(N__16637),
            .in3(N__30159),
            .lcout(),
            .ltout(\tok.n4604_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i49_4_lut_LC_8_3_5 .C_ON=1'b0;
    defparam \tok.i49_4_lut_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.i49_4_lut_LC_8_3_5 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.i49_4_lut_LC_8_3_5  (
            .in0(N__17600),
            .in1(N__29034),
            .in2(N__16634),
            .in3(N__28548),
            .lcout(\tok.n34_adj_719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_LC_8_3_6 .C_ON=1'b0;
    defparam \tok.i125_4_lut_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_LC_8_3_6 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \tok.i125_4_lut_LC_8_3_6  (
            .in0(N__30444),
            .in1(N__18598),
            .in2(N__24233),
            .in3(N__30158),
            .lcout(\tok.n83_adj_704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_125_LC_8_3_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_125_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_125_LC_8_3_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_125_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__29031),
            .in2(_gnd_net_),
            .in3(N__30443),
            .lcout(\tok.n101_adj_776 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4567_4_lut_LC_8_4_0 .C_ON=1'b0;
    defparam \tok.i4567_4_lut_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4567_4_lut_LC_8_4_0 .LUT_INIT=16'b0100100010000000;
    LogicCell40 \tok.i4567_4_lut_LC_8_4_0  (
            .in0(N__29866),
            .in1(N__29008),
            .in2(N__30442),
            .in3(N__30154),
            .lcout(),
            .ltout(\tok.n4610_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i58_4_lut_LC_8_4_1 .C_ON=1'b0;
    defparam \tok.i58_4_lut_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.i58_4_lut_LC_8_4_1 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \tok.i58_4_lut_LC_8_4_1  (
            .in0(N__30155),
            .in1(N__16670),
            .in2(N__16619),
            .in3(N__28530),
            .lcout(\tok.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_131_LC_8_4_2 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_131_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_131_LC_8_4_2 .LUT_INIT=16'b0101000010001000;
    LogicCell40 \tok.i125_4_lut_adj_131_LC_8_4_2  (
            .in0(N__30423),
            .in1(N__16607),
            .in2(N__18744),
            .in3(N__30156),
            .lcout(),
            .ltout(\tok.n83_adj_796_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4604_2_lut_3_lut_LC_8_4_3 .C_ON=1'b0;
    defparam \tok.i4604_2_lut_3_lut_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4604_2_lut_3_lut_LC_8_4_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \tok.i4604_2_lut_3_lut_LC_8_4_3  (
            .in0(N__29009),
            .in1(_gnd_net_),
            .in2(N__16583),
            .in3(N__29867),
            .lcout(\tok.n4602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_133_LC_8_4_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_133_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_133_LC_8_4_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_133_LC_8_4_4  (
            .in0(N__25183),
            .in1(N__18880),
            .in2(N__25259),
            .in3(N__18698),
            .lcout(n92_adj_872),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i2_LC_8_4_5 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i2_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i2_LC_8_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.uart.capture_i0_i2_LC_8_4_5  (
            .in0(N__16975),
            .in1(N__16718),
            .in2(_gnd_net_),
            .in3(N__16964),
            .lcout(capture_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26236),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_adj_73_LC_8_4_6 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_adj_73_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_adj_73_LC_8_4_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \tok.i1_2_lut_3_lut_adj_73_LC_8_4_6  (
            .in0(N__28679),
            .in1(N__28828),
            .in2(_gnd_net_),
            .in3(N__28018),
            .lcout(\tok.n847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i59_3_lut_LC_8_4_7 .C_ON=1'b0;
    defparam \tok.i59_3_lut_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \tok.i59_3_lut_LC_8_4_7 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \tok.i59_3_lut_LC_8_4_7  (
            .in0(N__29007),
            .in1(N__30419),
            .in2(_gnd_net_),
            .in3(N__29865),
            .lcout(\tok.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.n602_bdd_4_lut_4749_LC_8_5_0 .C_ON=1'b0;
    defparam \tok.C_stk.n602_bdd_4_lut_4749_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.n602_bdd_4_lut_4749_LC_8_5_0 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \tok.C_stk.n602_bdd_4_lut_4749_LC_8_5_0  (
            .in0(N__18913),
            .in1(N__25107),
            .in2(N__26358),
            .in3(N__18802),
            .lcout(),
            .ltout(\tok.C_stk.n4906_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i6_LC_8_5_1 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i6_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i6_LC_8_5_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \tok.C_stk.head_i0_i6_LC_8_5_1  (
            .in0(N__24962),
            .in1(N__23098),
            .in2(N__16661),
            .in3(N__26352),
            .lcout(\tok.c_stk_r_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26241),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i4641_4_lut_LC_8_5_2 .C_ON=1'b0;
    defparam \tok.ram.i4641_4_lut_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i4641_4_lut_LC_8_5_2 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \tok.ram.i4641_4_lut_LC_8_5_2  (
            .in0(N__18911),
            .in1(N__26684),
            .in2(N__23106),
            .in3(N__25990),
            .lcout(),
            .ltout(\tok.ram.n4699_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5_4_lut_adj_25_LC_8_5_3 .C_ON=1'b0;
    defparam \tok.ram.i5_4_lut_adj_25_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5_4_lut_adj_25_LC_8_5_3 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.ram.i5_4_lut_adj_25_LC_8_5_3  (
            .in0(N__23099),
            .in1(N__25897),
            .in2(N__16658),
            .in3(N__29855),
            .lcout(),
            .ltout(\tok.n1_adj_760_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_104_LC_8_5_4 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_104_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_104_LC_8_5_4 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i27_4_lut_adj_104_LC_8_5_4  (
            .in0(N__16655),
            .in1(N__28550),
            .in2(N__16643),
            .in3(N__30147),
            .lcout(),
            .ltout(\tok.n13_adj_761_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_106_LC_8_5_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_106_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_106_LC_8_5_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_106_LC_8_5_5  (
            .in0(N__25260),
            .in1(N__25189),
            .in2(N__16640),
            .in3(N__18912),
            .lcout(n92_adj_871),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_LC_8_5_6 .C_ON=1'b0;
    defparam \tok.i26_3_lut_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_LC_8_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.i26_3_lut_LC_8_5_6  (
            .in0(N__18856),
            .in1(N__18840),
            .in2(_gnd_net_),
            .in3(N__23516),
            .lcout(\tok.tc_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.n602_bdd_4_lut_4719_LC_8_6_0 .C_ON=1'b0;
    defparam \tok.C_stk.n602_bdd_4_lut_4719_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.n602_bdd_4_lut_4719_LC_8_6_0 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \tok.C_stk.n602_bdd_4_lut_4719_LC_8_6_0  (
            .in0(N__26345),
            .in1(N__18643),
            .in2(N__25112),
            .in3(N__18765),
            .lcout(),
            .ltout(\tok.C_stk.n4870_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i1_LC_8_6_1 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i1_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i1_LC_8_6_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \tok.C_stk.head_i0_i1_LC_8_6_1  (
            .in0(N__16829),
            .in1(N__16788),
            .in2(N__16811),
            .in3(N__26346),
            .lcout(\tok.c_stk_r_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26247),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i4662_4_lut_LC_8_6_2 .C_ON=1'b0;
    defparam \tok.ram.i4662_4_lut_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i4662_4_lut_LC_8_6_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.ram.i4662_4_lut_LC_8_6_2  (
            .in0(N__26696),
            .in1(N__18641),
            .in2(N__16794),
            .in3(N__25983),
            .lcout(),
            .ltout(\tok.ram.n4714_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5_4_lut_adj_20_LC_8_6_3 .C_ON=1'b0;
    defparam \tok.ram.i5_4_lut_adj_20_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5_4_lut_adj_20_LC_8_6_3 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \tok.ram.i5_4_lut_adj_20_LC_8_6_3  (
            .in0(N__29847),
            .in1(N__25898),
            .in2(N__16808),
            .in3(N__16787),
            .lcout(),
            .ltout(\tok.n1_adj_717_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i18_4_lut_LC_8_6_4 .C_ON=1'b0;
    defparam \tok.i18_4_lut_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i18_4_lut_LC_8_6_4 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \tok.i18_4_lut_LC_8_6_4  (
            .in0(N__28554),
            .in1(N__16766),
            .in2(N__16754),
            .in3(N__30134),
            .lcout(),
            .ltout(\tok.n5_adj_718_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_74_LC_8_6_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_74_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_74_LC_8_6_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_74_LC_8_6_5  (
            .in0(N__18642),
            .in1(N__25261),
            .in2(N__16751),
            .in3(N__25190),
            .lcout(n92),
            .ltout(n92_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_147_LC_8_6_6 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_147_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_147_LC_8_6_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \tok.i26_3_lut_adj_147_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__23498),
            .in2(N__16748),
            .in3(N__18766),
            .lcout(\tok.tc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_182_LC_8_7_0 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_182_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_182_LC_8_7_0 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \tok.i2_4_lut_adj_182_LC_8_7_0  (
            .in0(N__16730),
            .in1(N__27275),
            .in2(N__22658),
            .in3(N__26435),
            .lcout(),
            .ltout(\tok.n6_adj_848_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_183_LC_8_7_1 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_183_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_183_LC_8_7_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i3_4_lut_adj_183_LC_8_7_1  (
            .in0(N__17008),
            .in1(N__17027),
            .in2(N__17015),
            .in3(N__27794),
            .lcout(),
            .ltout(\tok.n32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_184_LC_8_7_2 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_184_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_184_LC_8_7_2 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i3_4_lut_adj_184_LC_8_7_2  (
            .in0(N__29247),
            .in1(N__30410),
            .in2(N__17012),
            .in3(N__24269),
            .lcout(\tok.n10_adj_849 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i1_LC_8_7_3 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i1_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i1_LC_8_7_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.uart.rx_data_i0_i1_LC_8_7_3  (
            .in0(N__17009),
            .in1(_gnd_net_),
            .in2(N__16985),
            .in3(N__22113),
            .lcout(uart_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26251),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1549_3_lut_4_lut_LC_8_7_4 .C_ON=1'b0;
    defparam \tok.i1549_3_lut_4_lut_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1549_3_lut_4_lut_LC_8_7_4 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \tok.i1549_3_lut_4_lut_LC_8_7_4  (
            .in0(N__23867),
            .in1(N__18917),
            .in2(N__29284),
            .in3(N__21320),
            .lcout(\tok.table_wr_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.capture_i0_i1_LC_8_7_6 .C_ON=1'b0;
    defparam \tok.uart.capture_i0_i1_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \tok.uart.capture_i0_i1_LC_8_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.uart.capture_i0_i1_LC_8_7_6  (
            .in0(N__17172),
            .in1(N__16981),
            .in2(_gnd_net_),
            .in3(N__16953),
            .lcout(capture_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26251),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1697_3_lut_4_lut_LC_8_7_7 .C_ON=1'b0;
    defparam \tok.i1697_3_lut_4_lut_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1697_3_lut_4_lut_LC_8_7_7 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \tok.i1697_3_lut_4_lut_LC_8_7_7  (
            .in0(N__20059),
            .in1(N__29251),
            .in2(N__26036),
            .in3(N__23868),
            .lcout(\tok.table_wr_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_176_LC_8_8_0 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_176_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_176_LC_8_8_0 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \tok.i7_4_lut_adj_176_LC_8_8_0  (
            .in0(N__22016),
            .in1(N__29394),
            .in2(N__20069),
            .in3(N__17660),
            .lcout(),
            .ltout(\tok.n18_adj_844_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_180_LC_8_8_1 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_180_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_180_LC_8_8_1 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \tok.i9_4_lut_adj_180_LC_8_8_1  (
            .in0(N__24067),
            .in1(N__17186),
            .in2(N__16874),
            .in3(N__21060),
            .lcout(),
            .ltout(\tok.n20_adj_846_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_181_LC_8_8_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_181_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_181_LC_8_8_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.i1_4_lut_adj_181_LC_8_8_2  (
            .in0(N__16871),
            .in1(N__17488),
            .in2(N__16859),
            .in3(N__17216),
            .lcout(\tok.A_15_N_113_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_3_lut_LC_8_8_3 .C_ON=1'b0;
    defparam \tok.i4_3_lut_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4_3_lut_LC_8_8_3 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \tok.i4_3_lut_LC_8_8_3  (
            .in0(N__29850),
            .in1(_gnd_net_),
            .in2(N__19970),
            .in3(N__24712),
            .lcout(\tok.n15_adj_847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_175_LC_8_8_4 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_175_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_175_LC_8_8_4 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \tok.i1_4_lut_adj_175_LC_8_8_4  (
            .in0(N__27046),
            .in1(N__26791),
            .in2(N__17210),
            .in3(N__29849),
            .lcout(\tok.n12_adj_843 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i0_LC_8_8_5 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i0_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i0_LC_8_8_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.uart.rx_data_i0_i0_LC_8_8_5  (
            .in0(N__17173),
            .in1(N__22122),
            .in2(_gnd_net_),
            .in3(N__17156),
            .lcout(uart_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26256),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_3_lut_adj_82_LC_8_9_0 .C_ON=1'b0;
    defparam \tok.i5_3_lut_adj_82_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i5_3_lut_adj_82_LC_8_9_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \tok.i5_3_lut_adj_82_LC_8_9_0  (
            .in0(N__27217),
            .in1(N__17144),
            .in2(_gnd_net_),
            .in3(N__20411),
            .lcout(\tok.n16_adj_730 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_155_i16_2_lut_3_lut_LC_8_9_1 .C_ON=1'b0;
    defparam \tok.equal_155_i16_2_lut_3_lut_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.equal_155_i16_2_lut_3_lut_LC_8_9_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \tok.equal_155_i16_2_lut_3_lut_LC_8_9_1  (
            .in0(N__28075),
            .in1(N__29221),
            .in2(_gnd_net_),
            .in3(N__28117),
            .lcout(\tok.n400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2649_3_lut_4_lut_LC_8_9_2 .C_ON=1'b0;
    defparam \tok.i2649_3_lut_4_lut_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2649_3_lut_4_lut_LC_8_9_2 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \tok.i2649_3_lut_4_lut_LC_8_9_2  (
            .in0(N__27216),
            .in1(N__17036),
            .in2(N__29267),
            .in3(N__23865),
            .lcout(\tok.n2724 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1771_3_lut_4_lut_LC_8_9_3 .C_ON=1'b0;
    defparam \tok.i1771_3_lut_4_lut_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1771_3_lut_4_lut_LC_8_9_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \tok.i1771_3_lut_4_lut_LC_8_9_3  (
            .in0(N__23866),
            .in1(N__18677),
            .in2(N__29576),
            .in3(N__29226),
            .lcout(\tok.table_wr_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2562_3_lut_4_lut_LC_8_9_4 .C_ON=1'b0;
    defparam \tok.i2562_3_lut_4_lut_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2562_3_lut_4_lut_LC_8_9_4 .LUT_INIT=16'b1011101110110000;
    LogicCell40 \tok.i2562_3_lut_4_lut_LC_8_9_4  (
            .in0(N__24622),
            .in1(N__28076),
            .in2(N__29266),
            .in3(N__26410),
            .lcout(\tok.n2614 ),
            .ltout(\tok.n2614_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2564_3_lut_4_lut_LC_8_9_5 .C_ON=1'b0;
    defparam \tok.i2564_3_lut_4_lut_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2564_3_lut_4_lut_LC_8_9_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \tok.i2564_3_lut_4_lut_LC_8_9_5  (
            .in0(N__28130),
            .in1(N__29222),
            .in2(N__17030),
            .in3(N__28118),
            .lcout(\tok.n2616 ),
            .ltout(\tok.n2616_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_186_LC_8_9_6 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_186_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_186_LC_8_9_6 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \tok.i5_4_lut_adj_186_LC_8_9_6  (
            .in0(N__20162),
            .in1(N__22028),
            .in2(N__17585),
            .in3(N__17582),
            .lcout(\tok.n12_adj_851 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_adj_185_LC_8_9_7 .C_ON=1'b0;
    defparam \tok.i1_3_lut_adj_185_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_adj_185_LC_8_9_7 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i1_3_lut_adj_185_LC_8_9_7  (
            .in0(N__17564),
            .in1(N__20078),
            .in2(_gnd_net_),
            .in3(N__27215),
            .lcout(\tok.n8_adj_850 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A__15__I_16_i5_3_lut_LC_8_10_0 .C_ON=1'b0;
    defparam \tok.A__15__I_16_i5_3_lut_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.A__15__I_16_i5_3_lut_LC_8_10_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.A__15__I_16_i5_3_lut_LC_8_10_0  (
            .in0(N__27392),
            .in1(N__17736),
            .in2(_gnd_net_),
            .in3(N__17411),
            .lcout(\tok.A_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_163_LC_8_10_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_163_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_163_LC_8_10_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.i1_4_lut_adj_163_LC_8_10_1  (
            .in0(N__23018),
            .in1(N__24278),
            .in2(N__17519),
            .in3(N__17606),
            .lcout(\tok.A_15_N_113_4 ),
            .ltout(\tok.A_15_N_113_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i5_LC_8_10_2 .C_ON=1'b0;
    defparam \tok.A_i5_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \tok.A_i5_LC_8_10_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.A_i5_LC_8_10_2  (
            .in0(N__17348),
            .in1(_gnd_net_),
            .in2(N__17405),
            .in3(N__24394),
            .lcout(\tok.A_low_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26265),
            .ce(N__17239),
            .sr(N__19130));
    defparam \tok.i4681_2_lut_LC_8_10_3 .C_ON=1'b0;
    defparam \tok.i4681_2_lut_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4681_2_lut_LC_8_10_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \tok.i4681_2_lut_LC_8_10_3  (
            .in0(N__17737),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17346),
            .lcout(\tok.n950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.A_i1_LC_8_10_4 .C_ON=1'b0;
    defparam \tok.A_i1_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \tok.A_i1_LC_8_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A_i1_LC_8_10_4  (
            .in0(N__17347),
            .in1(N__29572),
            .in2(_gnd_net_),
            .in3(N__17402),
            .lcout(\tok.A_low_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26265),
            .ce(N__17239),
            .sr(N__19130));
    defparam \tok.A_i7_LC_8_10_5 .C_ON=1'b0;
    defparam \tok.A_i7_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \tok.A_i7_LC_8_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.A_i7_LC_8_10_5  (
            .in0(N__21323),
            .in1(N__17349),
            .in2(_gnd_net_),
            .in3(N__17396),
            .lcout(\tok.A_low_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26265),
            .ce(N__17239),
            .sr(N__19130));
    defparam \tok.A_i4_LC_8_10_6 .C_ON=1'b0;
    defparam \tok.A_i4_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \tok.A_i4_LC_8_10_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \tok.A_i4_LC_8_10_6  (
            .in0(N__17693),
            .in1(_gnd_net_),
            .in2(N__17374),
            .in3(N__21546),
            .lcout(\tok.A_low_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26265),
            .ce(N__17239),
            .sr(N__19130));
    defparam \tok.A__15__I_16_i4_3_lut_LC_8_10_7 .C_ON=1'b0;
    defparam \tok.A__15__I_16_i4_3_lut_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.A__15__I_16_i4_3_lut_LC_8_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.A__15__I_16_i4_3_lut_LC_8_10_7  (
            .in0(N__17735),
            .in1(N__17692),
            .in2(_gnd_net_),
            .in3(N__21796),
            .lcout(\tok.A_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4375_4_lut_LC_8_11_0 .C_ON=1'b0;
    defparam \tok.i4375_4_lut_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4375_4_lut_LC_8_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \tok.i4375_4_lut_LC_8_11_0  (
            .in0(N__27228),
            .in1(N__26485),
            .in2(N__26597),
            .in3(N__24268),
            .lcout(),
            .ltout(\tok.n4528_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_LC_8_11_1 .C_ON=1'b0;
    defparam \tok.i6_4_lut_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_LC_8_11_1 .LUT_INIT=16'b1111111101001111;
    LogicCell40 \tok.i6_4_lut_LC_8_11_1  (
            .in0(N__29278),
            .in1(N__27713),
            .in2(N__17678),
            .in3(N__17651),
            .lcout(\tok.n892 ),
            .ltout(\tok.n892_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_174_LC_8_11_2 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_174_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_174_LC_8_11_2 .LUT_INIT=16'b1111111100011101;
    LogicCell40 \tok.i2_4_lut_adj_174_LC_8_11_2  (
            .in0(N__26562),
            .in1(N__21989),
            .in2(N__17675),
            .in3(N__17672),
            .lcout(\tok.n13_adj_842 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_4_lut_adj_165_LC_8_11_3 .C_ON=1'b0;
    defparam \tok.i1_3_lut_4_lut_adj_165_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_4_lut_adj_165_LC_8_11_3 .LUT_INIT=16'b0011101100110011;
    LogicCell40 \tok.i1_3_lut_4_lut_adj_165_LC_8_11_3  (
            .in0(N__29820),
            .in1(N__24456),
            .in2(N__24621),
            .in3(N__27986),
            .lcout(\tok.n8_adj_666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i8_1_lut_2_lut_4_lut_LC_8_11_4 .C_ON=1'b0;
    defparam \tok.i8_1_lut_2_lut_4_lut_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i8_1_lut_2_lut_4_lut_LC_8_11_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \tok.i8_1_lut_2_lut_4_lut_LC_8_11_4  (
            .in0(N__30390),
            .in1(N__29819),
            .in2(N__28013),
            .in3(N__30111),
            .lcout(\tok.n8_adj_777 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i54_3_lut_LC_8_11_5 .C_ON=1'b0;
    defparam \tok.i54_3_lut_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i54_3_lut_LC_8_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.i54_3_lut_LC_8_11_5  (
            .in0(N__27423),
            .in1(N__26563),
            .in2(_gnd_net_),
            .in3(N__17888),
            .lcout(),
            .ltout(\tok.n4502_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4_4_lut_adj_159_LC_8_11_6 .C_ON=1'b0;
    defparam \tok.i4_4_lut_adj_159_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i4_4_lut_adj_159_LC_8_11_6 .LUT_INIT=16'b0010111100111111;
    LogicCell40 \tok.i4_4_lut_adj_159_LC_8_11_6  (
            .in0(N__26919),
            .in1(N__26814),
            .in2(N__17609),
            .in3(N__29036),
            .lcout(\tok.n12_adj_830 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4678_4_lut_4_lut_LC_8_11_7 .C_ON=1'b0;
    defparam \tok.i4678_4_lut_4_lut_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i4678_4_lut_4_lut_LC_8_11_7 .LUT_INIT=16'b0000101000111111;
    LogicCell40 \tok.i4678_4_lut_4_lut_LC_8_11_7  (
            .in0(N__30112),
            .in1(N__27987),
            .in2(N__29864),
            .in3(N__30391),
            .lcout(\tok.n4607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_11_i9_2_lut_LC_8_12_0 .C_ON=1'b0;
    defparam \tok.select_73_Select_11_i9_2_lut_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_11_i9_2_lut_LC_8_12_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tok.select_73_Select_11_i9_2_lut_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__20870),
            .in2(_gnd_net_),
            .in3(N__29421),
            .lcout(\tok.n9_adj_689 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_99_i9_2_lut_LC_8_12_1 .C_ON=1'b0;
    defparam \tok.or_99_i9_2_lut_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i9_2_lut_LC_8_12_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \tok.or_99_i9_2_lut_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__28324),
            .in2(_gnd_net_),
            .in3(N__27399),
            .lcout(),
            .ltout(\tok.n181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_35_LC_8_12_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_35_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_35_LC_8_12_2 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \tok.i1_4_lut_adj_35_LC_8_12_2  (
            .in0(N__24844),
            .in1(N__17893),
            .in2(N__17963),
            .in3(N__26796),
            .lcout(),
            .ltout(\tok.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_LC_8_12_3 .C_ON=1'b0;
    defparam \tok.i9_4_lut_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_LC_8_12_3 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \tok.i9_4_lut_LC_8_12_3  (
            .in0(N__28283),
            .in1(N__21813),
            .in2(N__17960),
            .in3(N__24725),
            .lcout(),
            .ltout(\tok.n20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4670_4_lut_LC_8_12_4 .C_ON=1'b0;
    defparam \tok.i4670_4_lut_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4670_4_lut_LC_8_12_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.i4670_4_lut_LC_8_12_4  (
            .in0(N__17957),
            .in1(N__21560),
            .in2(N__17948),
            .in3(N__17945),
            .lcout(\tok.n4684 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_99_i13_2_lut_LC_8_12_5 .C_ON=1'b0;
    defparam \tok.or_99_i13_2_lut_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i13_2_lut_LC_8_12_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \tok.or_99_i13_2_lut_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__28323),
            .in2(_gnd_net_),
            .in3(N__24843),
            .lcout(),
            .ltout(\tok.n177_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_61_LC_8_12_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_61_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_61_LC_8_12_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \tok.i1_4_lut_adj_61_LC_8_12_6  (
            .in0(N__22994),
            .in1(N__17892),
            .in2(N__17834),
            .in3(N__26795),
            .lcout(),
            .ltout(\tok.n12_adj_696_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i9_4_lut_adj_64_LC_8_12_7 .C_ON=1'b0;
    defparam \tok.i9_4_lut_adj_64_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.i9_4_lut_adj_64_LC_8_12_7 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \tok.i9_4_lut_adj_64_LC_8_12_7  (
            .in0(N__19826),
            .in1(N__27323),
            .in2(N__17831),
            .in3(N__24724),
            .lcout(\tok.n20_adj_700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_2_lut_LC_8_13_0 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_2_lut_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_2_lut_LC_8_13_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_2_lut_LC_8_13_0  (
            .in0(N__17786),
            .in1(N__17785),
            .in2(N__19405),
            .in3(N__17753),
            .lcout(\tok.n33_adj_663 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\tok.n3888 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_3_lut_LC_8_13_1 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_3_lut_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_3_lut_LC_8_13_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_3_lut_LC_8_13_1  (
            .in0(N__18407),
            .in1(N__18406),
            .in2(N__19430),
            .in3(N__18368),
            .lcout(\tok.n33_adj_841 ),
            .ltout(),
            .carryin(\tok.n3888 ),
            .carryout(\tok.n3889 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_4_lut_LC_8_13_2 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_4_lut_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_4_lut_LC_8_13_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_4_lut_LC_8_13_2  (
            .in0(N__18333),
            .in1(N__18332),
            .in2(N__19406),
            .in3(N__18299),
            .lcout(\tok.n33_adj_665 ),
            .ltout(),
            .carryin(\tok.n3889 ),
            .carryout(\tok.n3890 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_5_lut_LC_8_13_3 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_5_lut_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_5_lut_LC_8_13_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_5_lut_LC_8_13_3  (
            .in0(N__18263),
            .in1(N__18262),
            .in2(N__19431),
            .in3(N__18224),
            .lcout(\tok.n33_adj_755 ),
            .ltout(),
            .carryin(\tok.n3890 ),
            .carryout(\tok.n3891 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_6_lut_LC_8_13_4 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_6_lut_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_6_lut_LC_8_13_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_6_lut_LC_8_13_4  (
            .in0(N__18213),
            .in1(N__18212),
            .in2(N__19407),
            .in3(N__18140),
            .lcout(\tok.n33_adj_852 ),
            .ltout(),
            .carryin(\tok.n3891 ),
            .carryout(\tok.n3892 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_7_lut_LC_8_13_5 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_7_lut_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_7_lut_LC_8_13_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_7_lut_LC_8_13_5  (
            .in0(N__18113),
            .in1(N__18112),
            .in2(N__19432),
            .in3(N__18074),
            .lcout(\tok.n33_adj_817 ),
            .ltout(),
            .carryin(\tok.n3892 ),
            .carryout(\tok.n3893 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_8_lut_LC_8_13_6 .C_ON=1'b1;
    defparam \tok.idx_7__I_0_8_lut_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_8_lut_LC_8_13_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_8_lut_LC_8_13_6  (
            .in0(N__19214),
            .in1(N__19215),
            .in2(N__19408),
            .in3(N__18071),
            .lcout(\tok.n33 ),
            .ltout(),
            .carryin(\tok.n3893 ),
            .carryout(\tok.n3894 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_7__I_0_9_lut_LC_8_13_7 .C_ON=1'b0;
    defparam \tok.idx_7__I_0_9_lut_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.idx_7__I_0_9_lut_LC_8_13_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \tok.idx_7__I_0_9_lut_LC_8_13_7  (
            .in0(N__18044),
            .in1(N__18045),
            .in2(N__19433),
            .in3(N__18002),
            .lcout(\tok.n33_adj_643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i12_LC_9_2_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i12_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i12_LC_9_2_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i12_LC_9_2_0  (
            .in0(N__25708),
            .in1(N__17990),
            .in2(_gnd_net_),
            .in3(N__25327),
            .lcout(\tok.tail_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26231),
            .ce(N__25471),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i18_LC_9_2_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i18_LC_9_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i18_LC_9_2_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i18_LC_9_2_1  (
            .in0(N__25751),
            .in1(N__18536),
            .in2(_gnd_net_),
            .in3(N__25714),
            .lcout(\tok.C_stk.tail_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26231),
            .ce(N__25471),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i15_LC_9_2_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i15_LC_9_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i15_LC_9_2_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i15_LC_9_2_2  (
            .in0(N__25709),
            .in1(N__22838),
            .in2(_gnd_net_),
            .in3(N__18562),
            .lcout(\tok.tail_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26231),
            .ce(N__25471),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i0_LC_9_2_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i0_LC_9_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i0_LC_9_2_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.C_stk.tail_i0_i0_LC_9_2_3  (
            .in0(N__22874),
            .in1(N__25712),
            .in2(_gnd_net_),
            .in3(N__18604),
            .lcout(\tok.C_stk.tail_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26231),
            .ce(N__25471),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i7_LC_9_2_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i7_LC_9_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i7_LC_9_2_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \tok.C_stk.tail_i0_i7_LC_9_2_4  (
            .in0(N__25711),
            .in1(_gnd_net_),
            .in2(N__22855),
            .in3(N__18746),
            .lcout(\tok.C_stk.tail_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26231),
            .ce(N__25471),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i4_LC_9_2_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i4_LC_9_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i4_LC_9_2_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.C_stk.tail_i0_i4_LC_9_2_5  (
            .in0(N__18524),
            .in1(N__25713),
            .in2(_gnd_net_),
            .in3(N__30538),
            .lcout(\tok.C_stk.tail_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26231),
            .ce(N__25471),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i44_LC_9_2_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i44_LC_9_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i44_LC_9_2_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i44_LC_9_2_6  (
            .in0(N__25710),
            .in1(N__23231),
            .in2(_gnd_net_),
            .in3(N__18511),
            .lcout(\tok.tail_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26231),
            .ce(N__25471),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i48_LC_9_2_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i48_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i48_LC_9_2_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i48_LC_9_2_7  (
            .in0(N__18500),
            .in1(N__18481),
            .in2(_gnd_net_),
            .in3(N__25715),
            .lcout(\tok.tail_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26231),
            .ce(N__25471),
            .sr(_gnd_net_));
    defparam \tok.i4634_2_lut_3_lut_LC_9_3_0 .C_ON=1'b0;
    defparam \tok.i4634_2_lut_3_lut_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4634_2_lut_3_lut_LC_9_3_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.i4634_2_lut_3_lut_LC_9_3_0  (
            .in0(N__18449),
            .in1(N__29035),
            .in2(_gnd_net_),
            .in3(N__29857),
            .lcout(),
            .ltout(\tok.n4694_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_LC_9_3_1 .C_ON=1'b0;
    defparam \tok.i27_4_lut_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_LC_9_3_1 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \tok.i27_4_lut_LC_9_3_1  (
            .in0(N__18572),
            .in1(N__28549),
            .in2(N__18440),
            .in3(N__30161),
            .lcout(),
            .ltout(\tok.n13_adj_713_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_71_LC_9_3_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_71_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_71_LC_9_3_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_71_LC_9_3_2  (
            .in0(N__18672),
            .in1(N__25251),
            .in2(N__18611),
            .in3(N__25191),
            .lcout(n10_adj_875),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.n602_bdd_4_lut_4739_LC_9_3_3 .C_ON=1'b0;
    defparam \tok.C_stk.n602_bdd_4_lut_4739_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.n602_bdd_4_lut_4739_LC_9_3_3 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \tok.C_stk.n602_bdd_4_lut_4739_LC_9_3_3  (
            .in0(N__25106),
            .in1(N__26347),
            .in2(N__19469),
            .in3(N__18673),
            .lcout(),
            .ltout(\tok.C_stk.n4894_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i0_LC_9_3_4 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i0_LC_9_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i0_LC_9_3_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \tok.C_stk.head_i0_i0_LC_9_3_4  (
            .in0(N__26348),
            .in1(N__22888),
            .in2(N__18608),
            .in3(N__18602),
            .lcout(\tok.c_stk_r_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26237),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i4666_4_lut_LC_9_3_5 .C_ON=1'b0;
    defparam \tok.ram.i4666_4_lut_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i4666_4_lut_LC_9_3_5 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.ram.i4666_4_lut_LC_9_3_5  (
            .in0(N__26695),
            .in1(N__18671),
            .in2(N__18605),
            .in3(N__25996),
            .lcout(),
            .ltout(\tok.ram.n4717_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5_4_lut_LC_9_3_6 .C_ON=1'b0;
    defparam \tok.ram.i5_4_lut_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5_4_lut_LC_9_3_6 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.ram.i5_4_lut_LC_9_3_6  (
            .in0(N__18603),
            .in1(N__25884),
            .in2(N__18575),
            .in3(N__29856),
            .lcout(\tok.n1_adj_712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.n602_bdd_4_lut_LC_9_4_0 .C_ON=1'b0;
    defparam \tok.C_stk.n602_bdd_4_lut_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.n602_bdd_4_lut_LC_9_4_0 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \tok.C_stk.n602_bdd_4_lut_LC_9_4_0  (
            .in0(N__18879),
            .in1(N__25101),
            .in2(N__18845),
            .in3(N__26359),
            .lcout(),
            .ltout(\tok.C_stk.n4912_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i7_LC_9_4_1 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i7_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i7_LC_9_4_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \tok.C_stk.head_i0_i7_LC_9_4_1  (
            .in0(N__26360),
            .in1(N__18566),
            .in2(N__18551),
            .in3(N__18743),
            .lcout(\tok.c_stk_r_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26242),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_137_LC_9_4_2 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_137_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_137_LC_9_4_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.i26_3_lut_adj_137_LC_9_4_2  (
            .in0(N__18803),
            .in1(N__23518),
            .in2(_gnd_net_),
            .in3(N__18814),
            .lcout(\tok.tc_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i4637_4_lut_LC_9_4_3 .C_ON=1'b0;
    defparam \tok.ram.i4637_4_lut_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i4637_4_lut_LC_9_4_3 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \tok.ram.i4637_4_lut_LC_9_4_3  (
            .in0(N__26694),
            .in1(N__25995),
            .in2(N__18745),
            .in3(N__18878),
            .lcout(),
            .ltout(\tok.ram.n4696_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5_4_lut_adj_26_LC_9_4_4 .C_ON=1'b0;
    defparam \tok.ram.i5_4_lut_adj_26_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5_4_lut_adj_26_LC_9_4_4 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.ram.i5_4_lut_adj_26_LC_9_4_4  (
            .in0(N__25873),
            .in1(N__18739),
            .in2(N__18710),
            .in3(N__29873),
            .lcout(),
            .ltout(\tok.n1_adj_798_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_132_LC_9_4_5 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_132_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_132_LC_9_4_5 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i27_4_lut_adj_132_LC_9_4_5  (
            .in0(N__18707),
            .in1(N__28531),
            .in2(N__18701),
            .in3(N__30160),
            .lcout(\tok.n13_adj_799 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_148_LC_9_4_6 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_148_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_148_LC_9_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.i26_3_lut_adj_148_LC_9_4_6  (
            .in0(N__19468),
            .in1(N__19480),
            .in2(_gnd_net_),
            .in3(N__23517),
            .lcout(\tok.tc_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_2_lut_LC_9_5_0 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_2_lut_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_2_lut_LC_9_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_2_lut_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__19454),
            .in2(_gnd_net_),
            .in3(N__18653),
            .lcout(\tok.tc_plus_1_0 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\tok.n3895 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_3_lut_LC_9_5_1 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_3_lut_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_3_lut_LC_9_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_3_lut_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__18764),
            .in2(_gnd_net_),
            .in3(N__18626),
            .lcout(\tok.tc_plus_1_1 ),
            .ltout(),
            .carryin(\tok.n3895 ),
            .carryout(\tok.n3896 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_4_lut_LC_9_5_2 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_4_lut_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_4_lut_LC_9_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_4_lut_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__25034),
            .in2(_gnd_net_),
            .in3(N__18623),
            .lcout(\tok.tc_plus_1_2 ),
            .ltout(),
            .carryin(\tok.n3896 ),
            .carryout(\tok.n3897 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_5_lut_LC_9_5_3 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_5_lut_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_5_lut_LC_9_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_5_lut_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__23555),
            .in2(_gnd_net_),
            .in3(N__18620),
            .lcout(\tok.tc_plus_1_3 ),
            .ltout(),
            .carryin(\tok.n3897 ),
            .carryout(\tok.n3898 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_6_lut_LC_9_5_4 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_6_lut_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_6_lut_LC_9_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_6_lut_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__25352),
            .in2(_gnd_net_),
            .in3(N__18617),
            .lcout(\tok.tc_plus_1_4 ),
            .ltout(),
            .carryin(\tok.n3898 ),
            .carryout(\tok.n3899 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_7_lut_LC_9_5_5 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_7_lut_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_7_lut_LC_9_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_7_lut_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__23684),
            .in2(_gnd_net_),
            .in3(N__18614),
            .lcout(\tok.tc_plus_1_5 ),
            .ltout(),
            .carryin(\tok.n3899 ),
            .carryout(\tok.n3900 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_8_lut_LC_9_5_6 .C_ON=1'b1;
    defparam \tok.tc_7__I_0_8_lut_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_8_lut_LC_9_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_8_lut_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__18794),
            .in2(_gnd_net_),
            .in3(N__18896),
            .lcout(\tok.tc_plus_1_6 ),
            .ltout(),
            .carryin(\tok.n3900 ),
            .carryout(\tok.n3901 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_7__I_0_9_lut_LC_9_5_7 .C_ON=1'b0;
    defparam \tok.tc_7__I_0_9_lut_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.tc_7__I_0_9_lut_LC_9_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.tc_7__I_0_9_lut_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__18836),
            .in2(_gnd_net_),
            .in3(N__18893),
            .lcout(\tok.tc_plus_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.tc_i7_LC_9_6_0 .C_ON=1'b0;
    defparam \tok.tc_i7_LC_9_6_0 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i7_LC_9_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.tc_i7_LC_9_6_0  (
            .in0(N__23502),
            .in1(N__18860),
            .in2(_gnd_net_),
            .in3(N__18841),
            .lcout(c_stk_w_7_N_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26252),
            .ce(),
            .sr(N__19151));
    defparam \tok.tc_i6_LC_9_6_1 .C_ON=1'b0;
    defparam \tok.tc_i6_LC_9_6_1 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i6_LC_9_6_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.tc_i6_LC_9_6_1  (
            .in0(N__18801),
            .in1(N__23505),
            .in2(_gnd_net_),
            .in3(N__18815),
            .lcout(c_stk_w_7_N_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26252),
            .ce(),
            .sr(N__19151));
    defparam \tok.tc_i5_LC_9_6_2 .C_ON=1'b0;
    defparam \tok.tc_i5_LC_9_6_2 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i5_LC_9_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.tc_i5_LC_9_6_2  (
            .in0(N__23501),
            .in1(N__23711),
            .in2(_gnd_net_),
            .in3(N__23691),
            .lcout(c_stk_w_7_N_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26252),
            .ce(),
            .sr(N__19151));
    defparam \tok.tc_i4_LC_9_6_3 .C_ON=1'b0;
    defparam \tok.tc_i4_LC_9_6_3 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i4_LC_9_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.tc_i4_LC_9_6_3  (
            .in0(N__25151),
            .in1(N__25359),
            .in2(_gnd_net_),
            .in3(N__23506),
            .lcout(c_stk_w_7_N_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26252),
            .ce(),
            .sr(N__19151));
    defparam \tok.tc_i3_LC_9_6_4 .C_ON=1'b0;
    defparam \tok.tc_i3_LC_9_6_4 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i3_LC_9_6_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.tc_i3_LC_9_6_4  (
            .in0(N__23500),
            .in1(_gnd_net_),
            .in2(N__23585),
            .in3(N__23562),
            .lcout(c_stk_w_7_N_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26252),
            .ce(),
            .sr(N__19151));
    defparam \tok.tc_i2_LC_9_6_5 .C_ON=1'b0;
    defparam \tok.tc_i2_LC_9_6_5 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i2_LC_9_6_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.tc_i2_LC_9_6_5  (
            .in0(N__23654),
            .in1(N__23504),
            .in2(_gnd_net_),
            .in3(N__25041),
            .lcout(c_stk_w_7_N_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26252),
            .ce(),
            .sr(N__19151));
    defparam \tok.tc_i1_LC_9_6_6 .C_ON=1'b0;
    defparam \tok.tc_i1_LC_9_6_6 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i1_LC_9_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.tc_i1_LC_9_6_6  (
            .in0(N__23499),
            .in1(N__18773),
            .in2(_gnd_net_),
            .in3(N__18767),
            .lcout(c_stk_w_7_N_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26252),
            .ce(),
            .sr(N__19151));
    defparam \tok.tc_i0_LC_9_6_7 .C_ON=1'b0;
    defparam \tok.tc_i0_LC_9_6_7 .SEQ_MODE=4'b1011;
    defparam \tok.tc_i0_LC_9_6_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \tok.tc_i0_LC_9_6_7  (
            .in0(N__19484),
            .in1(N__23503),
            .in2(_gnd_net_),
            .in3(N__19461),
            .lcout(c_stk_w_7_N_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26252),
            .ce(),
            .sr(N__19151));
    defparam \tok.i1_2_lut_adj_37_LC_9_7_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_37_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_37_LC_9_7_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \tok.i1_2_lut_adj_37_LC_9_7_0  (
            .in0(N__22261),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19377),
            .lcout(\tok.n5_adj_655 ),
            .ltout(\tok.n5_adj_655_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_38_LC_9_7_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_38_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_38_LC_9_7_1 .LUT_INIT=16'b1011101010111011;
    LogicCell40 \tok.i1_4_lut_adj_38_LC_9_7_1  (
            .in0(N__19005),
            .in1(N__18989),
            .in2(N__19349),
            .in3(N__22450),
            .lcout(stall_),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_105_LC_9_7_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_105_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_105_LC_9_7_2 .LUT_INIT=16'b0010001000101111;
    LogicCell40 \tok.i1_4_lut_adj_105_LC_9_7_2  (
            .in0(N__19346),
            .in1(N__24066),
            .in2(N__19312),
            .in3(N__27050),
            .lcout(\tok.uart_stall ),
            .ltout(\tok.uart_stall_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2655_2_lut_LC_9_7_3 .C_ON=1'b0;
    defparam \tok.i2655_2_lut_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2655_2_lut_LC_9_7_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \tok.i2655_2_lut_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19283),
            .in3(N__18990),
            .lcout(\tok.n2732 ),
            .ltout(\tok.n2732_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.idx_i6_LC_9_7_4 .C_ON=1'b0;
    defparam \tok.idx_i6_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \tok.idx_i6_LC_9_7_4 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \tok.idx_i6_LC_9_7_4  (
            .in0(N__19184),
            .in1(N__18940),
            .in2(N__19232),
            .in3(N__22748),
            .lcout(\tok.n43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26257),
            .ce(),
            .sr(N__19143));
    defparam \tok.stall_200_LC_9_7_6 .C_ON=1'b0;
    defparam \tok.stall_200_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \tok.stall_200_LC_9_7_6 .LUT_INIT=16'b1111111100001101;
    LogicCell40 \tok.stall_200_LC_9_7_6  (
            .in0(N__22451),
            .in1(N__19157),
            .in2(N__18995),
            .in3(N__19007),
            .lcout(\tok.stall ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26257),
            .ce(),
            .sr(N__19143));
    defparam \tok.i1_4_lut_adj_179_LC_9_7_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_179_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_179_LC_9_7_7 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \tok.i1_4_lut_adj_179_LC_9_7_7  (
            .in0(N__19006),
            .in1(N__22262),
            .in2(N__22489),
            .in3(N__18991),
            .lcout(\tok.n4431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_2_lut_LC_9_8_0 .C_ON=1'b1;
    defparam \tok.add_104_2_lut_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_2_lut_LC_9_8_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \tok.add_104_2_lut_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__26900),
            .in2(N__29574),
            .in3(N__27661),
            .lcout(\tok.n5_adj_682 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\tok.n3925 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_3_lut_LC_9_8_1 .C_ON=1'b1;
    defparam \tok.add_104_3_lut_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_3_lut_LC_9_8_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_3_lut_LC_9_8_1  (
            .in0(N__27660),
            .in1(N__24173),
            .in2(N__20169),
            .in3(N__20072),
            .lcout(\tok.n4_adj_790 ),
            .ltout(),
            .carryin(\tok.n3925 ),
            .carryout(\tok.n3926 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_4_lut_LC_9_8_2 .C_ON=1'b1;
    defparam \tok.add_104_4_lut_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_4_lut_LC_9_8_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_4_lut_LC_9_8_2  (
            .in0(N__27667),
            .in1(N__21981),
            .in2(N__20060),
            .in3(N__19961),
            .lcout(\tok.n5_adj_789 ),
            .ltout(),
            .carryin(\tok.n3926 ),
            .carryout(\tok.n3927 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_5_lut_LC_9_8_3 .C_ON=1'b1;
    defparam \tok.add_104_5_lut_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_5_lut_LC_9_8_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_5_lut_LC_9_8_3  (
            .in0(N__27657),
            .in1(N__21824),
            .in2(N__21544),
            .in3(N__19958),
            .lcout(\tok.n23_adj_788 ),
            .ltout(),
            .carryin(\tok.n3927 ),
            .carryout(\tok.n3928 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_6_lut_LC_9_8_4 .C_ON=1'b1;
    defparam \tok.add_104_6_lut_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_6_lut_LC_9_8_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_6_lut_LC_9_8_4  (
            .in0(N__27666),
            .in1(N__27411),
            .in2(N__24389),
            .in3(N__19955),
            .lcout(\tok.n13_adj_787 ),
            .ltout(),
            .carryin(\tok.n3928 ),
            .carryout(\tok.n3929 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_7_lut_LC_9_8_5 .C_ON=1'b1;
    defparam \tok.add_104_7_lut_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_7_lut_LC_9_8_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_7_lut_LC_9_8_5  (
            .in0(N__27659),
            .in1(N__22389),
            .in2(N__19951),
            .in3(N__19844),
            .lcout(\tok.n5_adj_775 ),
            .ltout(),
            .carryin(\tok.n3929 ),
            .carryout(\tok.n3930 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_8_lut_LC_9_8_6 .C_ON=1'b1;
    defparam \tok.add_104_8_lut_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_8_lut_LC_9_8_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_8_lut_LC_9_8_6  (
            .in0(N__27668),
            .in1(N__28232),
            .in2(N__21321),
            .in3(N__19829),
            .lcout(\tok.n5_adj_773 ),
            .ltout(),
            .carryin(\tok.n3930 ),
            .carryout(\tok.n3931 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_9_lut_LC_9_8_7 .C_ON=1'b1;
    defparam \tok.add_104_9_lut_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_9_lut_LC_9_8_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_9_lut_LC_9_8_7  (
            .in0(N__27658),
            .in1(N__19775),
            .in2(N__19678),
            .in3(N__19574),
            .lcout(\tok.n5_adj_752 ),
            .ltout(),
            .carryin(\tok.n3931 ),
            .carryout(\tok.n3932 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_10_lut_LC_9_9_0 .C_ON=1'b1;
    defparam \tok.add_104_10_lut_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_10_lut_LC_9_9_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_10_lut_LC_9_9_0  (
            .in0(N__27653),
            .in1(N__19562),
            .in2(N__24856),
            .in3(N__19487),
            .lcout(\tok.n5 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\tok.n3933 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_11_lut_LC_9_9_1 .C_ON=1'b1;
    defparam \tok.add_104_11_lut_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_11_lut_LC_9_9_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_11_lut_LC_9_9_1  (
            .in0(N__27664),
            .in1(N__22656),
            .in2(N__21182),
            .in3(N__21071),
            .lcout(\tok.n21 ),
            .ltout(),
            .carryin(\tok.n3933 ),
            .carryout(\tok.n3934 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_12_lut_LC_9_9_2 .C_ON=1'b1;
    defparam \tok.add_104_12_lut_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_12_lut_LC_9_9_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_12_lut_LC_9_9_2  (
            .in0(N__27656),
            .in1(N__21055),
            .in2(N__20965),
            .in3(N__20873),
            .lcout(\tok.n5_adj_668 ),
            .ltout(),
            .carryin(\tok.n3934 ),
            .carryout(\tok.n3935 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_13_lut_LC_9_9_3 .C_ON=1'b1;
    defparam \tok.add_104_13_lut_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_13_lut_LC_9_9_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_13_lut_LC_9_9_3  (
            .in0(N__27663),
            .in1(N__21434),
            .in2(N__20869),
            .in3(N__20765),
            .lcout(\tok.n5_adj_690 ),
            .ltout(),
            .carryin(\tok.n3935 ),
            .carryout(\tok.n3936 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_14_lut_LC_9_9_4 .C_ON=1'b1;
    defparam \tok.add_104_14_lut_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_14_lut_LC_9_9_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_14_lut_LC_9_9_4  (
            .in0(N__27654),
            .in1(N__23005),
            .in2(N__20760),
            .in3(N__20684),
            .lcout(\tok.n5_adj_694 ),
            .ltout(),
            .carryin(\tok.n3936 ),
            .carryout(\tok.n3937 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_15_lut_LC_9_9_5 .C_ON=1'b1;
    defparam \tok.add_104_15_lut_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_15_lut_LC_9_9_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_15_lut_LC_9_9_5  (
            .in0(N__27665),
            .in1(N__20676),
            .in2(N__20595),
            .in3(N__20513),
            .lcout(\tok.n5_adj_710 ),
            .ltout(),
            .carryin(\tok.n3937 ),
            .carryout(\tok.n3938 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_16_lut_LC_9_9_6 .C_ON=1'b1;
    defparam \tok.add_104_16_lut_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_16_lut_LC_9_9_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_16_lut_LC_9_9_6  (
            .in0(N__27655),
            .in1(N__20510),
            .in2(N__24014),
            .in3(N__20405),
            .lcout(\tok.n5_adj_729 ),
            .ltout(),
            .carryin(\tok.n3938 ),
            .carryout(\tok.n3939 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.add_104_17_lut_LC_9_9_7 .C_ON=1'b0;
    defparam \tok.add_104_17_lut_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.add_104_17_lut_LC_9_9_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.add_104_17_lut_LC_9_9_7  (
            .in0(N__27662),
            .in1(N__20399),
            .in2(N__20321),
            .in3(N__20216),
            .lcout(\tok.n5_adj_750 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_167_LC_9_10_0 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_167_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_167_LC_9_10_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_167_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__20198),
            .in2(_gnd_net_),
            .in3(N__20183),
            .lcout(),
            .ltout(\tok.n5_adj_837_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_168_LC_9_10_1 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_168_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_168_LC_9_10_1 .LUT_INIT=16'b1111111101010100;
    LogicCell40 \tok.i3_4_lut_adj_168_LC_9_10_1  (
            .in0(N__29293),
            .in1(N__21347),
            .in2(N__21554),
            .in3(N__22004),
            .lcout(),
            .ltout(\tok.n10_adj_838_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_170_LC_9_10_2 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_170_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_170_LC_9_10_2 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i5_4_lut_adj_170_LC_9_10_2  (
            .in0(N__21545),
            .in1(N__21461),
            .in2(N__21452),
            .in3(N__29392),
            .lcout(\tok.n12_adj_840 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_166_LC_9_10_3 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_166_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_166_LC_9_10_3 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \tok.i2_4_lut_adj_166_LC_9_10_3  (
            .in0(N__27781),
            .in1(N__21435),
            .in2(N__21194),
            .in3(N__27571),
            .lcout(\tok.n6_adj_835 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_99_LC_9_10_4 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_99_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_99_LC_9_10_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i1_2_lut_adj_99_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__29292),
            .in2(_gnd_net_),
            .in3(N__27780),
            .lcout(\tok.n109 ),
            .ltout(\tok.n109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_120_LC_9_10_5 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_120_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_120_LC_9_10_5 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \tok.i6_4_lut_adj_120_LC_9_10_5  (
            .in0(N__29393),
            .in1(N__21341),
            .in2(N__21326),
            .in3(N__21319),
            .lcout(\tok.n18_adj_782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_102_LC_9_10_6 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_102_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_102_LC_9_10_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i1_2_lut_adj_102_LC_9_10_6  (
            .in0(N__27570),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29294),
            .lcout(\tok.n101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i3_LC_9_10_7 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i3_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i3_LC_9_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.rx_data_i0_i3_LC_9_10_7  (
            .in0(N__21193),
            .in1(N__21221),
            .in2(_gnd_net_),
            .in3(N__22123),
            .lcout(uart_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26268),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_2_lut_LC_9_11_0 .C_ON=1'b1;
    defparam \tok.i1_2_lut_2_lut_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_2_lut_LC_9_11_0 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \tok.i1_2_lut_2_lut_LC_9_11_0  (
            .in0(N__30322),
            .in1(N__30020),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n40 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\tok.n3902 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_3_lut_LC_9_11_1 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_3_lut_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_3_lut_LC_9_11_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_100_add_2_3_lut_LC_9_11_1  (
            .in0(N__22176),
            .in1(N__30323),
            .in2(_gnd_net_),
            .in3(N__22019),
            .lcout(\tok.n13_adj_816 ),
            .ltout(),
            .carryin(\tok.n3902 ),
            .carryout(\tok.n3903 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_4_lut_LC_9_11_2 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_4_lut_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_4_lut_LC_9_11_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_100_add_2_4_lut_LC_9_11_2  (
            .in0(N__22177),
            .in1(N__29824),
            .in2(_gnd_net_),
            .in3(N__22007),
            .lcout(\tok.n2_adj_811 ),
            .ltout(),
            .carryin(\tok.n3903 ),
            .carryout(\tok.n3904 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_5_lut_LC_9_11_3 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_5_lut_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_5_lut_LC_9_11_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \tok.sub_100_add_2_5_lut_LC_9_11_3  (
            .in0(N__22175),
            .in1(N__27988),
            .in2(N__21689),
            .in3(N__21998),
            .lcout(\tok.n26_adj_808 ),
            .ltout(),
            .carryin(\tok.n3904 ),
            .carryout(\tok.n3905 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_6_lut_LC_9_11_4 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_6_lut_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_6_lut_LC_9_11_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_100_add_2_6_lut_LC_9_11_4  (
            .in0(N__26882),
            .in1(N__28973),
            .in2(_gnd_net_),
            .in3(N__21995),
            .lcout(\tok.n36 ),
            .ltout(),
            .carryin(\tok.n3905 ),
            .carryout(\tok.n3906 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_7_lut_LC_9_11_5 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_7_lut_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_7_lut_LC_9_11_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_100_add_2_7_lut_LC_9_11_5  (
            .in0(N__24180),
            .in1(N__28658),
            .in2(_gnd_net_),
            .in3(N__21992),
            .lcout(\tok.n211 ),
            .ltout(),
            .carryin(\tok.n3906 ),
            .carryout(\tok.n3907 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_8_lut_LC_9_11_6 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_8_lut_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_8_lut_LC_9_11_6 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_100_add_2_8_lut_LC_9_11_6  (
            .in0(N__21986),
            .in1(N__28505),
            .in2(N__21691),
            .in3(N__21854),
            .lcout(\tok.n210 ),
            .ltout(),
            .carryin(\tok.n3907 ),
            .carryout(\tok.n3908 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_9_lut_LC_9_11_7 .C_ON=1'b1;
    defparam \tok.sub_100_add_2_9_lut_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_9_lut_LC_9_11_7 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \tok.sub_100_add_2_9_lut_LC_9_11_7  (
            .in0(N__21794),
            .in1(N__28808),
            .in2(N__21690),
            .in3(N__21704),
            .lcout(\tok.n209 ),
            .ltout(),
            .carryin(\tok.n3908 ),
            .carryout(\tok.n3909 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.sub_100_add_2_10_lut_LC_9_12_0 .C_ON=1'b0;
    defparam \tok.sub_100_add_2_10_lut_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \tok.sub_100_add_2_10_lut_LC_9_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \tok.sub_100_add_2_10_lut_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__21665),
            .in2(_gnd_net_),
            .in3(N__21563),
            .lcout(\tok.n191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2546_2_lut_LC_9_12_1 .C_ON=1'b0;
    defparam \tok.i2546_2_lut_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \tok.i2546_2_lut_LC_9_12_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i2546_2_lut_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__24845),
            .in2(_gnd_net_),
            .in3(N__26599),
            .lcout(\tok.n2598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_5_i2_2_lut_LC_9_12_2 .C_ON=1'b0;
    defparam \tok.select_73_Select_5_i2_2_lut_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_5_i2_2_lut_LC_9_12_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \tok.select_73_Select_5_i2_2_lut_LC_9_12_2  (
            .in0(N__22811),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24471),
            .lcout(\tok.n2_adj_810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4623_3_lut_LC_9_12_3 .C_ON=1'b0;
    defparam \tok.i4623_3_lut_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4623_3_lut_LC_9_12_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \tok.i4623_3_lut_LC_9_12_3  (
            .in0(N__22796),
            .in1(N__22787),
            .in2(_gnd_net_),
            .in3(N__22775),
            .lcout(\tok.n4663 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_LC_9_12_4 .C_ON=1'b0;
    defparam \tok.i50_4_lut_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_LC_9_12_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \tok.i50_4_lut_LC_9_12_4  (
            .in0(N__22490),
            .in1(N__28252),
            .in2(N__22283),
            .in3(N__22754),
            .lcout(\tok.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.inv_106_i7_1_lut_LC_9_12_6 .C_ON=1'b0;
    defparam \tok.inv_106_i7_1_lut_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \tok.inv_106_i7_1_lut_LC_9_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.inv_106_i7_1_lut_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28251),
            .lcout(\tok.n296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_13_i2_3_lut_LC_9_12_7 .C_ON=1'b0;
    defparam \tok.select_73_Select_13_i2_3_lut_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_13_i2_3_lut_LC_9_12_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \tok.select_73_Select_13_i2_3_lut_LC_9_12_7  (
            .in0(N__24472),
            .in1(N__22697),
            .in2(_gnd_net_),
            .in3(N__22657),
            .lcout(\tok.n2_adj_703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i50_4_lut_adj_218_LC_9_13_1 .C_ON=1'b0;
    defparam \tok.i50_4_lut_adj_218_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \tok.i50_4_lut_adj_218_LC_9_13_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \tok.i50_4_lut_adj_218_LC_9_13_1  (
            .in0(N__22491),
            .in1(N__22393),
            .in2(N__22281),
            .in3(N__22196),
            .lcout(\tok.n27_adj_868 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i25_1_lut_LC_9_13_2 .C_ON=1'b0;
    defparam \tok.i25_1_lut_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \tok.i25_1_lut_LC_9_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \tok.i25_1_lut_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24469),
            .lcout(\tok.n82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.uart.rx_data_i0_i4_LC_9_13_3 .C_ON=1'b0;
    defparam \tok.uart.rx_data_i0_i4_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \tok.uart.rx_data_i0_i4_LC_9_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.uart.rx_data_i0_i4_LC_9_13_3  (
            .in0(N__23057),
            .in1(N__22148),
            .in2(_gnd_net_),
            .in3(N__22124),
            .lcout(uart_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26270),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_3_lut_adj_156_LC_9_13_4 .C_ON=1'b0;
    defparam \tok.i2_3_lut_adj_156_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_3_lut_adj_156_LC_9_13_4 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \tok.i2_3_lut_adj_156_LC_9_13_4  (
            .in0(N__23069),
            .in1(N__23003),
            .in2(_gnd_net_),
            .in3(N__27575),
            .lcout(),
            .ltout(\tok.n6_adj_827_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_157_LC_9_13_5 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_157_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_157_LC_9_13_5 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i3_4_lut_adj_157_LC_9_13_5  (
            .in0(N__23056),
            .in1(N__23048),
            .in2(N__23033),
            .in3(N__27795),
            .lcout(),
            .ltout(\tok.n33_adj_828_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_160_LC_9_13_6 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_160_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_160_LC_9_13_6 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \tok.i3_4_lut_adj_160_LC_9_13_6  (
            .in0(N__23030),
            .in1(N__29285),
            .in2(N__23021),
            .in3(N__24470),
            .lcout(\tok.n11_adj_831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2462_2_lut_LC_9_13_7 .C_ON=1'b0;
    defparam \tok.i2462_2_lut_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2462_2_lut_LC_9_13_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \tok.i2462_2_lut_LC_9_13_7  (
            .in0(N__23004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26600),
            .lcout(\tok.n2514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i8_LC_11_2_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i8_LC_11_2_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i8_LC_11_2_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i8_LC_11_2_0  (
            .in0(N__25727),
            .in1(N__23180),
            .in2(_gnd_net_),
            .in3(N__22892),
            .lcout(\tok.tail_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26238),
            .ce(N__25465),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i16_LC_11_2_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i16_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i16_LC_11_2_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i16_LC_11_2_1  (
            .in0(N__22867),
            .in1(N__23155),
            .in2(_gnd_net_),
            .in3(N__25728),
            .lcout(\tok.C_stk.tail_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26238),
            .ce(N__25465),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i23_LC_11_2_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i23_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i23_LC_11_2_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i23_LC_11_2_2  (
            .in0(N__25724),
            .in1(N__22820),
            .in2(_gnd_net_),
            .in3(N__22856),
            .lcout(\tok.C_stk.tail_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26238),
            .ce(N__25465),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i31_LC_11_2_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i31_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i31_LC_11_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i31_LC_11_2_3  (
            .in0(N__22831),
            .in1(N__23198),
            .in2(_gnd_net_),
            .in3(N__25730),
            .lcout(\tok.tail_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26238),
            .ce(N__25465),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i39_LC_11_2_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i39_LC_11_2_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i39_LC_11_2_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i39_LC_11_2_4  (
            .in0(N__25725),
            .in1(N__23189),
            .in2(_gnd_net_),
            .in3(N__22819),
            .lcout(\tok.C_stk.tail_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26238),
            .ce(N__25465),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i47_LC_11_2_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i47_LC_11_2_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i47_LC_11_2_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i47_LC_11_2_5  (
            .in0(N__23290),
            .in1(N__23197),
            .in2(_gnd_net_),
            .in3(N__25731),
            .lcout(\tok.tail_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26238),
            .ce(N__25465),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i55_LC_11_2_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i55_LC_11_2_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i55_LC_11_2_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i55_LC_11_2_6  (
            .in0(N__25726),
            .in1(N__23270),
            .in2(_gnd_net_),
            .in3(N__23188),
            .lcout(\tok.tail_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26238),
            .ce(N__25465),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i24_LC_11_2_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i24_LC_11_2_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i24_LC_11_2_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i24_LC_11_2_7  (
            .in0(N__23179),
            .in1(N__23171),
            .in2(_gnd_net_),
            .in3(N__25729),
            .lcout(\tok.tail_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26238),
            .ce(N__25465),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i30_LC_11_3_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i30_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i30_LC_11_3_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i30_LC_11_3_0  (
            .in0(N__24974),
            .in1(N__23129),
            .in2(_gnd_net_),
            .in3(N__25620),
            .lcout(\tok.tail_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26243),
            .ce(N__25466),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i38_LC_11_3_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i38_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i38_LC_11_3_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \tok.C_stk.tail_i0_i38_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__23137),
            .in2(N__25706),
            .in3(N__23119),
            .lcout(\tok.C_stk.tail_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26243),
            .ce(N__25466),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i22_LC_11_3_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i22_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i22_LC_11_3_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \tok.C_stk.tail_i0_i22_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__25619),
            .in2(N__23141),
            .in3(N__24940),
            .lcout(\tok.C_stk.tail_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26243),
            .ce(N__25466),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i46_LC_11_3_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i46_LC_11_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i46_LC_11_3_3 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \tok.C_stk.tail_i0_i46_LC_11_3_3  (
            .in0(N__23128),
            .in1(N__23254),
            .in2(N__25707),
            .in3(_gnd_net_),
            .lcout(\tok.tail_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26243),
            .ce(N__25466),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i54_LC_11_3_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i54_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i54_LC_11_3_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i54_LC_11_3_4  (
            .in0(N__23120),
            .in1(N__23242),
            .in2(_gnd_net_),
            .in3(N__25622),
            .lcout(\tok.tail_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26243),
            .ce(N__25466),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i6_LC_11_3_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i6_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i6_LC_11_3_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \tok.C_stk.tail_i0_i6_LC_11_3_5  (
            .in0(N__24941),
            .in1(_gnd_net_),
            .in2(N__25704),
            .in3(N__23111),
            .lcout(\tok.C_stk.tail_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26243),
            .ce(N__25466),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i52_LC_11_3_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i52_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i52_LC_11_3_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i52_LC_11_3_6  (
            .in0(N__23210),
            .in1(N__23348),
            .in2(_gnd_net_),
            .in3(N__25621),
            .lcout(\tok.tail_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26243),
            .ce(N__25466),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i10_LC_11_3_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i10_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i10_LC_11_3_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \tok.C_stk.tail_i0_i10_LC_11_3_7  (
            .in0(N__23330),
            .in1(N__26374),
            .in2(N__25705),
            .in3(_gnd_net_),
            .lcout(\tok.tail_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26243),
            .ce(N__25466),
            .sr(_gnd_net_));
    defparam \tok.i547_3_lut_4_lut_LC_11_4_0 .C_ON=1'b0;
    defparam \tok.i547_3_lut_4_lut_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \tok.i547_3_lut_4_lut_LC_11_4_0 .LUT_INIT=16'b1000101010101010;
    LogicCell40 \tok.i547_3_lut_4_lut_LC_11_4_0  (
            .in0(N__25459),
            .in1(N__24623),
            .in2(N__23312),
            .in3(N__28074),
            .lcout(\tok.n602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.i545_2_lut_LC_11_4_1 .C_ON=1'b0;
    defparam \tok.C_stk.i545_2_lut_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.i545_2_lut_LC_11_4_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.C_stk.i545_2_lut_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__23311),
            .in2(_gnd_net_),
            .in3(N__25458),
            .lcout(\tok.C_stk.n600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i63_LC_11_4_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i63_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i63_LC_11_4_3 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i63_LC_11_4_3  (
            .in0(N__23266),
            .in1(N__25697),
            .in2(N__23291),
            .in3(N__25464),
            .lcout(\tok.tail_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26248),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i62_LC_11_4_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i62_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i62_LC_11_4_4 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \tok.C_stk.tail_i0_i62_LC_11_4_4  (
            .in0(N__25461),
            .in1(N__23255),
            .in2(N__25733),
            .in3(N__23243),
            .lcout(\tok.tail_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26248),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i61_LC_11_4_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i61_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i61_LC_11_4_5 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i61_LC_11_4_5  (
            .in0(N__25015),
            .in1(N__25696),
            .in2(N__24995),
            .in3(N__25463),
            .lcout(\tok.tail_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26248),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i60_LC_11_4_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i60_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i60_LC_11_4_6 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \tok.C_stk.tail_i0_i60_LC_11_4_6  (
            .in0(N__25460),
            .in1(N__23230),
            .in2(N__25732),
            .in3(N__23209),
            .lcout(\tok.tail_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26248),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i59_LC_11_4_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i59_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i59_LC_11_4_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i59_LC_11_4_7  (
            .in0(N__24895),
            .in1(N__25695),
            .in2(N__24875),
            .in3(N__25462),
            .lcout(\tok.tail_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26248),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.n602_bdd_4_lut_4744_LC_11_5_0 .C_ON=1'b0;
    defparam \tok.C_stk.n602_bdd_4_lut_4744_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.n602_bdd_4_lut_4744_LC_11_5_0 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \tok.C_stk.n602_bdd_4_lut_4744_LC_11_5_0  (
            .in0(N__25074),
            .in1(N__26304),
            .in2(N__23699),
            .in3(N__23373),
            .lcout(),
            .ltout(\tok.C_stk.n4900_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i5_LC_11_5_1 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i5_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i5_LC_11_5_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \tok.C_stk.head_i0_i5_LC_11_5_1  (
            .in0(N__26305),
            .in1(N__24560),
            .in2(N__23438),
            .in3(N__24584),
            .lcout(\tok.c_stk_r_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26253),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_98_LC_11_5_2 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_98_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_98_LC_11_5_2 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_98_LC_11_5_2  (
            .in0(N__24583),
            .in1(N__30380),
            .in2(N__23435),
            .in3(N__30151),
            .lcout(),
            .ltout(\tok.n83_adj_742_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4619_2_lut_3_lut_LC_11_5_3 .C_ON=1'b0;
    defparam \tok.i4619_2_lut_3_lut_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4619_2_lut_3_lut_LC_11_5_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i4619_2_lut_3_lut_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__28962),
            .in2(N__23402),
            .in3(N__29800),
            .lcout(),
            .ltout(\tok.n4651_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_100_LC_11_5_4 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_100_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_100_LC_11_5_4 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \tok.i27_4_lut_adj_100_LC_11_5_4  (
            .in0(N__23393),
            .in1(N__28504),
            .in2(N__23399),
            .in3(N__30152),
            .lcout(\tok.n13_adj_758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.n602_bdd_4_lut_4729_LC_11_5_5 .C_ON=1'b0;
    defparam \tok.C_stk.n602_bdd_4_lut_4729_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.n602_bdd_4_lut_4729_LC_11_5_5 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \tok.C_stk.n602_bdd_4_lut_4729_LC_11_5_5  (
            .in0(N__26303),
            .in1(N__25073),
            .in2(N__23570),
            .in3(N__23615),
            .lcout(\tok.C_stk.n4882 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i4645_4_lut_LC_11_5_6 .C_ON=1'b0;
    defparam \tok.ram.i4645_4_lut_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i4645_4_lut_LC_11_5_6 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \tok.ram.i4645_4_lut_LC_11_5_6  (
            .in0(N__26683),
            .in1(N__25994),
            .in2(N__24589),
            .in3(N__23372),
            .lcout(),
            .ltout(\tok.ram.n4702_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5_4_lut_adj_24_LC_11_5_7 .C_ON=1'b0;
    defparam \tok.ram.i5_4_lut_adj_24_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5_4_lut_adj_24_LC_11_5_7 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \tok.ram.i5_4_lut_adj_24_LC_11_5_7  (
            .in0(N__24585),
            .in1(N__25899),
            .in2(N__23396),
            .in3(N__29799),
            .lcout(\tok.n1_adj_757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i4654_4_lut_LC_11_6_0 .C_ON=1'b0;
    defparam \tok.ram.i4654_4_lut_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i4654_4_lut_LC_11_6_0 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.ram.i4654_4_lut_LC_11_6_0  (
            .in0(N__26650),
            .in1(N__23619),
            .in2(N__30489),
            .in3(N__25978),
            .lcout(\tok.ram.n4708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_101_LC_11_6_1 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_101_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_101_LC_11_6_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_101_LC_11_6_1  (
            .in0(N__25265),
            .in1(N__25204),
            .in2(N__23387),
            .in3(N__23717),
            .lcout(n10_adj_873),
            .ltout(n10_adj_873_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_138_LC_11_6_2 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_138_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_138_LC_11_6_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.i26_3_lut_adj_138_LC_11_6_2  (
            .in0(N__23521),
            .in1(_gnd_net_),
            .in2(N__23702),
            .in3(N__23692),
            .lcout(\tok.tc_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_81_LC_11_6_3 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_81_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_81_LC_11_6_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \tok.i1_4_lut_adj_81_LC_11_6_3  (
            .in0(N__25916),
            .in1(N__25203),
            .in2(N__25275),
            .in3(N__26032),
            .lcout(n10_adj_874),
            .ltout(n10_adj_874_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_143_LC_11_6_4 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_143_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_143_LC_11_6_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.i26_3_lut_adj_143_LC_11_6_4  (
            .in0(N__23520),
            .in1(_gnd_net_),
            .in2(N__23642),
            .in3(N__25043),
            .lcout(\tok.tc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_88_LC_11_6_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_88_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_88_LC_11_6_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \tok.i1_4_lut_adj_88_LC_11_6_5  (
            .in0(N__23620),
            .in1(N__25205),
            .in2(N__25276),
            .in3(N__25832),
            .lcout(n92_adj_870),
            .ltout(n92_adj_870_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_141_LC_11_6_6 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_141_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_141_LC_11_6_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \tok.i26_3_lut_adj_141_LC_11_6_6  (
            .in0(N__23519),
            .in1(_gnd_net_),
            .in2(N__23573),
            .in3(N__23563),
            .lcout(\tok.tc_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i26_3_lut_adj_139_LC_11_6_7 .C_ON=1'b0;
    defparam \tok.i26_3_lut_adj_139_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \tok.i26_3_lut_adj_139_LC_11_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.i26_3_lut_adj_139_LC_11_6_7  (
            .in0(N__25144),
            .in1(N__25363),
            .in2(_gnd_net_),
            .in3(N__23522),
            .lcout(\tok.tc_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_113_i9_2_lut_LC_11_7_0 .C_ON=1'b0;
    defparam \tok.equal_113_i9_2_lut_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.equal_113_i9_2_lut_LC_11_7_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \tok.equal_113_i9_2_lut_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__30286),
            .in2(_gnd_net_),
            .in3(N__29968),
            .lcout(\tok.n9_adj_645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_220_i11_2_lut_4_lut_LC_11_7_1 .C_ON=1'b0;
    defparam \tok.T_7__I_0_220_i11_2_lut_4_lut_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_220_i11_2_lut_4_lut_LC_11_7_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \tok.T_7__I_0_220_i11_2_lut_4_lut_LC_11_7_1  (
            .in0(N__30288),
            .in1(N__29683),
            .in2(N__30040),
            .in3(N__27884),
            .lcout(\tok.n11_adj_648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_142_i14_2_lut_3_lut_4_lut_LC_11_7_2 .C_ON=1'b0;
    defparam \tok.equal_142_i14_2_lut_3_lut_4_lut_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.equal_142_i14_2_lut_3_lut_4_lut_LC_11_7_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \tok.equal_142_i14_2_lut_3_lut_4_lut_LC_11_7_2  (
            .in0(N__28400),
            .in1(N__28590),
            .in2(N__28773),
            .in3(N__28904),
            .lcout(\tok.n14_adj_650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_119_i10_2_lut_LC_11_7_3 .C_ON=1'b0;
    defparam \tok.equal_119_i10_2_lut_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.equal_119_i10_2_lut_LC_11_7_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \tok.equal_119_i10_2_lut_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__29681),
            .in2(_gnd_net_),
            .in3(N__27880),
            .lcout(\tok.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_120_i14_2_lut_3_lut_4_lut_LC_11_7_4 .C_ON=1'b0;
    defparam \tok.equal_120_i14_2_lut_3_lut_4_lut_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.equal_120_i14_2_lut_3_lut_4_lut_LC_11_7_4 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \tok.equal_120_i14_2_lut_3_lut_4_lut_LC_11_7_4  (
            .in0(N__28402),
            .in1(N__28594),
            .in2(N__28774),
            .in3(N__28905),
            .lcout(\tok.n14_adj_702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_121_i9_2_lut_LC_11_7_5 .C_ON=1'b0;
    defparam \tok.equal_121_i9_2_lut_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.equal_121_i9_2_lut_LC_11_7_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \tok.equal_121_i9_2_lut_LC_11_7_5  (
            .in0(N__30287),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29967),
            .lcout(\tok.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4403_3_lut_4_lut_LC_11_7_6 .C_ON=1'b0;
    defparam \tok.i4403_3_lut_4_lut_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i4403_3_lut_4_lut_LC_11_7_6 .LUT_INIT=16'b1111011111110111;
    LogicCell40 \tok.i4403_3_lut_4_lut_LC_11_7_6  (
            .in0(N__29682),
            .in1(N__29969),
            .in2(N__27927),
            .in3(_gnd_net_),
            .lcout(\tok.n4558 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_11_7_7 .C_ON=1'b0;
    defparam \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_11_7_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \tok.equal_130_i14_2_lut_3_lut_4_lut_LC_11_7_7  (
            .in0(N__28903),
            .in1(N__28739),
            .in2(N__28625),
            .in3(N__28401),
            .lcout(\tok.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_119_i11_2_lut_4_lut_LC_11_8_0 .C_ON=1'b0;
    defparam \tok.equal_119_i11_2_lut_4_lut_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \tok.equal_119_i11_2_lut_4_lut_LC_11_8_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \tok.equal_119_i11_2_lut_4_lut_LC_11_8_0  (
            .in0(N__29674),
            .in1(N__30279),
            .in2(N__27923),
            .in3(N__29962),
            .lcout(\tok.n11_adj_647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_1_lut_2_lut_4_lut_LC_11_8_1 .C_ON=1'b0;
    defparam \tok.i5_1_lut_2_lut_4_lut_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5_1_lut_2_lut_4_lut_LC_11_8_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \tok.i5_1_lut_2_lut_4_lut_LC_11_8_1  (
            .in0(N__29966),
            .in1(N__27879),
            .in2(N__30345),
            .in3(N__29680),
            .lcout(\tok.n9_adj_797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4315_2_lut_4_lut_LC_11_8_2 .C_ON=1'b0;
    defparam \tok.i4315_2_lut_4_lut_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \tok.i4315_2_lut_4_lut_LC_11_8_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \tok.i4315_2_lut_4_lut_LC_11_8_2  (
            .in0(N__29679),
            .in1(N__30282),
            .in2(N__27926),
            .in3(N__29965),
            .lcout(\tok.n4464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2534_2_lut_LC_11_8_3 .C_ON=1'b0;
    defparam \tok.i2534_2_lut_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2534_2_lut_LC_11_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.i2534_2_lut_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__29676),
            .in2(_gnd_net_),
            .in3(N__27868),
            .lcout(\tok.n2586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_121_i11_2_lut_4_lut_LC_11_8_4 .C_ON=1'b0;
    defparam \tok.equal_121_i11_2_lut_4_lut_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.equal_121_i11_2_lut_4_lut_LC_11_8_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.equal_121_i11_2_lut_4_lut_LC_11_8_4  (
            .in0(N__29677),
            .in1(N__30280),
            .in2(N__27924),
            .in3(N__29963),
            .lcout(\tok.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_4_lut_adj_154_LC_11_8_5 .C_ON=1'b0;
    defparam \tok.i1_2_lut_4_lut_adj_154_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_4_lut_adj_154_LC_11_8_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \tok.i1_2_lut_4_lut_adj_154_LC_11_8_5  (
            .in0(N__28906),
            .in1(N__28746),
            .in2(N__28634),
            .in3(N__28416),
            .lcout(\tok.n14_adj_825 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_114_i11_2_lut_4_lut_LC_11_8_6 .C_ON=1'b0;
    defparam \tok.equal_114_i11_2_lut_4_lut_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.equal_114_i11_2_lut_4_lut_LC_11_8_6 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \tok.equal_114_i11_2_lut_4_lut_LC_11_8_6  (
            .in0(N__29678),
            .in1(N__30281),
            .in2(N__27925),
            .in3(N__29964),
            .lcout(\tok.n11_adj_649 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_123_i10_2_lut_LC_11_8_7 .C_ON=1'b0;
    defparam \tok.equal_123_i10_2_lut_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.equal_123_i10_2_lut_LC_11_8_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.equal_123_i10_2_lut_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__27869),
            .in2(_gnd_net_),
            .in3(N__29675),
            .lcout(\tok.n10_adj_646 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4417_4_lut_4_lut_LC_11_9_0 .C_ON=1'b0;
    defparam \tok.i4417_4_lut_4_lut_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \tok.i4417_4_lut_4_lut_LC_11_9_0 .LUT_INIT=16'b1110111111010101;
    LogicCell40 \tok.i4417_4_lut_4_lut_LC_11_9_0  (
            .in0(N__30289),
            .in1(N__29684),
            .in2(N__27928),
            .in3(N__29973),
            .lcout(),
            .ltout(\tok.n4575_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_32_LC_11_9_1 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_32_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_32_LC_11_9_1 .LUT_INIT=16'b0011111110111111;
    LogicCell40 \tok.i3_4_lut_adj_32_LC_11_9_1  (
            .in0(N__23773),
            .in1(N__23801),
            .in2(N__23780),
            .in3(N__27266),
            .lcout(\tok.n4424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4373_4_lut_LC_11_9_2 .C_ON=1'b0;
    defparam \tok.i4373_4_lut_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \tok.i4373_4_lut_LC_11_9_2 .LUT_INIT=16'b1111111100111011;
    LogicCell40 \tok.i4373_4_lut_LC_11_9_2  (
            .in0(N__23756),
            .in1(N__26441),
            .in2(N__27596),
            .in3(N__27500),
            .lcout(\tok.n83 ),
            .ltout(\tok.n83_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2669_2_lut_LC_11_9_3 .C_ON=1'b0;
    defparam \tok.i2669_2_lut_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i2669_2_lut_LC_11_9_3 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \tok.i2669_2_lut_LC_11_9_3  (
            .in0(N__26730),
            .in1(_gnd_net_),
            .in2(N__23777),
            .in3(_gnd_net_),
            .lcout(\tok.n2746 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4413_4_lut_4_lut_LC_11_9_4 .C_ON=1'b0;
    defparam \tok.i4413_4_lut_4_lut_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i4413_4_lut_4_lut_LC_11_9_4 .LUT_INIT=16'b1110111111110011;
    LogicCell40 \tok.i4413_4_lut_4_lut_LC_11_9_4  (
            .in0(N__30291),
            .in1(N__29685),
            .in2(N__27930),
            .in3(N__29974),
            .lcout(),
            .ltout(\tok.n4571_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_34_LC_11_9_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_34_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_34_LC_11_9_5 .LUT_INIT=16'b1011111100111111;
    LogicCell40 \tok.i1_4_lut_adj_34_LC_11_9_5  (
            .in0(N__23774),
            .in1(N__29121),
            .in2(N__23759),
            .in3(N__28056),
            .lcout(\tok.n4393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_3_lut_3_lut_LC_11_9_6 .C_ON=1'b0;
    defparam \tok.i1_3_lut_3_lut_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_3_lut_3_lut_LC_11_9_6 .LUT_INIT=16'b1111101011110101;
    LogicCell40 \tok.i1_3_lut_3_lut_LC_11_9_6  (
            .in0(N__30290),
            .in1(_gnd_net_),
            .in2(N__27929),
            .in3(N__29975),
            .lcout(),
            .ltout(\tok.n4460_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2651_4_lut_LC_11_9_7 .C_ON=1'b0;
    defparam \tok.i2651_4_lut_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2651_4_lut_LC_11_9_7 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \tok.i2651_4_lut_LC_11_9_7  (
            .in0(N__27289),
            .in1(N__29122),
            .in2(N__24500),
            .in3(N__26455),
            .lcout(\tok.n2726 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_158_LC_11_10_0 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_158_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_158_LC_11_10_0 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \tok.i2_4_lut_adj_158_LC_11_10_0  (
            .in0(N__24659),
            .in1(N__29436),
            .in2(N__24393),
            .in3(N__28971),
            .lcout(),
            .ltout(\tok.n10_adj_829_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_162_LC_11_10_1 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_162_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_162_LC_11_10_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \tok.i5_4_lut_adj_162_LC_11_10_1  (
            .in0(N__30571),
            .in1(N__24293),
            .in2(N__24281),
            .in3(N__27188),
            .lcout(\tok.n13_adj_833 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_169_LC_11_10_2 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_169_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_169_LC_11_10_2 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \tok.i1_4_lut_adj_169_LC_11_10_2  (
            .in0(N__28001),
            .in1(N__30184),
            .in2(N__27218),
            .in3(N__24261),
            .lcout(\tok.n8_adj_839 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i6_4_lut_adj_55_LC_11_10_7 .C_ON=1'b0;
    defparam \tok.i6_4_lut_adj_55_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i6_4_lut_adj_55_LC_11_10_7 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \tok.i6_4_lut_adj_55_LC_11_10_7  (
            .in0(N__24068),
            .in1(N__24857),
            .in2(N__24226),
            .in3(N__27192),
            .lcout(\tok.n18_adj_681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.xor_103_i7_2_lut_LC_11_11_1 .C_ON=1'b0;
    defparam \tok.xor_103_i7_2_lut_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \tok.xor_103_i7_2_lut_LC_11_11_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tok.xor_103_i7_2_lut_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__24186),
            .in2(_gnd_net_),
            .in3(N__28543),
            .lcout(),
            .ltout(\tok.n244_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i5_4_lut_adj_122_LC_11_11_2 .C_ON=1'b0;
    defparam \tok.i5_4_lut_adj_122_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \tok.i5_4_lut_adj_122_LC_11_11_2 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \tok.i5_4_lut_adj_122_LC_11_11_2  (
            .in0(N__24069),
            .in1(N__23983),
            .in2(N__23912),
            .in3(N__24703),
            .lcout(\tok.n17_adj_785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.select_73_Select_13_i3_2_lut_LC_11_11_4 .C_ON=1'b0;
    defparam \tok.select_73_Select_13_i3_2_lut_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.select_73_Select_13_i3_2_lut_LC_11_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \tok.select_73_Select_13_i3_2_lut_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__24855),
            .in2(_gnd_net_),
            .in3(N__24704),
            .lcout(\tok.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_4_lut_adj_172_LC_11_11_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_4_lut_adj_172_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_4_lut_adj_172_LC_11_11_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \tok.i1_4_lut_4_lut_adj_172_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__28000),
            .in2(_gnd_net_),
            .in3(N__29782),
            .lcout(\tok.n40_adj_661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4329_2_lut_3_lut_LC_11_11_7 .C_ON=1'b0;
    defparam \tok.i4329_2_lut_3_lut_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \tok.i4329_2_lut_3_lut_LC_11_11_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \tok.i4329_2_lut_3_lut_LC_11_11_7  (
            .in0(N__30393),
            .in1(N__27530),
            .in2(_gnd_net_),
            .in3(N__30109),
            .lcout(\tok.n4478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i13_LC_12_3_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i13_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i13_LC_12_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i13_LC_12_3_0  (
            .in0(N__24533),
            .in1(N__24553),
            .in2(_gnd_net_),
            .in3(N__25639),
            .lcout(\tok.tail_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26249),
            .ce(N__25467),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i5_LC_12_3_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i5_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i5_LC_12_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i5_LC_12_3_1  (
            .in0(N__25638),
            .in1(N__24542),
            .in2(_gnd_net_),
            .in3(N__24590),
            .lcout(\tok.C_stk.tail_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26249),
            .ce(N__25467),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i21_LC_12_3_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i21_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i21_LC_12_3_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \tok.C_stk.tail_i0_i21_LC_12_3_2  (
            .in0(N__24541),
            .in1(_gnd_net_),
            .in2(N__24524),
            .in3(N__25640),
            .lcout(\tok.C_stk.tail_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26249),
            .ce(N__25467),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i29_LC_12_3_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i29_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i29_LC_12_3_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \tok.C_stk.tail_i0_i29_LC_12_3_3  (
            .in0(N__25636),
            .in1(N__24532),
            .in2(_gnd_net_),
            .in3(N__24509),
            .lcout(\tok.tail_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26249),
            .ce(N__25467),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i37_LC_12_3_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i37_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i37_LC_12_3_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i37_LC_12_3_4  (
            .in0(N__24520),
            .in1(N__25004),
            .in2(_gnd_net_),
            .in3(N__25641),
            .lcout(\tok.C_stk.tail_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26249),
            .ce(N__25467),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i45_LC_12_3_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i45_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i45_LC_12_3_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i45_LC_12_3_5  (
            .in0(N__25637),
            .in1(N__24985),
            .in2(_gnd_net_),
            .in3(N__24508),
            .lcout(\tok.tail_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26249),
            .ce(N__25467),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i53_LC_12_3_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i53_LC_12_3_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i53_LC_12_3_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i53_LC_12_3_6  (
            .in0(N__25016),
            .in1(N__25003),
            .in2(_gnd_net_),
            .in3(N__25642),
            .lcout(\tok.tail_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26249),
            .ce(N__25467),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i14_LC_12_3_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i14_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i14_LC_12_3_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i14_LC_12_3_7  (
            .in0(N__25635),
            .in1(N__24973),
            .in2(_gnd_net_),
            .in3(N__24952),
            .lcout(\tok.tail_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26249),
            .ce(N__25467),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i11_LC_12_4_0 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i11_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i11_LC_12_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i11_LC_12_4_0  (
            .in0(N__25716),
            .in1(N__24923),
            .in2(_gnd_net_),
            .in3(N__25132),
            .lcout(\tok.tail_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26254),
            .ce(N__25472),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i3_LC_12_4_1 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i3_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i3_LC_12_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.C_stk.tail_i0_i3_LC_12_4_1  (
            .in0(N__24932),
            .in1(N__25721),
            .in2(_gnd_net_),
            .in3(N__30487),
            .lcout(\tok.C_stk.tail_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26254),
            .ce(N__25472),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i19_LC_12_4_2 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i19_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i19_LC_12_4_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i19_LC_12_4_2  (
            .in0(N__25717),
            .in1(N__24914),
            .in2(_gnd_net_),
            .in3(N__24931),
            .lcout(\tok.C_stk.tail_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26254),
            .ce(N__25472),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i27_LC_12_4_3 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i27_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i27_LC_12_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \tok.C_stk.tail_i0_i27_LC_12_4_3  (
            .in0(N__24922),
            .in1(N__24905),
            .in2(_gnd_net_),
            .in3(N__25722),
            .lcout(\tok.tail_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26254),
            .ce(N__25472),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i35_LC_12_4_4 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i35_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i35_LC_12_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i35_LC_12_4_4  (
            .in0(N__25718),
            .in1(N__24884),
            .in2(_gnd_net_),
            .in3(N__24913),
            .lcout(\tok.C_stk.tail_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26254),
            .ce(N__25472),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i43_LC_12_4_5 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i43_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i43_LC_12_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \tok.C_stk.tail_i0_i43_LC_12_4_5  (
            .in0(N__24868),
            .in1(N__24904),
            .in2(_gnd_net_),
            .in3(N__25723),
            .lcout(\tok.tail_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26254),
            .ce(N__25472),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i51_LC_12_4_6 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i51_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i51_LC_12_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \tok.C_stk.tail_i0_i51_LC_12_4_6  (
            .in0(N__25719),
            .in1(N__24896),
            .in2(_gnd_net_),
            .in3(N__24883),
            .lcout(\tok.tail_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26254),
            .ce(N__25472),
            .sr(_gnd_net_));
    defparam \tok.C_stk.tail_i0_i2_LC_12_4_7 .C_ON=1'b0;
    defparam \tok.C_stk.tail_i0_i2_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.tail_i0_i2_LC_12_4_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \tok.C_stk.tail_i0_i2_LC_12_4_7  (
            .in0(N__25747),
            .in1(N__25720),
            .in2(_gnd_net_),
            .in3(N__25826),
            .lcout(\tok.C_stk.tail_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26254),
            .ce(N__25472),
            .sr(_gnd_net_));
    defparam \tok.C_stk.n602_bdd_4_lut_4734_LC_12_5_0 .C_ON=1'b0;
    defparam \tok.C_stk.n602_bdd_4_lut_4734_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.n602_bdd_4_lut_4734_LC_12_5_0 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \tok.C_stk.n602_bdd_4_lut_4734_LC_12_5_0  (
            .in0(N__26322),
            .in1(N__25297),
            .in2(N__25105),
            .in3(N__25364),
            .lcout(),
            .ltout(\tok.C_stk.n4888_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i4_LC_12_5_1 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i4_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i4_LC_12_5_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \tok.C_stk.head_i0_i4_LC_12_5_1  (
            .in0(N__25334),
            .in1(N__30536),
            .in2(N__25316),
            .in3(N__26324),
            .lcout(\tok.c_stk_r_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26260),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i4650_4_lut_LC_12_5_2 .C_ON=1'b0;
    defparam \tok.ram.i4650_4_lut_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i4650_4_lut_LC_12_5_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.ram.i4650_4_lut_LC_12_5_2  (
            .in0(N__26682),
            .in1(N__25295),
            .in2(N__30539),
            .in3(N__26000),
            .lcout(),
            .ltout(\tok.ram.n4705_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5_4_lut_adj_23_LC_12_5_3 .C_ON=1'b0;
    defparam \tok.ram.i5_4_lut_adj_23_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5_4_lut_adj_23_LC_12_5_3 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \tok.ram.i5_4_lut_adj_23_LC_12_5_3  (
            .in0(N__29851),
            .in1(N__30535),
            .in2(N__25313),
            .in3(N__25910),
            .lcout(),
            .ltout(\tok.n1_adj_745_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_92_LC_12_5_4 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_92_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_92_LC_12_5_4 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i27_4_lut_adj_92_LC_12_5_4  (
            .in0(N__27704),
            .in1(N__28556),
            .in2(N__25310),
            .in3(N__30153),
            .lcout(),
            .ltout(\tok.n13_adj_746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_93_LC_12_5_5 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_93_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_93_LC_12_5_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \tok.i1_4_lut_adj_93_LC_12_5_5  (
            .in0(N__25296),
            .in1(N__25277),
            .in2(N__25208),
            .in3(N__25202),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i3_LC_12_5_6 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i3_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i3_LC_12_5_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \tok.C_stk.head_i0_i3_LC_12_5_6  (
            .in0(N__26323),
            .in1(N__25133),
            .in2(N__25121),
            .in3(N__30488),
            .lcout(\tok.c_stk_r_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26260),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.n602_bdd_4_lut_4724_LC_12_6_0 .C_ON=1'b0;
    defparam \tok.C_stk.n602_bdd_4_lut_4724_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \tok.C_stk.n602_bdd_4_lut_4724_LC_12_6_0 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \tok.C_stk.n602_bdd_4_lut_4724_LC_12_6_0  (
            .in0(N__26330),
            .in1(N__26031),
            .in2(N__25111),
            .in3(N__25042),
            .lcout(),
            .ltout(\tok.C_stk.n4876_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.C_stk.head_i0_i2_LC_12_6_1 .C_ON=1'b0;
    defparam \tok.C_stk.head_i0_i2_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \tok.C_stk.head_i0_i2_LC_12_6_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \tok.C_stk.head_i0_i2_LC_12_6_1  (
            .in0(N__26378),
            .in1(N__25821),
            .in2(N__26363),
            .in3(N__26331),
            .lcout(\tok.c_stk_r_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26262),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i4658_4_lut_LC_12_6_2 .C_ON=1'b0;
    defparam \tok.ram.i4658_4_lut_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i4658_4_lut_LC_12_6_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \tok.ram.i4658_4_lut_LC_12_6_2  (
            .in0(N__26673),
            .in1(N__26030),
            .in2(N__25825),
            .in3(N__25979),
            .lcout(),
            .ltout(\tok.ram.n4711_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5_4_lut_adj_21_LC_12_6_3 .C_ON=1'b0;
    defparam \tok.ram.i5_4_lut_adj_21_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5_4_lut_adj_21_LC_12_6_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \tok.ram.i5_4_lut_adj_21_LC_12_6_3  (
            .in0(N__25909),
            .in1(N__25820),
            .in2(N__25922),
            .in3(N__29863),
            .lcout(),
            .ltout(\tok.n1_adj_724_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i27_4_lut_adj_78_LC_12_6_4 .C_ON=1'b0;
    defparam \tok.i27_4_lut_adj_78_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \tok.i27_4_lut_adj_78_LC_12_6_4 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \tok.i27_4_lut_adj_78_LC_12_6_4  (
            .in0(N__25757),
            .in1(N__28532),
            .in2(N__25919),
            .in3(N__30136),
            .lcout(\tok.n13_adj_725 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i5_4_lut_adj_22_LC_12_6_5 .C_ON=1'b0;
    defparam \tok.ram.i5_4_lut_adj_22_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i5_4_lut_adj_22_LC_12_6_5 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \tok.ram.i5_4_lut_adj_22_LC_12_6_5  (
            .in0(N__25908),
            .in1(N__25844),
            .in2(N__30493),
            .in3(N__29862),
            .lcout(\tok.n1_adj_736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i18_4_lut_adj_87_LC_12_7_0 .C_ON=1'b0;
    defparam \tok.i18_4_lut_adj_87_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \tok.i18_4_lut_adj_87_LC_12_7_0 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \tok.i18_4_lut_adj_87_LC_12_7_0  (
            .in0(N__30105),
            .in1(N__25838),
            .in2(N__29606),
            .in3(N__28459),
            .lcout(\tok.n5_adj_737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_75_LC_12_7_1 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_75_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_75_LC_12_7_1 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \tok.i125_4_lut_adj_75_LC_12_7_1  (
            .in0(N__30384),
            .in1(N__25816),
            .in2(N__25796),
            .in3(N__30104),
            .lcout(),
            .ltout(\tok.n83_adj_721_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4632_2_lut_3_lut_LC_12_7_2 .C_ON=1'b0;
    defparam \tok.i4632_2_lut_3_lut_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.i4632_2_lut_3_lut_LC_12_7_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \tok.i4632_2_lut_3_lut_LC_12_7_2  (
            .in0(N__29859),
            .in1(_gnd_net_),
            .in2(N__25760),
            .in3(N__28941),
            .lcout(\tok.n4692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i2_4_lut_4_lut_LC_12_7_3 .C_ON=1'b0;
    defparam \tok.ram.i2_4_lut_4_lut_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i2_4_lut_4_lut_LC_12_7_3 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \tok.ram.i2_4_lut_4_lut_LC_12_7_3  (
            .in0(N__30381),
            .in1(N__29858),
            .in2(N__28012),
            .in3(N__30102),
            .lcout(),
            .ltout(\tok.ram.n14_adj_631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i2581_4_lut_LC_12_7_4 .C_ON=1'b0;
    defparam \tok.ram.i2581_4_lut_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i2581_4_lut_LC_12_7_4 .LUT_INIT=16'b1110111011101010;
    LogicCell40 \tok.ram.i2581_4_lut_LC_12_7_4  (
            .in0(N__26497),
            .in1(N__27556),
            .in2(N__26819),
            .in3(N__28057),
            .lcout(\tok.n2635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_130_LC_12_7_5 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_130_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_130_LC_12_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i1_2_lut_adj_130_LC_12_7_5  (
            .in0(N__30383),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28940),
            .lcout(\tok.n4_adj_795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_adj_150_LC_12_7_6 .C_ON=1'b0;
    defparam \tok.i1_2_lut_adj_150_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_adj_150_LC_12_7_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \tok.i1_2_lut_adj_150_LC_12_7_6  (
            .in0(N__30103),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30382),
            .lcout(\tok.n41 ),
            .ltout(\tok.n41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_adj_45_LC_12_7_7 .C_ON=1'b0;
    defparam \tok.i2_4_lut_adj_45_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_adj_45_LC_12_7_7 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \tok.i2_4_lut_adj_45_LC_12_7_7  (
            .in0(N__28058),
            .in1(N__29597),
            .in2(N__26627),
            .in3(N__28939),
            .lcout(\tok.n884 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_157_i15_2_lut_3_lut_LC_12_8_1 .C_ON=1'b0;
    defparam \tok.equal_157_i15_2_lut_3_lut_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \tok.equal_157_i15_2_lut_3_lut_LC_12_8_1 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \tok.equal_157_i15_2_lut_3_lut_LC_12_8_1  (
            .in0(N__28055),
            .in1(N__28103),
            .in2(_gnd_net_),
            .in3(N__26498),
            .lcout(\tok.n15_adj_662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4415_4_lut_LC_12_8_3 .C_ON=1'b0;
    defparam \tok.i4415_4_lut_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4415_4_lut_LC_12_8_3 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \tok.i4415_4_lut_LC_12_8_3  (
            .in0(N__28104),
            .in1(N__27528),
            .in2(N__26456),
            .in3(N__27267),
            .lcout(\tok.n4573 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2_4_lut_LC_12_8_4 .C_ON=1'b0;
    defparam \tok.i2_4_lut_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \tok.i2_4_lut_LC_12_8_4 .LUT_INIT=16'b0100110011111111;
    LogicCell40 \tok.i2_4_lut_LC_12_8_4  (
            .in0(N__28102),
            .in1(N__28054),
            .in2(N__26434),
            .in3(N__26397),
            .lcout(),
            .ltout(\tok.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_LC_12_8_5 .C_ON=1'b0;
    defparam \tok.i3_4_lut_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_LC_12_8_5 .LUT_INIT=16'b1111010011110101;
    LogicCell40 \tok.i3_4_lut_LC_12_8_5  (
            .in0(N__27690),
            .in1(N__30352),
            .in2(N__26381),
            .in3(N__30044),
            .lcout(),
            .ltout(\tok.n4422_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_33_LC_12_8_6 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_33_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_33_LC_12_8_6 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \tok.i1_4_lut_adj_33_LC_12_8_6  (
            .in0(N__27589),
            .in1(N__27538),
            .in2(N__27578),
            .in3(N__27555),
            .lcout(),
            .ltout(\tok.n51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_4_lut_adj_36_LC_12_8_7 .C_ON=1'b0;
    defparam \tok.i1_4_lut_adj_36_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_4_lut_adj_36_LC_12_8_7 .LUT_INIT=16'b1111001111110001;
    LogicCell40 \tok.i1_4_lut_adj_36_LC_12_8_7  (
            .in0(N__27539),
            .in1(N__27529),
            .in2(N__27509),
            .in3(N__27506),
            .lcout(\tok.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_adj_60_LC_12_9_3 .C_ON=1'b0;
    defparam \tok.i3_3_lut_adj_60_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_adj_60_LC_12_9_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \tok.i3_3_lut_adj_60_LC_12_9_3  (
            .in0(N__27494),
            .in1(N__27479),
            .in2(_gnd_net_),
            .in3(N__27168),
            .lcout(),
            .ltout(\tok.n14_adj_695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_adj_62_LC_12_9_4 .C_ON=1'b0;
    defparam \tok.i7_4_lut_adj_62_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_adj_62_LC_12_9_4 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \tok.i7_4_lut_adj_62_LC_12_9_4  (
            .in0(N__27045),
            .in1(N__27470),
            .in2(N__27455),
            .in3(N__27448),
            .lcout(\tok.n18_adj_698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i2458_2_lut_LC_12_9_5 .C_ON=1'b0;
    defparam \tok.i2458_2_lut_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \tok.i2458_2_lut_LC_12_9_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \tok.i2458_2_lut_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__30412),
            .in2(_gnd_net_),
            .in3(N__30113),
            .lcout(\tok.n2177 ),
            .ltout(\tok.n2177_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.ram.i1_3_lut_LC_12_9_6 .C_ON=1'b0;
    defparam \tok.ram.i1_3_lut_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \tok.ram.i1_3_lut_LC_12_9_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \tok.ram.i1_3_lut_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__27290),
            .in2(N__27278),
            .in3(N__27268),
            .lcout(\tok.n132 ),
            .ltout(\tok.n132_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_LC_12_9_7 .C_ON=1'b0;
    defparam \tok.i3_3_lut_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_LC_12_9_7 .LUT_INIT=16'b1111111100001100;
    LogicCell40 \tok.i3_3_lut_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__27122),
            .in2(N__27110),
            .in3(N__27107),
            .lcout(\tok.n14_adj_651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i7_4_lut_LC_12_10_0 .C_ON=1'b0;
    defparam \tok.i7_4_lut_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \tok.i7_4_lut_LC_12_10_0 .LUT_INIT=16'b1110111111101110;
    LogicCell40 \tok.i7_4_lut_LC_12_10_0  (
            .in0(N__27098),
            .in1(N__27083),
            .in2(N__27061),
            .in3(N__26933),
            .lcout(\tok.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.or_99_i11_2_lut_LC_12_10_4 .C_ON=1'b0;
    defparam \tok.or_99_i11_2_lut_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \tok.or_99_i11_2_lut_LC_12_10_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \tok.or_99_i11_2_lut_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__28299),
            .in2(_gnd_net_),
            .in3(N__28260),
            .lcout(\tok.n179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_117_i10_2_lut_LC_12_10_5 .C_ON=1'b0;
    defparam \tok.equal_117_i10_2_lut_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \tok.equal_117_i10_2_lut_LC_12_10_5 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \tok.equal_117_i10_2_lut_LC_12_10_5  (
            .in0(N__27979),
            .in1(N__29802),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tok.n10_adj_675 ),
            .ltout(\tok.n10_adj_675_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4335_3_lut_4_lut_4_lut_LC_12_10_6 .C_ON=1'b0;
    defparam \tok.i4335_3_lut_4_lut_4_lut_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \tok.i4335_3_lut_4_lut_4_lut_LC_12_10_6 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \tok.i4335_3_lut_4_lut_4_lut_LC_12_10_6  (
            .in0(N__27762),
            .in1(N__28116),
            .in2(N__28079),
            .in3(N__28073),
            .lcout(\tok.n4484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_4_lut_adj_152_LC_12_10_7 .C_ON=1'b0;
    defparam \tok.i1_2_lut_4_lut_adj_152_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_4_lut_adj_152_LC_12_10_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \tok.i1_2_lut_4_lut_adj_152_LC_12_10_7  (
            .in0(N__30392),
            .in1(N__29801),
            .in2(N__28011),
            .in3(N__30110),
            .lcout(\tok.n2178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_4_lut_adj_42_LC_12_11_6 .C_ON=1'b0;
    defparam \tok.i3_4_lut_adj_42_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \tok.i3_4_lut_adj_42_LC_12_11_6 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \tok.i3_4_lut_adj_42_LC_12_11_6  (
            .in0(N__27737),
            .in1(N__27728),
            .in2(N__27722),
            .in3(N__27698),
            .lcout(\tok.n42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4585_2_lut_3_lut_LC_13_6_3 .C_ON=1'b0;
    defparam \tok.i4585_2_lut_3_lut_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \tok.i4585_2_lut_3_lut_LC_13_6_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \tok.i4585_2_lut_3_lut_LC_13_6_3  (
            .in0(N__30500),
            .in1(N__28990),
            .in2(_gnd_net_),
            .in3(N__29860),
            .lcout(\tok.n4688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.T_7__I_0_233_i14_2_lut_3_lut_4_lut_LC_13_7_1 .C_ON=1'b0;
    defparam \tok.T_7__I_0_233_i14_2_lut_3_lut_4_lut_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \tok.T_7__I_0_233_i14_2_lut_3_lut_4_lut_LC_13_7_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \tok.T_7__I_0_233_i14_2_lut_3_lut_4_lut_LC_13_7_1  (
            .in0(N__28449),
            .in1(N__28626),
            .in2(N__28807),
            .in3(N__28934),
            .lcout(\tok.n14_adj_658 ),
            .ltout(\tok.n14_adj_658_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.equal_154_i16_3_lut_4_lut_LC_13_7_2 .C_ON=1'b0;
    defparam \tok.equal_154_i16_3_lut_4_lut_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \tok.equal_154_i16_3_lut_4_lut_LC_13_7_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \tok.equal_154_i16_3_lut_4_lut_LC_13_7_2  (
            .in0(N__27691),
            .in1(N__30385),
            .in2(N__27671),
            .in3(N__30106),
            .lcout(\tok.n399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_90_LC_13_7_3 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_90_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_90_LC_13_7_3 .LUT_INIT=16'b0100101001000000;
    LogicCell40 \tok.i125_4_lut_adj_90_LC_13_7_3  (
            .in0(N__30107),
            .in1(N__30572),
            .in2(N__30418),
            .in3(N__30537),
            .lcout(\tok.n83_adj_743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i125_4_lut_adj_84_LC_13_7_4 .C_ON=1'b0;
    defparam \tok.i125_4_lut_adj_84_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \tok.i125_4_lut_adj_84_LC_13_7_4 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \tok.i125_4_lut_adj_84_LC_13_7_4  (
            .in0(N__30494),
            .in1(N__30389),
            .in2(N__30194),
            .in3(N__30108),
            .lcout(),
            .ltout(\tok.n83_adj_733_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4584_2_lut_3_lut_LC_13_7_5 .C_ON=1'b0;
    defparam \tok.i4584_2_lut_3_lut_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \tok.i4584_2_lut_3_lut_LC_13_7_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \tok.i4584_2_lut_3_lut_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__28935),
            .in2(N__29876),
            .in3(N__29861),
            .lcout(\tok.n4627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i1_2_lut_3_lut_LC_13_7_6 .C_ON=1'b0;
    defparam \tok.i1_2_lut_3_lut_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \tok.i1_2_lut_3_lut_LC_13_7_6 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \tok.i1_2_lut_3_lut_LC_13_7_6  (
            .in0(N__28627),
            .in1(N__28775),
            .in2(_gnd_net_),
            .in3(N__28450),
            .lcout(\tok.n883 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i3_3_lut_adj_53_LC_13_7_7 .C_ON=1'b0;
    defparam \tok.i3_3_lut_adj_53_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \tok.i3_3_lut_adj_53_LC_13_7_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \tok.i3_3_lut_adj_53_LC_13_7_7  (
            .in0(N__29591),
            .in1(N__29573),
            .in2(_gnd_net_),
            .in3(N__29457),
            .lcout(\tok.n15_adj_680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i4710_2_lut_LC_13_8_7 .C_ON=1'b0;
    defparam \tok.i4710_2_lut_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \tok.i4710_2_lut_LC_13_8_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \tok.i4710_2_lut_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__29149),
            .in2(_gnd_net_),
            .in3(N__29126),
            .lcout(\tok.write_flag ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tok.i244_2_lut_3_lut_4_lut_LC_13_11_4 .C_ON=1'b0;
    defparam \tok.i244_2_lut_3_lut_4_lut_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \tok.i244_2_lut_3_lut_4_lut_LC_13_11_4 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \tok.i244_2_lut_3_lut_4_lut_LC_13_11_4  (
            .in0(N__28989),
            .in1(N__28830),
            .in2(N__28699),
            .in3(N__28542),
            .lcout(\tok.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
